VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 1100.000 ;
  PIN custom_settings[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.720 4.000 596.320 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 606.600 4.000 607.200 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.920 4.000 623.520 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.800 4.000 498.400 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.680 4.000 509.280 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.120 4.000 514.720 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.000 4.000 525.600 ;
    END
  END custom_settings[9]
  PIN io_in_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 10.210 1096.000 10.490 1100.000 ;
    END
  END io_in_0
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 253.000 4.000 253.600 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END io_oeb[9]
  PIN io_oeb_6502
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 353.640 200.000 354.240 ;
    END
  END io_oeb_6502
  PIN io_oeb_as1802
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 946.600 200.000 947.200 ;
    END
  END io_oeb_as1802
  PIN io_oeb_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END io_oeb_scrapcpu[0]
  PIN io_oeb_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 900.360 4.000 900.960 ;
    END
  END io_oeb_scrapcpu[10]
  PIN io_oeb_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 905.800 4.000 906.400 ;
    END
  END io_oeb_scrapcpu[11]
  PIN io_oeb_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END io_oeb_scrapcpu[12]
  PIN io_oeb_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 916.680 4.000 917.280 ;
    END
  END io_oeb_scrapcpu[13]
  PIN io_oeb_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.120 4.000 922.720 ;
    END
  END io_oeb_scrapcpu[14]
  PIN io_oeb_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 927.560 4.000 928.160 ;
    END
  END io_oeb_scrapcpu[15]
  PIN io_oeb_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.000 4.000 933.600 ;
    END
  END io_oeb_scrapcpu[16]
  PIN io_oeb_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 938.440 4.000 939.040 ;
    END
  END io_oeb_scrapcpu[17]
  PIN io_oeb_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.880 4.000 944.480 ;
    END
  END io_oeb_scrapcpu[18]
  PIN io_oeb_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 949.320 4.000 949.920 ;
    END
  END io_oeb_scrapcpu[19]
  PIN io_oeb_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 851.400 4.000 852.000 ;
    END
  END io_oeb_scrapcpu[1]
  PIN io_oeb_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 954.760 4.000 955.360 ;
    END
  END io_oeb_scrapcpu[20]
  PIN io_oeb_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END io_oeb_scrapcpu[21]
  PIN io_oeb_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END io_oeb_scrapcpu[22]
  PIN io_oeb_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 971.080 4.000 971.680 ;
    END
  END io_oeb_scrapcpu[23]
  PIN io_oeb_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 976.520 4.000 977.120 ;
    END
  END io_oeb_scrapcpu[24]
  PIN io_oeb_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 981.960 4.000 982.560 ;
    END
  END io_oeb_scrapcpu[25]
  PIN io_oeb_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 987.400 4.000 988.000 ;
    END
  END io_oeb_scrapcpu[26]
  PIN io_oeb_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END io_oeb_scrapcpu[27]
  PIN io_oeb_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 998.280 4.000 998.880 ;
    END
  END io_oeb_scrapcpu[28]
  PIN io_oeb_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1003.720 4.000 1004.320 ;
    END
  END io_oeb_scrapcpu[29]
  PIN io_oeb_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END io_oeb_scrapcpu[2]
  PIN io_oeb_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.160 4.000 1009.760 ;
    END
  END io_oeb_scrapcpu[30]
  PIN io_oeb_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1014.600 4.000 1015.200 ;
    END
  END io_oeb_scrapcpu[31]
  PIN io_oeb_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.040 4.000 1020.640 ;
    END
  END io_oeb_scrapcpu[32]
  PIN io_oeb_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END io_oeb_scrapcpu[33]
  PIN io_oeb_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.920 4.000 1031.520 ;
    END
  END io_oeb_scrapcpu[34]
  PIN io_oeb_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END io_oeb_scrapcpu[35]
  PIN io_oeb_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END io_oeb_scrapcpu[3]
  PIN io_oeb_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END io_oeb_scrapcpu[4]
  PIN io_oeb_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END io_oeb_scrapcpu[5]
  PIN io_oeb_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END io_oeb_scrapcpu[6]
  PIN io_oeb_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END io_oeb_scrapcpu[7]
  PIN io_oeb_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 889.480 4.000 890.080 ;
    END
  END io_oeb_scrapcpu[8]
  PIN io_oeb_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.920 4.000 895.520 ;
    END
  END io_oeb_scrapcpu[9]
  PIN io_oeb_vliw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END io_oeb_vliw[0]
  PIN io_oeb_vliw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END io_oeb_vliw[10]
  PIN io_oeb_vliw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END io_oeb_vliw[11]
  PIN io_oeb_vliw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END io_oeb_vliw[12]
  PIN io_oeb_vliw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END io_oeb_vliw[13]
  PIN io_oeb_vliw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.280 4.000 726.880 ;
    END
  END io_oeb_vliw[14]
  PIN io_oeb_vliw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END io_oeb_vliw[15]
  PIN io_oeb_vliw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.160 4.000 737.760 ;
    END
  END io_oeb_vliw[16]
  PIN io_oeb_vliw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 742.600 4.000 743.200 ;
    END
  END io_oeb_vliw[17]
  PIN io_oeb_vliw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END io_oeb_vliw[18]
  PIN io_oeb_vliw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 753.480 4.000 754.080 ;
    END
  END io_oeb_vliw[19]
  PIN io_oeb_vliw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END io_oeb_vliw[1]
  PIN io_oeb_vliw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.920 4.000 759.520 ;
    END
  END io_oeb_vliw[20]
  PIN io_oeb_vliw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END io_oeb_vliw[21]
  PIN io_oeb_vliw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END io_oeb_vliw[22]
  PIN io_oeb_vliw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END io_oeb_vliw[23]
  PIN io_oeb_vliw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END io_oeb_vliw[24]
  PIN io_oeb_vliw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END io_oeb_vliw[25]
  PIN io_oeb_vliw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 791.560 4.000 792.160 ;
    END
  END io_oeb_vliw[26]
  PIN io_oeb_vliw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END io_oeb_vliw[27]
  PIN io_oeb_vliw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END io_oeb_vliw[28]
  PIN io_oeb_vliw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END io_oeb_vliw[29]
  PIN io_oeb_vliw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END io_oeb_vliw[2]
  PIN io_oeb_vliw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END io_oeb_vliw[30]
  PIN io_oeb_vliw[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 818.760 4.000 819.360 ;
    END
  END io_oeb_vliw[31]
  PIN io_oeb_vliw[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END io_oeb_vliw[32]
  PIN io_oeb_vliw[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END io_oeb_vliw[33]
  PIN io_oeb_vliw[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 835.080 4.000 835.680 ;
    END
  END io_oeb_vliw[34]
  PIN io_oeb_vliw[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 4.000 841.120 ;
    END
  END io_oeb_vliw[35]
  PIN io_oeb_vliw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END io_oeb_vliw[3]
  PIN io_oeb_vliw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END io_oeb_vliw[4]
  PIN io_oeb_vliw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END io_oeb_vliw[5]
  PIN io_oeb_vliw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END io_oeb_vliw[6]
  PIN io_oeb_vliw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END io_oeb_vliw[7]
  PIN io_oeb_vliw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END io_oeb_vliw[8]
  PIN io_oeb_vliw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END io_oeb_vliw[9]
  PIN io_oeb_z80[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 652.840 200.000 653.440 ;
    END
  END io_oeb_z80[0]
  PIN io_oeb_z80[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 680.040 200.000 680.640 ;
    END
  END io_oeb_z80[10]
  PIN io_oeb_z80[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 682.760 200.000 683.360 ;
    END
  END io_oeb_z80[11]
  PIN io_oeb_z80[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 685.480 200.000 686.080 ;
    END
  END io_oeb_z80[12]
  PIN io_oeb_z80[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 688.200 200.000 688.800 ;
    END
  END io_oeb_z80[13]
  PIN io_oeb_z80[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 690.920 200.000 691.520 ;
    END
  END io_oeb_z80[14]
  PIN io_oeb_z80[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 693.640 200.000 694.240 ;
    END
  END io_oeb_z80[15]
  PIN io_oeb_z80[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 696.360 200.000 696.960 ;
    END
  END io_oeb_z80[16]
  PIN io_oeb_z80[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 699.080 200.000 699.680 ;
    END
  END io_oeb_z80[17]
  PIN io_oeb_z80[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 701.800 200.000 702.400 ;
    END
  END io_oeb_z80[18]
  PIN io_oeb_z80[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 704.520 200.000 705.120 ;
    END
  END io_oeb_z80[19]
  PIN io_oeb_z80[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 655.560 200.000 656.160 ;
    END
  END io_oeb_z80[1]
  PIN io_oeb_z80[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 707.240 200.000 707.840 ;
    END
  END io_oeb_z80[20]
  PIN io_oeb_z80[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 709.960 200.000 710.560 ;
    END
  END io_oeb_z80[21]
  PIN io_oeb_z80[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 712.680 200.000 713.280 ;
    END
  END io_oeb_z80[22]
  PIN io_oeb_z80[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 715.400 200.000 716.000 ;
    END
  END io_oeb_z80[23]
  PIN io_oeb_z80[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 718.120 200.000 718.720 ;
    END
  END io_oeb_z80[24]
  PIN io_oeb_z80[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 720.840 200.000 721.440 ;
    END
  END io_oeb_z80[25]
  PIN io_oeb_z80[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 723.560 200.000 724.160 ;
    END
  END io_oeb_z80[26]
  PIN io_oeb_z80[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 726.280 200.000 726.880 ;
    END
  END io_oeb_z80[27]
  PIN io_oeb_z80[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 729.000 200.000 729.600 ;
    END
  END io_oeb_z80[28]
  PIN io_oeb_z80[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 731.720 200.000 732.320 ;
    END
  END io_oeb_z80[29]
  PIN io_oeb_z80[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 658.280 200.000 658.880 ;
    END
  END io_oeb_z80[2]
  PIN io_oeb_z80[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 734.440 200.000 735.040 ;
    END
  END io_oeb_z80[30]
  PIN io_oeb_z80[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 737.160 200.000 737.760 ;
    END
  END io_oeb_z80[31]
  PIN io_oeb_z80[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 739.880 200.000 740.480 ;
    END
  END io_oeb_z80[32]
  PIN io_oeb_z80[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 742.600 200.000 743.200 ;
    END
  END io_oeb_z80[33]
  PIN io_oeb_z80[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 745.320 200.000 745.920 ;
    END
  END io_oeb_z80[34]
  PIN io_oeb_z80[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 748.040 200.000 748.640 ;
    END
  END io_oeb_z80[35]
  PIN io_oeb_z80[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 661.000 200.000 661.600 ;
    END
  END io_oeb_z80[3]
  PIN io_oeb_z80[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 663.720 200.000 664.320 ;
    END
  END io_oeb_z80[4]
  PIN io_oeb_z80[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 666.440 200.000 667.040 ;
    END
  END io_oeb_z80[5]
  PIN io_oeb_z80[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 669.160 200.000 669.760 ;
    END
  END io_oeb_z80[6]
  PIN io_oeb_z80[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 671.880 200.000 672.480 ;
    END
  END io_oeb_z80[7]
  PIN io_oeb_z80[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 674.600 200.000 675.200 ;
    END
  END io_oeb_z80[8]
  PIN io_oeb_z80[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 677.320 200.000 677.920 ;
    END
  END io_oeb_z80[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 152.360 200.000 152.960 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 179.560 200.000 180.160 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 182.280 200.000 182.880 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 185.000 200.000 185.600 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.720 200.000 188.320 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 190.440 200.000 191.040 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 193.160 200.000 193.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 195.880 200.000 196.480 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 198.600 200.000 199.200 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 201.320 200.000 201.920 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 204.040 200.000 204.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 155.080 200.000 155.680 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 206.760 200.000 207.360 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 209.480 200.000 210.080 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 212.200 200.000 212.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 214.920 200.000 215.520 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 217.640 200.000 218.240 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 220.360 200.000 220.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 223.080 200.000 223.680 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 225.800 200.000 226.400 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 228.520 200.000 229.120 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 231.240 200.000 231.840 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 157.800 200.000 158.400 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 233.960 200.000 234.560 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 236.680 200.000 237.280 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 239.400 200.000 240.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 242.120 200.000 242.720 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 244.840 200.000 245.440 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 247.560 200.000 248.160 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 250.280 200.000 250.880 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 253.000 200.000 253.600 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 160.520 200.000 161.120 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 163.240 200.000 163.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 165.960 200.000 166.560 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 200.000 169.280 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 171.400 200.000 172.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 174.120 200.000 174.720 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.840 200.000 177.440 ;
    END
  END io_out[9]
  PIN io_out_6502[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 255.720 200.000 256.320 ;
    END
  END io_out_6502[0]
  PIN io_out_6502[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 282.920 200.000 283.520 ;
    END
  END io_out_6502[10]
  PIN io_out_6502[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 285.640 200.000 286.240 ;
    END
  END io_out_6502[11]
  PIN io_out_6502[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 288.360 200.000 288.960 ;
    END
  END io_out_6502[12]
  PIN io_out_6502[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 291.080 200.000 291.680 ;
    END
  END io_out_6502[13]
  PIN io_out_6502[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 293.800 200.000 294.400 ;
    END
  END io_out_6502[14]
  PIN io_out_6502[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 296.520 200.000 297.120 ;
    END
  END io_out_6502[15]
  PIN io_out_6502[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 299.240 200.000 299.840 ;
    END
  END io_out_6502[16]
  PIN io_out_6502[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 301.960 200.000 302.560 ;
    END
  END io_out_6502[17]
  PIN io_out_6502[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 304.680 200.000 305.280 ;
    END
  END io_out_6502[18]
  PIN io_out_6502[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 307.400 200.000 308.000 ;
    END
  END io_out_6502[19]
  PIN io_out_6502[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 258.440 200.000 259.040 ;
    END
  END io_out_6502[1]
  PIN io_out_6502[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 310.120 200.000 310.720 ;
    END
  END io_out_6502[20]
  PIN io_out_6502[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 312.840 200.000 313.440 ;
    END
  END io_out_6502[21]
  PIN io_out_6502[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 315.560 200.000 316.160 ;
    END
  END io_out_6502[22]
  PIN io_out_6502[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 318.280 200.000 318.880 ;
    END
  END io_out_6502[23]
  PIN io_out_6502[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 321.000 200.000 321.600 ;
    END
  END io_out_6502[24]
  PIN io_out_6502[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 323.720 200.000 324.320 ;
    END
  END io_out_6502[25]
  PIN io_out_6502[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 326.440 200.000 327.040 ;
    END
  END io_out_6502[26]
  PIN io_out_6502[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 329.160 200.000 329.760 ;
    END
  END io_out_6502[27]
  PIN io_out_6502[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 331.880 200.000 332.480 ;
    END
  END io_out_6502[28]
  PIN io_out_6502[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 334.600 200.000 335.200 ;
    END
  END io_out_6502[29]
  PIN io_out_6502[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 261.160 200.000 261.760 ;
    END
  END io_out_6502[2]
  PIN io_out_6502[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 337.320 200.000 337.920 ;
    END
  END io_out_6502[30]
  PIN io_out_6502[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 340.040 200.000 340.640 ;
    END
  END io_out_6502[31]
  PIN io_out_6502[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 342.760 200.000 343.360 ;
    END
  END io_out_6502[32]
  PIN io_out_6502[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 345.480 200.000 346.080 ;
    END
  END io_out_6502[33]
  PIN io_out_6502[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 348.200 200.000 348.800 ;
    END
  END io_out_6502[34]
  PIN io_out_6502[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 350.920 200.000 351.520 ;
    END
  END io_out_6502[35]
  PIN io_out_6502[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 263.880 200.000 264.480 ;
    END
  END io_out_6502[3]
  PIN io_out_6502[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 266.600 200.000 267.200 ;
    END
  END io_out_6502[4]
  PIN io_out_6502[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 269.320 200.000 269.920 ;
    END
  END io_out_6502[5]
  PIN io_out_6502[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 272.040 200.000 272.640 ;
    END
  END io_out_6502[6]
  PIN io_out_6502[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 274.760 200.000 275.360 ;
    END
  END io_out_6502[7]
  PIN io_out_6502[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 277.480 200.000 278.080 ;
    END
  END io_out_6502[8]
  PIN io_out_6502[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 280.200 200.000 280.800 ;
    END
  END io_out_6502[9]
  PIN io_out_as1802[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 848.680 200.000 849.280 ;
    END
  END io_out_as1802[0]
  PIN io_out_as1802[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 875.880 200.000 876.480 ;
    END
  END io_out_as1802[10]
  PIN io_out_as1802[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 878.600 200.000 879.200 ;
    END
  END io_out_as1802[11]
  PIN io_out_as1802[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 881.320 200.000 881.920 ;
    END
  END io_out_as1802[12]
  PIN io_out_as1802[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 884.040 200.000 884.640 ;
    END
  END io_out_as1802[13]
  PIN io_out_as1802[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 886.760 200.000 887.360 ;
    END
  END io_out_as1802[14]
  PIN io_out_as1802[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 889.480 200.000 890.080 ;
    END
  END io_out_as1802[15]
  PIN io_out_as1802[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 892.200 200.000 892.800 ;
    END
  END io_out_as1802[16]
  PIN io_out_as1802[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 894.920 200.000 895.520 ;
    END
  END io_out_as1802[17]
  PIN io_out_as1802[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 897.640 200.000 898.240 ;
    END
  END io_out_as1802[18]
  PIN io_out_as1802[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 900.360 200.000 900.960 ;
    END
  END io_out_as1802[19]
  PIN io_out_as1802[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 851.400 200.000 852.000 ;
    END
  END io_out_as1802[1]
  PIN io_out_as1802[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 903.080 200.000 903.680 ;
    END
  END io_out_as1802[20]
  PIN io_out_as1802[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 905.800 200.000 906.400 ;
    END
  END io_out_as1802[21]
  PIN io_out_as1802[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 908.520 200.000 909.120 ;
    END
  END io_out_as1802[22]
  PIN io_out_as1802[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 911.240 200.000 911.840 ;
    END
  END io_out_as1802[23]
  PIN io_out_as1802[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 913.960 200.000 914.560 ;
    END
  END io_out_as1802[24]
  PIN io_out_as1802[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 916.680 200.000 917.280 ;
    END
  END io_out_as1802[25]
  PIN io_out_as1802[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 919.400 200.000 920.000 ;
    END
  END io_out_as1802[26]
  PIN io_out_as1802[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 922.120 200.000 922.720 ;
    END
  END io_out_as1802[27]
  PIN io_out_as1802[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 924.840 200.000 925.440 ;
    END
  END io_out_as1802[28]
  PIN io_out_as1802[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 927.560 200.000 928.160 ;
    END
  END io_out_as1802[29]
  PIN io_out_as1802[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 854.120 200.000 854.720 ;
    END
  END io_out_as1802[2]
  PIN io_out_as1802[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 930.280 200.000 930.880 ;
    END
  END io_out_as1802[30]
  PIN io_out_as1802[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 933.000 200.000 933.600 ;
    END
  END io_out_as1802[31]
  PIN io_out_as1802[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 935.720 200.000 936.320 ;
    END
  END io_out_as1802[32]
  PIN io_out_as1802[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 938.440 200.000 939.040 ;
    END
  END io_out_as1802[33]
  PIN io_out_as1802[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 941.160 200.000 941.760 ;
    END
  END io_out_as1802[34]
  PIN io_out_as1802[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 943.880 200.000 944.480 ;
    END
  END io_out_as1802[35]
  PIN io_out_as1802[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 856.840 200.000 857.440 ;
    END
  END io_out_as1802[3]
  PIN io_out_as1802[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 859.560 200.000 860.160 ;
    END
  END io_out_as1802[4]
  PIN io_out_as1802[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 862.280 200.000 862.880 ;
    END
  END io_out_as1802[5]
  PIN io_out_as1802[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 865.000 200.000 865.600 ;
    END
  END io_out_as1802[6]
  PIN io_out_as1802[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 867.720 200.000 868.320 ;
    END
  END io_out_as1802[7]
  PIN io_out_as1802[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 870.440 200.000 871.040 ;
    END
  END io_out_as1802[8]
  PIN io_out_as1802[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 873.160 200.000 873.760 ;
    END
  END io_out_as1802[9]
  PIN io_out_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 750.760 200.000 751.360 ;
    END
  END io_out_scrapcpu[0]
  PIN io_out_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 777.960 200.000 778.560 ;
    END
  END io_out_scrapcpu[10]
  PIN io_out_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 780.680 200.000 781.280 ;
    END
  END io_out_scrapcpu[11]
  PIN io_out_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 783.400 200.000 784.000 ;
    END
  END io_out_scrapcpu[12]
  PIN io_out_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 786.120 200.000 786.720 ;
    END
  END io_out_scrapcpu[13]
  PIN io_out_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 788.840 200.000 789.440 ;
    END
  END io_out_scrapcpu[14]
  PIN io_out_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 791.560 200.000 792.160 ;
    END
  END io_out_scrapcpu[15]
  PIN io_out_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 794.280 200.000 794.880 ;
    END
  END io_out_scrapcpu[16]
  PIN io_out_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 797.000 200.000 797.600 ;
    END
  END io_out_scrapcpu[17]
  PIN io_out_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 799.720 200.000 800.320 ;
    END
  END io_out_scrapcpu[18]
  PIN io_out_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 802.440 200.000 803.040 ;
    END
  END io_out_scrapcpu[19]
  PIN io_out_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 753.480 200.000 754.080 ;
    END
  END io_out_scrapcpu[1]
  PIN io_out_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 805.160 200.000 805.760 ;
    END
  END io_out_scrapcpu[20]
  PIN io_out_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 807.880 200.000 808.480 ;
    END
  END io_out_scrapcpu[21]
  PIN io_out_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 810.600 200.000 811.200 ;
    END
  END io_out_scrapcpu[22]
  PIN io_out_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 813.320 200.000 813.920 ;
    END
  END io_out_scrapcpu[23]
  PIN io_out_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 816.040 200.000 816.640 ;
    END
  END io_out_scrapcpu[24]
  PIN io_out_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 818.760 200.000 819.360 ;
    END
  END io_out_scrapcpu[25]
  PIN io_out_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 821.480 200.000 822.080 ;
    END
  END io_out_scrapcpu[26]
  PIN io_out_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 824.200 200.000 824.800 ;
    END
  END io_out_scrapcpu[27]
  PIN io_out_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 826.920 200.000 827.520 ;
    END
  END io_out_scrapcpu[28]
  PIN io_out_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 829.640 200.000 830.240 ;
    END
  END io_out_scrapcpu[29]
  PIN io_out_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 756.200 200.000 756.800 ;
    END
  END io_out_scrapcpu[2]
  PIN io_out_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 832.360 200.000 832.960 ;
    END
  END io_out_scrapcpu[30]
  PIN io_out_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 835.080 200.000 835.680 ;
    END
  END io_out_scrapcpu[31]
  PIN io_out_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 837.800 200.000 838.400 ;
    END
  END io_out_scrapcpu[32]
  PIN io_out_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 840.520 200.000 841.120 ;
    END
  END io_out_scrapcpu[33]
  PIN io_out_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 843.240 200.000 843.840 ;
    END
  END io_out_scrapcpu[34]
  PIN io_out_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 845.960 200.000 846.560 ;
    END
  END io_out_scrapcpu[35]
  PIN io_out_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 758.920 200.000 759.520 ;
    END
  END io_out_scrapcpu[3]
  PIN io_out_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 761.640 200.000 762.240 ;
    END
  END io_out_scrapcpu[4]
  PIN io_out_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 764.360 200.000 764.960 ;
    END
  END io_out_scrapcpu[5]
  PIN io_out_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 767.080 200.000 767.680 ;
    END
  END io_out_scrapcpu[6]
  PIN io_out_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 769.800 200.000 770.400 ;
    END
  END io_out_scrapcpu[7]
  PIN io_out_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 772.520 200.000 773.120 ;
    END
  END io_out_scrapcpu[8]
  PIN io_out_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 775.240 200.000 775.840 ;
    END
  END io_out_scrapcpu[9]
  PIN io_out_vliw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 1096.000 19.690 1100.000 ;
    END
  END io_out_vliw[0]
  PIN io_out_vliw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 65.410 1096.000 65.690 1100.000 ;
    END
  END io_out_vliw[10]
  PIN io_out_vliw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 70.010 1096.000 70.290 1100.000 ;
    END
  END io_out_vliw[11]
  PIN io_out_vliw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 1096.000 74.890 1100.000 ;
    END
  END io_out_vliw[12]
  PIN io_out_vliw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 79.210 1096.000 79.490 1100.000 ;
    END
  END io_out_vliw[13]
  PIN io_out_vliw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 83.810 1096.000 84.090 1100.000 ;
    END
  END io_out_vliw[14]
  PIN io_out_vliw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 88.410 1096.000 88.690 1100.000 ;
    END
  END io_out_vliw[15]
  PIN io_out_vliw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 93.010 1096.000 93.290 1100.000 ;
    END
  END io_out_vliw[16]
  PIN io_out_vliw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 97.610 1096.000 97.890 1100.000 ;
    END
  END io_out_vliw[17]
  PIN io_out_vliw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 102.210 1096.000 102.490 1100.000 ;
    END
  END io_out_vliw[18]
  PIN io_out_vliw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 106.810 1096.000 107.090 1100.000 ;
    END
  END io_out_vliw[19]
  PIN io_out_vliw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 24.010 1096.000 24.290 1100.000 ;
    END
  END io_out_vliw[1]
  PIN io_out_vliw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 111.410 1096.000 111.690 1100.000 ;
    END
  END io_out_vliw[20]
  PIN io_out_vliw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 116.010 1096.000 116.290 1100.000 ;
    END
  END io_out_vliw[21]
  PIN io_out_vliw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 120.610 1096.000 120.890 1100.000 ;
    END
  END io_out_vliw[22]
  PIN io_out_vliw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 125.210 1096.000 125.490 1100.000 ;
    END
  END io_out_vliw[23]
  PIN io_out_vliw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 129.810 1096.000 130.090 1100.000 ;
    END
  END io_out_vliw[24]
  PIN io_out_vliw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 134.410 1096.000 134.690 1100.000 ;
    END
  END io_out_vliw[25]
  PIN io_out_vliw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 139.010 1096.000 139.290 1100.000 ;
    END
  END io_out_vliw[26]
  PIN io_out_vliw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 143.610 1096.000 143.890 1100.000 ;
    END
  END io_out_vliw[27]
  PIN io_out_vliw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 148.210 1096.000 148.490 1100.000 ;
    END
  END io_out_vliw[28]
  PIN io_out_vliw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 152.810 1096.000 153.090 1100.000 ;
    END
  END io_out_vliw[29]
  PIN io_out_vliw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 28.610 1096.000 28.890 1100.000 ;
    END
  END io_out_vliw[2]
  PIN io_out_vliw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 157.410 1096.000 157.690 1100.000 ;
    END
  END io_out_vliw[30]
  PIN io_out_vliw[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 162.010 1096.000 162.290 1100.000 ;
    END
  END io_out_vliw[31]
  PIN io_out_vliw[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 166.610 1096.000 166.890 1100.000 ;
    END
  END io_out_vliw[32]
  PIN io_out_vliw[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 171.210 1096.000 171.490 1100.000 ;
    END
  END io_out_vliw[33]
  PIN io_out_vliw[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 175.810 1096.000 176.090 1100.000 ;
    END
  END io_out_vliw[34]
  PIN io_out_vliw[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 180.410 1096.000 180.690 1100.000 ;
    END
  END io_out_vliw[35]
  PIN io_out_vliw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 33.210 1096.000 33.490 1100.000 ;
    END
  END io_out_vliw[3]
  PIN io_out_vliw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 37.810 1096.000 38.090 1100.000 ;
    END
  END io_out_vliw[4]
  PIN io_out_vliw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 42.410 1096.000 42.690 1100.000 ;
    END
  END io_out_vliw[5]
  PIN io_out_vliw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 47.010 1096.000 47.290 1100.000 ;
    END
  END io_out_vliw[6]
  PIN io_out_vliw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 1096.000 51.890 1100.000 ;
    END
  END io_out_vliw[7]
  PIN io_out_vliw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 56.210 1096.000 56.490 1100.000 ;
    END
  END io_out_vliw[8]
  PIN io_out_vliw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 60.810 1096.000 61.090 1100.000 ;
    END
  END io_out_vliw[9]
  PIN io_out_z80[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 552.200 200.000 552.800 ;
    END
  END io_out_z80[0]
  PIN io_out_z80[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 579.400 200.000 580.000 ;
    END
  END io_out_z80[10]
  PIN io_out_z80[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 582.120 200.000 582.720 ;
    END
  END io_out_z80[11]
  PIN io_out_z80[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 584.840 200.000 585.440 ;
    END
  END io_out_z80[12]
  PIN io_out_z80[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 587.560 200.000 588.160 ;
    END
  END io_out_z80[13]
  PIN io_out_z80[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 590.280 200.000 590.880 ;
    END
  END io_out_z80[14]
  PIN io_out_z80[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 593.000 200.000 593.600 ;
    END
  END io_out_z80[15]
  PIN io_out_z80[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 595.720 200.000 596.320 ;
    END
  END io_out_z80[16]
  PIN io_out_z80[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 598.440 200.000 599.040 ;
    END
  END io_out_z80[17]
  PIN io_out_z80[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 601.160 200.000 601.760 ;
    END
  END io_out_z80[18]
  PIN io_out_z80[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 603.880 200.000 604.480 ;
    END
  END io_out_z80[19]
  PIN io_out_z80[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 554.920 200.000 555.520 ;
    END
  END io_out_z80[1]
  PIN io_out_z80[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 606.600 200.000 607.200 ;
    END
  END io_out_z80[20]
  PIN io_out_z80[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 609.320 200.000 609.920 ;
    END
  END io_out_z80[21]
  PIN io_out_z80[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 612.040 200.000 612.640 ;
    END
  END io_out_z80[22]
  PIN io_out_z80[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 614.760 200.000 615.360 ;
    END
  END io_out_z80[23]
  PIN io_out_z80[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 617.480 200.000 618.080 ;
    END
  END io_out_z80[24]
  PIN io_out_z80[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 620.200 200.000 620.800 ;
    END
  END io_out_z80[25]
  PIN io_out_z80[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 622.920 200.000 623.520 ;
    END
  END io_out_z80[26]
  PIN io_out_z80[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 625.640 200.000 626.240 ;
    END
  END io_out_z80[27]
  PIN io_out_z80[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 628.360 200.000 628.960 ;
    END
  END io_out_z80[28]
  PIN io_out_z80[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 631.080 200.000 631.680 ;
    END
  END io_out_z80[29]
  PIN io_out_z80[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 557.640 200.000 558.240 ;
    END
  END io_out_z80[2]
  PIN io_out_z80[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 633.800 200.000 634.400 ;
    END
  END io_out_z80[30]
  PIN io_out_z80[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 636.520 200.000 637.120 ;
    END
  END io_out_z80[31]
  PIN io_out_z80[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 639.240 200.000 639.840 ;
    END
  END io_out_z80[32]
  PIN io_out_z80[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 641.960 200.000 642.560 ;
    END
  END io_out_z80[33]
  PIN io_out_z80[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 644.680 200.000 645.280 ;
    END
  END io_out_z80[34]
  PIN io_out_z80[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 647.400 200.000 648.000 ;
    END
  END io_out_z80[35]
  PIN io_out_z80[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 560.360 200.000 560.960 ;
    END
  END io_out_z80[3]
  PIN io_out_z80[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 563.080 200.000 563.680 ;
    END
  END io_out_z80[4]
  PIN io_out_z80[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 565.800 200.000 566.400 ;
    END
  END io_out_z80[5]
  PIN io_out_z80[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 568.520 200.000 569.120 ;
    END
  END io_out_z80[6]
  PIN io_out_z80[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 571.240 200.000 571.840 ;
    END
  END io_out_z80[7]
  PIN io_out_z80[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 573.960 200.000 574.560 ;
    END
  END io_out_z80[8]
  PIN io_out_z80[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 576.680 200.000 577.280 ;
    END
  END io_out_z80[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 443.400 200.000 444.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 470.600 200.000 471.200 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 473.320 200.000 473.920 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 476.040 200.000 476.640 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 478.760 200.000 479.360 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 481.480 200.000 482.080 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 484.200 200.000 484.800 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 486.920 200.000 487.520 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 489.640 200.000 490.240 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 492.360 200.000 492.960 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 495.080 200.000 495.680 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 446.120 200.000 446.720 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 497.800 200.000 498.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 500.520 200.000 501.120 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 503.240 200.000 503.840 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 505.960 200.000 506.560 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 508.680 200.000 509.280 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 511.400 200.000 512.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 514.120 200.000 514.720 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 516.840 200.000 517.440 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 519.560 200.000 520.160 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 522.280 200.000 522.880 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 448.840 200.000 449.440 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 525.000 200.000 525.600 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 527.720 200.000 528.320 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 530.440 200.000 531.040 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 533.160 200.000 533.760 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 535.880 200.000 536.480 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 538.600 200.000 539.200 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 541.320 200.000 541.920 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 544.040 200.000 544.640 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 546.760 200.000 547.360 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 549.480 200.000 550.080 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 451.560 200.000 452.160 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 454.280 200.000 454.880 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 457.000 200.000 457.600 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 459.720 200.000 460.320 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 462.440 200.000 463.040 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 465.160 200.000 465.760 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 467.880 200.000 468.480 ;
    END
  END la_data_out[9]
  PIN rst_6502
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END rst_6502
  PIN rst_as1802
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 189.610 1096.000 189.890 1100.000 ;
    END
  END rst_as1802
  PIN rst_scrapcpu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 185.010 1096.000 185.290 1100.000 ;
    END
  END rst_scrapcpu
  PIN rst_vliw
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 14.810 1096.000 15.090 1100.000 ;
    END
  END rst_vliw
  PIN rst_z80
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 650.120 200.000 650.720 ;
    END
  END rst_z80
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1088.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 0.000 64.310 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 0.000 177.930 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.120 4.000 378.720 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.760 4.000 411.360 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 443.400 4.000 444.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 356.360 200.000 356.960 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 383.560 200.000 384.160 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 386.280 200.000 386.880 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 389.000 200.000 389.600 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 391.720 200.000 392.320 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 394.440 200.000 395.040 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 397.160 200.000 397.760 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 399.880 200.000 400.480 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 402.600 200.000 403.200 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 405.320 200.000 405.920 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 408.040 200.000 408.640 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 359.080 200.000 359.680 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 410.760 200.000 411.360 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 413.480 200.000 414.080 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 416.200 200.000 416.800 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 418.920 200.000 419.520 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 421.640 200.000 422.240 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 424.360 200.000 424.960 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 427.080 200.000 427.680 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 429.800 200.000 430.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 432.520 200.000 433.120 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 435.240 200.000 435.840 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 361.800 200.000 362.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 437.960 200.000 438.560 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 440.680 200.000 441.280 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 364.520 200.000 365.120 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 367.240 200.000 367.840 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 369.960 200.000 370.560 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 372.680 200.000 373.280 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 375.400 200.000 376.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 378.120 200.000 378.720 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 380.840 200.000 381.440 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 1088.085 ;
      LAYER met1 ;
        RECT 0.530 10.640 199.570 1088.240 ;
      LAYER met2 ;
        RECT 0.550 1095.720 9.930 1096.570 ;
        RECT 10.770 1095.720 14.530 1096.570 ;
        RECT 15.370 1095.720 19.130 1096.570 ;
        RECT 19.970 1095.720 23.730 1096.570 ;
        RECT 24.570 1095.720 28.330 1096.570 ;
        RECT 29.170 1095.720 32.930 1096.570 ;
        RECT 33.770 1095.720 37.530 1096.570 ;
        RECT 38.370 1095.720 42.130 1096.570 ;
        RECT 42.970 1095.720 46.730 1096.570 ;
        RECT 47.570 1095.720 51.330 1096.570 ;
        RECT 52.170 1095.720 55.930 1096.570 ;
        RECT 56.770 1095.720 60.530 1096.570 ;
        RECT 61.370 1095.720 65.130 1096.570 ;
        RECT 65.970 1095.720 69.730 1096.570 ;
        RECT 70.570 1095.720 74.330 1096.570 ;
        RECT 75.170 1095.720 78.930 1096.570 ;
        RECT 79.770 1095.720 83.530 1096.570 ;
        RECT 84.370 1095.720 88.130 1096.570 ;
        RECT 88.970 1095.720 92.730 1096.570 ;
        RECT 93.570 1095.720 97.330 1096.570 ;
        RECT 98.170 1095.720 101.930 1096.570 ;
        RECT 102.770 1095.720 106.530 1096.570 ;
        RECT 107.370 1095.720 111.130 1096.570 ;
        RECT 111.970 1095.720 115.730 1096.570 ;
        RECT 116.570 1095.720 120.330 1096.570 ;
        RECT 121.170 1095.720 124.930 1096.570 ;
        RECT 125.770 1095.720 129.530 1096.570 ;
        RECT 130.370 1095.720 134.130 1096.570 ;
        RECT 134.970 1095.720 138.730 1096.570 ;
        RECT 139.570 1095.720 143.330 1096.570 ;
        RECT 144.170 1095.720 147.930 1096.570 ;
        RECT 148.770 1095.720 152.530 1096.570 ;
        RECT 153.370 1095.720 157.130 1096.570 ;
        RECT 157.970 1095.720 161.730 1096.570 ;
        RECT 162.570 1095.720 166.330 1096.570 ;
        RECT 167.170 1095.720 170.930 1096.570 ;
        RECT 171.770 1095.720 175.530 1096.570 ;
        RECT 176.370 1095.720 180.130 1096.570 ;
        RECT 180.970 1095.720 184.730 1096.570 ;
        RECT 185.570 1095.720 189.330 1096.570 ;
        RECT 190.170 1095.720 199.940 1096.570 ;
        RECT 0.550 4.280 199.940 1095.720 ;
        RECT 0.550 3.670 3.950 4.280 ;
        RECT 4.790 3.670 9.930 4.280 ;
        RECT 10.770 3.670 15.910 4.280 ;
        RECT 16.750 3.670 21.890 4.280 ;
        RECT 22.730 3.670 27.870 4.280 ;
        RECT 28.710 3.670 33.850 4.280 ;
        RECT 34.690 3.670 39.830 4.280 ;
        RECT 40.670 3.670 45.810 4.280 ;
        RECT 46.650 3.670 51.790 4.280 ;
        RECT 52.630 3.670 57.770 4.280 ;
        RECT 58.610 3.670 63.750 4.280 ;
        RECT 64.590 3.670 69.730 4.280 ;
        RECT 70.570 3.670 75.710 4.280 ;
        RECT 76.550 3.670 81.690 4.280 ;
        RECT 82.530 3.670 87.670 4.280 ;
        RECT 88.510 3.670 93.650 4.280 ;
        RECT 94.490 3.670 99.630 4.280 ;
        RECT 100.470 3.670 105.610 4.280 ;
        RECT 106.450 3.670 111.590 4.280 ;
        RECT 112.430 3.670 117.570 4.280 ;
        RECT 118.410 3.670 123.550 4.280 ;
        RECT 124.390 3.670 129.530 4.280 ;
        RECT 130.370 3.670 135.510 4.280 ;
        RECT 136.350 3.670 141.490 4.280 ;
        RECT 142.330 3.670 147.470 4.280 ;
        RECT 148.310 3.670 153.450 4.280 ;
        RECT 154.290 3.670 159.430 4.280 ;
        RECT 160.270 3.670 165.410 4.280 ;
        RECT 166.250 3.670 171.390 4.280 ;
        RECT 172.230 3.670 177.370 4.280 ;
        RECT 178.210 3.670 183.350 4.280 ;
        RECT 184.190 3.670 189.330 4.280 ;
        RECT 190.170 3.670 195.310 4.280 ;
        RECT 196.150 3.670 199.940 4.280 ;
      LAYER met3 ;
        RECT 0.525 1037.360 199.575 1088.165 ;
        RECT 4.400 1035.960 199.575 1037.360 ;
        RECT 0.525 1031.920 199.575 1035.960 ;
        RECT 4.400 1030.520 199.575 1031.920 ;
        RECT 0.525 1026.480 199.575 1030.520 ;
        RECT 4.400 1025.080 199.575 1026.480 ;
        RECT 0.525 1021.040 199.575 1025.080 ;
        RECT 4.400 1019.640 199.575 1021.040 ;
        RECT 0.525 1015.600 199.575 1019.640 ;
        RECT 4.400 1014.200 199.575 1015.600 ;
        RECT 0.525 1010.160 199.575 1014.200 ;
        RECT 4.400 1008.760 199.575 1010.160 ;
        RECT 0.525 1004.720 199.575 1008.760 ;
        RECT 4.400 1003.320 199.575 1004.720 ;
        RECT 0.525 999.280 199.575 1003.320 ;
        RECT 4.400 997.880 199.575 999.280 ;
        RECT 0.525 993.840 199.575 997.880 ;
        RECT 4.400 992.440 199.575 993.840 ;
        RECT 0.525 988.400 199.575 992.440 ;
        RECT 4.400 987.000 199.575 988.400 ;
        RECT 0.525 982.960 199.575 987.000 ;
        RECT 4.400 981.560 199.575 982.960 ;
        RECT 0.525 977.520 199.575 981.560 ;
        RECT 4.400 976.120 199.575 977.520 ;
        RECT 0.525 972.080 199.575 976.120 ;
        RECT 4.400 970.680 199.575 972.080 ;
        RECT 0.525 966.640 199.575 970.680 ;
        RECT 4.400 965.240 199.575 966.640 ;
        RECT 0.525 961.200 199.575 965.240 ;
        RECT 4.400 959.800 199.575 961.200 ;
        RECT 0.525 955.760 199.575 959.800 ;
        RECT 4.400 954.360 199.575 955.760 ;
        RECT 0.525 950.320 199.575 954.360 ;
        RECT 4.400 948.920 199.575 950.320 ;
        RECT 0.525 947.600 199.575 948.920 ;
        RECT 0.525 946.200 195.600 947.600 ;
        RECT 0.525 944.880 199.575 946.200 ;
        RECT 4.400 943.480 195.600 944.880 ;
        RECT 0.525 942.160 199.575 943.480 ;
        RECT 0.525 940.760 195.600 942.160 ;
        RECT 0.525 939.440 199.575 940.760 ;
        RECT 4.400 938.040 195.600 939.440 ;
        RECT 0.525 936.720 199.575 938.040 ;
        RECT 0.525 935.320 195.600 936.720 ;
        RECT 0.525 934.000 199.575 935.320 ;
        RECT 4.400 932.600 195.600 934.000 ;
        RECT 0.525 931.280 199.575 932.600 ;
        RECT 0.525 929.880 195.600 931.280 ;
        RECT 0.525 928.560 199.575 929.880 ;
        RECT 4.400 927.160 195.600 928.560 ;
        RECT 0.525 925.840 199.575 927.160 ;
        RECT 0.525 924.440 195.600 925.840 ;
        RECT 0.525 923.120 199.575 924.440 ;
        RECT 4.400 921.720 195.600 923.120 ;
        RECT 0.525 920.400 199.575 921.720 ;
        RECT 0.525 919.000 195.600 920.400 ;
        RECT 0.525 917.680 199.575 919.000 ;
        RECT 4.400 916.280 195.600 917.680 ;
        RECT 0.525 914.960 199.575 916.280 ;
        RECT 0.525 913.560 195.600 914.960 ;
        RECT 0.525 912.240 199.575 913.560 ;
        RECT 4.400 910.840 195.600 912.240 ;
        RECT 0.525 909.520 199.575 910.840 ;
        RECT 0.525 908.120 195.600 909.520 ;
        RECT 0.525 906.800 199.575 908.120 ;
        RECT 4.400 905.400 195.600 906.800 ;
        RECT 0.525 904.080 199.575 905.400 ;
        RECT 0.525 902.680 195.600 904.080 ;
        RECT 0.525 901.360 199.575 902.680 ;
        RECT 4.400 899.960 195.600 901.360 ;
        RECT 0.525 898.640 199.575 899.960 ;
        RECT 0.525 897.240 195.600 898.640 ;
        RECT 0.525 895.920 199.575 897.240 ;
        RECT 4.400 894.520 195.600 895.920 ;
        RECT 0.525 893.200 199.575 894.520 ;
        RECT 0.525 891.800 195.600 893.200 ;
        RECT 0.525 890.480 199.575 891.800 ;
        RECT 4.400 889.080 195.600 890.480 ;
        RECT 0.525 887.760 199.575 889.080 ;
        RECT 0.525 886.360 195.600 887.760 ;
        RECT 0.525 885.040 199.575 886.360 ;
        RECT 4.400 883.640 195.600 885.040 ;
        RECT 0.525 882.320 199.575 883.640 ;
        RECT 0.525 880.920 195.600 882.320 ;
        RECT 0.525 879.600 199.575 880.920 ;
        RECT 4.400 878.200 195.600 879.600 ;
        RECT 0.525 876.880 199.575 878.200 ;
        RECT 0.525 875.480 195.600 876.880 ;
        RECT 0.525 874.160 199.575 875.480 ;
        RECT 4.400 872.760 195.600 874.160 ;
        RECT 0.525 871.440 199.575 872.760 ;
        RECT 0.525 870.040 195.600 871.440 ;
        RECT 0.525 868.720 199.575 870.040 ;
        RECT 4.400 867.320 195.600 868.720 ;
        RECT 0.525 866.000 199.575 867.320 ;
        RECT 0.525 864.600 195.600 866.000 ;
        RECT 0.525 863.280 199.575 864.600 ;
        RECT 4.400 861.880 195.600 863.280 ;
        RECT 0.525 860.560 199.575 861.880 ;
        RECT 0.525 859.160 195.600 860.560 ;
        RECT 0.525 857.840 199.575 859.160 ;
        RECT 4.400 856.440 195.600 857.840 ;
        RECT 0.525 855.120 199.575 856.440 ;
        RECT 0.525 853.720 195.600 855.120 ;
        RECT 0.525 852.400 199.575 853.720 ;
        RECT 4.400 851.000 195.600 852.400 ;
        RECT 0.525 849.680 199.575 851.000 ;
        RECT 0.525 848.280 195.600 849.680 ;
        RECT 0.525 846.960 199.575 848.280 ;
        RECT 4.400 845.560 195.600 846.960 ;
        RECT 0.525 844.240 199.575 845.560 ;
        RECT 0.525 842.840 195.600 844.240 ;
        RECT 0.525 841.520 199.575 842.840 ;
        RECT 4.400 840.120 195.600 841.520 ;
        RECT 0.525 838.800 199.575 840.120 ;
        RECT 0.525 837.400 195.600 838.800 ;
        RECT 0.525 836.080 199.575 837.400 ;
        RECT 4.400 834.680 195.600 836.080 ;
        RECT 0.525 833.360 199.575 834.680 ;
        RECT 0.525 831.960 195.600 833.360 ;
        RECT 0.525 830.640 199.575 831.960 ;
        RECT 4.400 829.240 195.600 830.640 ;
        RECT 0.525 827.920 199.575 829.240 ;
        RECT 0.525 826.520 195.600 827.920 ;
        RECT 0.525 825.200 199.575 826.520 ;
        RECT 4.400 823.800 195.600 825.200 ;
        RECT 0.525 822.480 199.575 823.800 ;
        RECT 0.525 821.080 195.600 822.480 ;
        RECT 0.525 819.760 199.575 821.080 ;
        RECT 4.400 818.360 195.600 819.760 ;
        RECT 0.525 817.040 199.575 818.360 ;
        RECT 0.525 815.640 195.600 817.040 ;
        RECT 0.525 814.320 199.575 815.640 ;
        RECT 4.400 812.920 195.600 814.320 ;
        RECT 0.525 811.600 199.575 812.920 ;
        RECT 0.525 810.200 195.600 811.600 ;
        RECT 0.525 808.880 199.575 810.200 ;
        RECT 4.400 807.480 195.600 808.880 ;
        RECT 0.525 806.160 199.575 807.480 ;
        RECT 0.525 804.760 195.600 806.160 ;
        RECT 0.525 803.440 199.575 804.760 ;
        RECT 4.400 802.040 195.600 803.440 ;
        RECT 0.525 800.720 199.575 802.040 ;
        RECT 0.525 799.320 195.600 800.720 ;
        RECT 0.525 798.000 199.575 799.320 ;
        RECT 4.400 796.600 195.600 798.000 ;
        RECT 0.525 795.280 199.575 796.600 ;
        RECT 0.525 793.880 195.600 795.280 ;
        RECT 0.525 792.560 199.575 793.880 ;
        RECT 4.400 791.160 195.600 792.560 ;
        RECT 0.525 789.840 199.575 791.160 ;
        RECT 0.525 788.440 195.600 789.840 ;
        RECT 0.525 787.120 199.575 788.440 ;
        RECT 4.400 785.720 195.600 787.120 ;
        RECT 0.525 784.400 199.575 785.720 ;
        RECT 0.525 783.000 195.600 784.400 ;
        RECT 0.525 781.680 199.575 783.000 ;
        RECT 4.400 780.280 195.600 781.680 ;
        RECT 0.525 778.960 199.575 780.280 ;
        RECT 0.525 777.560 195.600 778.960 ;
        RECT 0.525 776.240 199.575 777.560 ;
        RECT 4.400 774.840 195.600 776.240 ;
        RECT 0.525 773.520 199.575 774.840 ;
        RECT 0.525 772.120 195.600 773.520 ;
        RECT 0.525 770.800 199.575 772.120 ;
        RECT 4.400 769.400 195.600 770.800 ;
        RECT 0.525 768.080 199.575 769.400 ;
        RECT 0.525 766.680 195.600 768.080 ;
        RECT 0.525 765.360 199.575 766.680 ;
        RECT 4.400 763.960 195.600 765.360 ;
        RECT 0.525 762.640 199.575 763.960 ;
        RECT 0.525 761.240 195.600 762.640 ;
        RECT 0.525 759.920 199.575 761.240 ;
        RECT 4.400 758.520 195.600 759.920 ;
        RECT 0.525 757.200 199.575 758.520 ;
        RECT 0.525 755.800 195.600 757.200 ;
        RECT 0.525 754.480 199.575 755.800 ;
        RECT 4.400 753.080 195.600 754.480 ;
        RECT 0.525 751.760 199.575 753.080 ;
        RECT 0.525 750.360 195.600 751.760 ;
        RECT 0.525 749.040 199.575 750.360 ;
        RECT 4.400 747.640 195.600 749.040 ;
        RECT 0.525 746.320 199.575 747.640 ;
        RECT 0.525 744.920 195.600 746.320 ;
        RECT 0.525 743.600 199.575 744.920 ;
        RECT 4.400 742.200 195.600 743.600 ;
        RECT 0.525 740.880 199.575 742.200 ;
        RECT 0.525 739.480 195.600 740.880 ;
        RECT 0.525 738.160 199.575 739.480 ;
        RECT 4.400 736.760 195.600 738.160 ;
        RECT 0.525 735.440 199.575 736.760 ;
        RECT 0.525 734.040 195.600 735.440 ;
        RECT 0.525 732.720 199.575 734.040 ;
        RECT 4.400 731.320 195.600 732.720 ;
        RECT 0.525 730.000 199.575 731.320 ;
        RECT 0.525 728.600 195.600 730.000 ;
        RECT 0.525 727.280 199.575 728.600 ;
        RECT 4.400 725.880 195.600 727.280 ;
        RECT 0.525 724.560 199.575 725.880 ;
        RECT 0.525 723.160 195.600 724.560 ;
        RECT 0.525 721.840 199.575 723.160 ;
        RECT 4.400 720.440 195.600 721.840 ;
        RECT 0.525 719.120 199.575 720.440 ;
        RECT 0.525 717.720 195.600 719.120 ;
        RECT 0.525 716.400 199.575 717.720 ;
        RECT 4.400 715.000 195.600 716.400 ;
        RECT 0.525 713.680 199.575 715.000 ;
        RECT 0.525 712.280 195.600 713.680 ;
        RECT 0.525 710.960 199.575 712.280 ;
        RECT 4.400 709.560 195.600 710.960 ;
        RECT 0.525 708.240 199.575 709.560 ;
        RECT 0.525 706.840 195.600 708.240 ;
        RECT 0.525 705.520 199.575 706.840 ;
        RECT 4.400 704.120 195.600 705.520 ;
        RECT 0.525 702.800 199.575 704.120 ;
        RECT 0.525 701.400 195.600 702.800 ;
        RECT 0.525 700.080 199.575 701.400 ;
        RECT 4.400 698.680 195.600 700.080 ;
        RECT 0.525 697.360 199.575 698.680 ;
        RECT 0.525 695.960 195.600 697.360 ;
        RECT 0.525 694.640 199.575 695.960 ;
        RECT 4.400 693.240 195.600 694.640 ;
        RECT 0.525 691.920 199.575 693.240 ;
        RECT 0.525 690.520 195.600 691.920 ;
        RECT 0.525 689.200 199.575 690.520 ;
        RECT 4.400 687.800 195.600 689.200 ;
        RECT 0.525 686.480 199.575 687.800 ;
        RECT 0.525 685.080 195.600 686.480 ;
        RECT 0.525 683.760 199.575 685.080 ;
        RECT 4.400 682.360 195.600 683.760 ;
        RECT 0.525 681.040 199.575 682.360 ;
        RECT 0.525 679.640 195.600 681.040 ;
        RECT 0.525 678.320 199.575 679.640 ;
        RECT 4.400 676.920 195.600 678.320 ;
        RECT 0.525 675.600 199.575 676.920 ;
        RECT 0.525 674.200 195.600 675.600 ;
        RECT 0.525 672.880 199.575 674.200 ;
        RECT 4.400 671.480 195.600 672.880 ;
        RECT 0.525 670.160 199.575 671.480 ;
        RECT 0.525 668.760 195.600 670.160 ;
        RECT 0.525 667.440 199.575 668.760 ;
        RECT 4.400 666.040 195.600 667.440 ;
        RECT 0.525 664.720 199.575 666.040 ;
        RECT 0.525 663.320 195.600 664.720 ;
        RECT 0.525 662.000 199.575 663.320 ;
        RECT 4.400 660.600 195.600 662.000 ;
        RECT 0.525 659.280 199.575 660.600 ;
        RECT 0.525 657.880 195.600 659.280 ;
        RECT 0.525 656.560 199.575 657.880 ;
        RECT 4.400 655.160 195.600 656.560 ;
        RECT 0.525 653.840 199.575 655.160 ;
        RECT 0.525 652.440 195.600 653.840 ;
        RECT 0.525 651.120 199.575 652.440 ;
        RECT 4.400 649.720 195.600 651.120 ;
        RECT 0.525 648.400 199.575 649.720 ;
        RECT 0.525 647.000 195.600 648.400 ;
        RECT 0.525 645.680 199.575 647.000 ;
        RECT 4.400 644.280 195.600 645.680 ;
        RECT 0.525 642.960 199.575 644.280 ;
        RECT 0.525 641.560 195.600 642.960 ;
        RECT 0.525 640.240 199.575 641.560 ;
        RECT 4.400 638.840 195.600 640.240 ;
        RECT 0.525 637.520 199.575 638.840 ;
        RECT 0.525 636.120 195.600 637.520 ;
        RECT 0.525 634.800 199.575 636.120 ;
        RECT 4.400 633.400 195.600 634.800 ;
        RECT 0.525 632.080 199.575 633.400 ;
        RECT 0.525 630.680 195.600 632.080 ;
        RECT 0.525 629.360 199.575 630.680 ;
        RECT 4.400 627.960 195.600 629.360 ;
        RECT 0.525 626.640 199.575 627.960 ;
        RECT 0.525 625.240 195.600 626.640 ;
        RECT 0.525 623.920 199.575 625.240 ;
        RECT 4.400 622.520 195.600 623.920 ;
        RECT 0.525 621.200 199.575 622.520 ;
        RECT 0.525 619.800 195.600 621.200 ;
        RECT 0.525 618.480 199.575 619.800 ;
        RECT 4.400 617.080 195.600 618.480 ;
        RECT 0.525 615.760 199.575 617.080 ;
        RECT 0.525 614.360 195.600 615.760 ;
        RECT 0.525 613.040 199.575 614.360 ;
        RECT 4.400 611.640 195.600 613.040 ;
        RECT 0.525 610.320 199.575 611.640 ;
        RECT 0.525 608.920 195.600 610.320 ;
        RECT 0.525 607.600 199.575 608.920 ;
        RECT 4.400 606.200 195.600 607.600 ;
        RECT 0.525 604.880 199.575 606.200 ;
        RECT 0.525 603.480 195.600 604.880 ;
        RECT 0.525 602.160 199.575 603.480 ;
        RECT 4.400 600.760 195.600 602.160 ;
        RECT 0.525 599.440 199.575 600.760 ;
        RECT 0.525 598.040 195.600 599.440 ;
        RECT 0.525 596.720 199.575 598.040 ;
        RECT 4.400 595.320 195.600 596.720 ;
        RECT 0.525 594.000 199.575 595.320 ;
        RECT 0.525 592.600 195.600 594.000 ;
        RECT 0.525 591.280 199.575 592.600 ;
        RECT 4.400 589.880 195.600 591.280 ;
        RECT 0.525 588.560 199.575 589.880 ;
        RECT 0.525 587.160 195.600 588.560 ;
        RECT 0.525 585.840 199.575 587.160 ;
        RECT 4.400 584.440 195.600 585.840 ;
        RECT 0.525 583.120 199.575 584.440 ;
        RECT 0.525 581.720 195.600 583.120 ;
        RECT 0.525 580.400 199.575 581.720 ;
        RECT 4.400 579.000 195.600 580.400 ;
        RECT 0.525 577.680 199.575 579.000 ;
        RECT 0.525 576.280 195.600 577.680 ;
        RECT 0.525 574.960 199.575 576.280 ;
        RECT 4.400 573.560 195.600 574.960 ;
        RECT 0.525 572.240 199.575 573.560 ;
        RECT 0.525 570.840 195.600 572.240 ;
        RECT 0.525 569.520 199.575 570.840 ;
        RECT 4.400 568.120 195.600 569.520 ;
        RECT 0.525 566.800 199.575 568.120 ;
        RECT 0.525 565.400 195.600 566.800 ;
        RECT 0.525 564.080 199.575 565.400 ;
        RECT 4.400 562.680 195.600 564.080 ;
        RECT 0.525 561.360 199.575 562.680 ;
        RECT 0.525 559.960 195.600 561.360 ;
        RECT 0.525 558.640 199.575 559.960 ;
        RECT 4.400 557.240 195.600 558.640 ;
        RECT 0.525 555.920 199.575 557.240 ;
        RECT 0.525 554.520 195.600 555.920 ;
        RECT 0.525 553.200 199.575 554.520 ;
        RECT 4.400 551.800 195.600 553.200 ;
        RECT 0.525 550.480 199.575 551.800 ;
        RECT 0.525 549.080 195.600 550.480 ;
        RECT 0.525 547.760 199.575 549.080 ;
        RECT 4.400 546.360 195.600 547.760 ;
        RECT 0.525 545.040 199.575 546.360 ;
        RECT 0.525 543.640 195.600 545.040 ;
        RECT 0.525 542.320 199.575 543.640 ;
        RECT 4.400 540.920 195.600 542.320 ;
        RECT 0.525 539.600 199.575 540.920 ;
        RECT 0.525 538.200 195.600 539.600 ;
        RECT 0.525 536.880 199.575 538.200 ;
        RECT 4.400 535.480 195.600 536.880 ;
        RECT 0.525 534.160 199.575 535.480 ;
        RECT 0.525 532.760 195.600 534.160 ;
        RECT 0.525 531.440 199.575 532.760 ;
        RECT 4.400 530.040 195.600 531.440 ;
        RECT 0.525 528.720 199.575 530.040 ;
        RECT 0.525 527.320 195.600 528.720 ;
        RECT 0.525 526.000 199.575 527.320 ;
        RECT 4.400 524.600 195.600 526.000 ;
        RECT 0.525 523.280 199.575 524.600 ;
        RECT 0.525 521.880 195.600 523.280 ;
        RECT 0.525 520.560 199.575 521.880 ;
        RECT 4.400 519.160 195.600 520.560 ;
        RECT 0.525 517.840 199.575 519.160 ;
        RECT 0.525 516.440 195.600 517.840 ;
        RECT 0.525 515.120 199.575 516.440 ;
        RECT 4.400 513.720 195.600 515.120 ;
        RECT 0.525 512.400 199.575 513.720 ;
        RECT 0.525 511.000 195.600 512.400 ;
        RECT 0.525 509.680 199.575 511.000 ;
        RECT 4.400 508.280 195.600 509.680 ;
        RECT 0.525 506.960 199.575 508.280 ;
        RECT 0.525 505.560 195.600 506.960 ;
        RECT 0.525 504.240 199.575 505.560 ;
        RECT 4.400 502.840 195.600 504.240 ;
        RECT 0.525 501.520 199.575 502.840 ;
        RECT 0.525 500.120 195.600 501.520 ;
        RECT 0.525 498.800 199.575 500.120 ;
        RECT 4.400 497.400 195.600 498.800 ;
        RECT 0.525 496.080 199.575 497.400 ;
        RECT 0.525 494.680 195.600 496.080 ;
        RECT 0.525 493.360 199.575 494.680 ;
        RECT 4.400 491.960 195.600 493.360 ;
        RECT 0.525 490.640 199.575 491.960 ;
        RECT 0.525 489.240 195.600 490.640 ;
        RECT 0.525 487.920 199.575 489.240 ;
        RECT 4.400 486.520 195.600 487.920 ;
        RECT 0.525 485.200 199.575 486.520 ;
        RECT 0.525 483.800 195.600 485.200 ;
        RECT 0.525 482.480 199.575 483.800 ;
        RECT 4.400 481.080 195.600 482.480 ;
        RECT 0.525 479.760 199.575 481.080 ;
        RECT 0.525 478.360 195.600 479.760 ;
        RECT 0.525 477.040 199.575 478.360 ;
        RECT 4.400 475.640 195.600 477.040 ;
        RECT 0.525 474.320 199.575 475.640 ;
        RECT 0.525 472.920 195.600 474.320 ;
        RECT 0.525 471.600 199.575 472.920 ;
        RECT 4.400 470.200 195.600 471.600 ;
        RECT 0.525 468.880 199.575 470.200 ;
        RECT 0.525 467.480 195.600 468.880 ;
        RECT 0.525 466.160 199.575 467.480 ;
        RECT 4.400 464.760 195.600 466.160 ;
        RECT 0.525 463.440 199.575 464.760 ;
        RECT 0.525 462.040 195.600 463.440 ;
        RECT 0.525 460.720 199.575 462.040 ;
        RECT 4.400 459.320 195.600 460.720 ;
        RECT 0.525 458.000 199.575 459.320 ;
        RECT 0.525 456.600 195.600 458.000 ;
        RECT 0.525 455.280 199.575 456.600 ;
        RECT 4.400 453.880 195.600 455.280 ;
        RECT 0.525 452.560 199.575 453.880 ;
        RECT 0.525 451.160 195.600 452.560 ;
        RECT 0.525 449.840 199.575 451.160 ;
        RECT 4.400 448.440 195.600 449.840 ;
        RECT 0.525 447.120 199.575 448.440 ;
        RECT 0.525 445.720 195.600 447.120 ;
        RECT 0.525 444.400 199.575 445.720 ;
        RECT 4.400 443.000 195.600 444.400 ;
        RECT 0.525 441.680 199.575 443.000 ;
        RECT 0.525 440.280 195.600 441.680 ;
        RECT 0.525 438.960 199.575 440.280 ;
        RECT 4.400 437.560 195.600 438.960 ;
        RECT 0.525 436.240 199.575 437.560 ;
        RECT 0.525 434.840 195.600 436.240 ;
        RECT 0.525 433.520 199.575 434.840 ;
        RECT 4.400 432.120 195.600 433.520 ;
        RECT 0.525 430.800 199.575 432.120 ;
        RECT 0.525 429.400 195.600 430.800 ;
        RECT 0.525 428.080 199.575 429.400 ;
        RECT 4.400 426.680 195.600 428.080 ;
        RECT 0.525 425.360 199.575 426.680 ;
        RECT 0.525 423.960 195.600 425.360 ;
        RECT 0.525 422.640 199.575 423.960 ;
        RECT 4.400 421.240 195.600 422.640 ;
        RECT 0.525 419.920 199.575 421.240 ;
        RECT 0.525 418.520 195.600 419.920 ;
        RECT 0.525 417.200 199.575 418.520 ;
        RECT 4.400 415.800 195.600 417.200 ;
        RECT 0.525 414.480 199.575 415.800 ;
        RECT 0.525 413.080 195.600 414.480 ;
        RECT 0.525 411.760 199.575 413.080 ;
        RECT 4.400 410.360 195.600 411.760 ;
        RECT 0.525 409.040 199.575 410.360 ;
        RECT 0.525 407.640 195.600 409.040 ;
        RECT 0.525 406.320 199.575 407.640 ;
        RECT 4.400 404.920 195.600 406.320 ;
        RECT 0.525 403.600 199.575 404.920 ;
        RECT 0.525 402.200 195.600 403.600 ;
        RECT 0.525 400.880 199.575 402.200 ;
        RECT 4.400 399.480 195.600 400.880 ;
        RECT 0.525 398.160 199.575 399.480 ;
        RECT 0.525 396.760 195.600 398.160 ;
        RECT 0.525 395.440 199.575 396.760 ;
        RECT 4.400 394.040 195.600 395.440 ;
        RECT 0.525 392.720 199.575 394.040 ;
        RECT 0.525 391.320 195.600 392.720 ;
        RECT 0.525 390.000 199.575 391.320 ;
        RECT 4.400 388.600 195.600 390.000 ;
        RECT 0.525 387.280 199.575 388.600 ;
        RECT 0.525 385.880 195.600 387.280 ;
        RECT 0.525 384.560 199.575 385.880 ;
        RECT 4.400 383.160 195.600 384.560 ;
        RECT 0.525 381.840 199.575 383.160 ;
        RECT 0.525 380.440 195.600 381.840 ;
        RECT 0.525 379.120 199.575 380.440 ;
        RECT 4.400 377.720 195.600 379.120 ;
        RECT 0.525 376.400 199.575 377.720 ;
        RECT 0.525 375.000 195.600 376.400 ;
        RECT 0.525 373.680 199.575 375.000 ;
        RECT 4.400 372.280 195.600 373.680 ;
        RECT 0.525 370.960 199.575 372.280 ;
        RECT 0.525 369.560 195.600 370.960 ;
        RECT 0.525 368.240 199.575 369.560 ;
        RECT 4.400 366.840 195.600 368.240 ;
        RECT 0.525 365.520 199.575 366.840 ;
        RECT 0.525 364.120 195.600 365.520 ;
        RECT 0.525 362.800 199.575 364.120 ;
        RECT 4.400 361.400 195.600 362.800 ;
        RECT 0.525 360.080 199.575 361.400 ;
        RECT 0.525 358.680 195.600 360.080 ;
        RECT 0.525 357.360 199.575 358.680 ;
        RECT 4.400 355.960 195.600 357.360 ;
        RECT 0.525 354.640 199.575 355.960 ;
        RECT 0.525 353.240 195.600 354.640 ;
        RECT 0.525 351.920 199.575 353.240 ;
        RECT 4.400 350.520 195.600 351.920 ;
        RECT 0.525 349.200 199.575 350.520 ;
        RECT 0.525 347.800 195.600 349.200 ;
        RECT 0.525 346.480 199.575 347.800 ;
        RECT 4.400 345.080 195.600 346.480 ;
        RECT 0.525 343.760 199.575 345.080 ;
        RECT 0.525 342.360 195.600 343.760 ;
        RECT 0.525 341.040 199.575 342.360 ;
        RECT 4.400 339.640 195.600 341.040 ;
        RECT 0.525 338.320 199.575 339.640 ;
        RECT 0.525 336.920 195.600 338.320 ;
        RECT 0.525 335.600 199.575 336.920 ;
        RECT 4.400 334.200 195.600 335.600 ;
        RECT 0.525 332.880 199.575 334.200 ;
        RECT 0.525 331.480 195.600 332.880 ;
        RECT 0.525 330.160 199.575 331.480 ;
        RECT 4.400 328.760 195.600 330.160 ;
        RECT 0.525 327.440 199.575 328.760 ;
        RECT 0.525 326.040 195.600 327.440 ;
        RECT 0.525 324.720 199.575 326.040 ;
        RECT 4.400 323.320 195.600 324.720 ;
        RECT 0.525 322.000 199.575 323.320 ;
        RECT 0.525 320.600 195.600 322.000 ;
        RECT 0.525 319.280 199.575 320.600 ;
        RECT 4.400 317.880 195.600 319.280 ;
        RECT 0.525 316.560 199.575 317.880 ;
        RECT 0.525 315.160 195.600 316.560 ;
        RECT 0.525 313.840 199.575 315.160 ;
        RECT 4.400 312.440 195.600 313.840 ;
        RECT 0.525 311.120 199.575 312.440 ;
        RECT 0.525 309.720 195.600 311.120 ;
        RECT 0.525 308.400 199.575 309.720 ;
        RECT 4.400 307.000 195.600 308.400 ;
        RECT 0.525 305.680 199.575 307.000 ;
        RECT 0.525 304.280 195.600 305.680 ;
        RECT 0.525 302.960 199.575 304.280 ;
        RECT 4.400 301.560 195.600 302.960 ;
        RECT 0.525 300.240 199.575 301.560 ;
        RECT 0.525 298.840 195.600 300.240 ;
        RECT 0.525 297.520 199.575 298.840 ;
        RECT 4.400 296.120 195.600 297.520 ;
        RECT 0.525 294.800 199.575 296.120 ;
        RECT 0.525 293.400 195.600 294.800 ;
        RECT 0.525 292.080 199.575 293.400 ;
        RECT 4.400 290.680 195.600 292.080 ;
        RECT 0.525 289.360 199.575 290.680 ;
        RECT 0.525 287.960 195.600 289.360 ;
        RECT 0.525 286.640 199.575 287.960 ;
        RECT 4.400 285.240 195.600 286.640 ;
        RECT 0.525 283.920 199.575 285.240 ;
        RECT 0.525 282.520 195.600 283.920 ;
        RECT 0.525 281.200 199.575 282.520 ;
        RECT 4.400 279.800 195.600 281.200 ;
        RECT 0.525 278.480 199.575 279.800 ;
        RECT 0.525 277.080 195.600 278.480 ;
        RECT 0.525 275.760 199.575 277.080 ;
        RECT 4.400 274.360 195.600 275.760 ;
        RECT 0.525 273.040 199.575 274.360 ;
        RECT 0.525 271.640 195.600 273.040 ;
        RECT 0.525 270.320 199.575 271.640 ;
        RECT 4.400 268.920 195.600 270.320 ;
        RECT 0.525 267.600 199.575 268.920 ;
        RECT 0.525 266.200 195.600 267.600 ;
        RECT 0.525 264.880 199.575 266.200 ;
        RECT 4.400 263.480 195.600 264.880 ;
        RECT 0.525 262.160 199.575 263.480 ;
        RECT 0.525 260.760 195.600 262.160 ;
        RECT 0.525 259.440 199.575 260.760 ;
        RECT 4.400 258.040 195.600 259.440 ;
        RECT 0.525 256.720 199.575 258.040 ;
        RECT 0.525 255.320 195.600 256.720 ;
        RECT 0.525 254.000 199.575 255.320 ;
        RECT 4.400 252.600 195.600 254.000 ;
        RECT 0.525 251.280 199.575 252.600 ;
        RECT 0.525 249.880 195.600 251.280 ;
        RECT 0.525 248.560 199.575 249.880 ;
        RECT 4.400 247.160 195.600 248.560 ;
        RECT 0.525 245.840 199.575 247.160 ;
        RECT 0.525 244.440 195.600 245.840 ;
        RECT 0.525 243.120 199.575 244.440 ;
        RECT 4.400 241.720 195.600 243.120 ;
        RECT 0.525 240.400 199.575 241.720 ;
        RECT 0.525 239.000 195.600 240.400 ;
        RECT 0.525 237.680 199.575 239.000 ;
        RECT 4.400 236.280 195.600 237.680 ;
        RECT 0.525 234.960 199.575 236.280 ;
        RECT 0.525 233.560 195.600 234.960 ;
        RECT 0.525 232.240 199.575 233.560 ;
        RECT 4.400 230.840 195.600 232.240 ;
        RECT 0.525 229.520 199.575 230.840 ;
        RECT 0.525 228.120 195.600 229.520 ;
        RECT 0.525 226.800 199.575 228.120 ;
        RECT 4.400 225.400 195.600 226.800 ;
        RECT 0.525 224.080 199.575 225.400 ;
        RECT 0.525 222.680 195.600 224.080 ;
        RECT 0.525 221.360 199.575 222.680 ;
        RECT 4.400 219.960 195.600 221.360 ;
        RECT 0.525 218.640 199.575 219.960 ;
        RECT 0.525 217.240 195.600 218.640 ;
        RECT 0.525 215.920 199.575 217.240 ;
        RECT 4.400 214.520 195.600 215.920 ;
        RECT 0.525 213.200 199.575 214.520 ;
        RECT 0.525 211.800 195.600 213.200 ;
        RECT 0.525 210.480 199.575 211.800 ;
        RECT 4.400 209.080 195.600 210.480 ;
        RECT 0.525 207.760 199.575 209.080 ;
        RECT 0.525 206.360 195.600 207.760 ;
        RECT 0.525 205.040 199.575 206.360 ;
        RECT 4.400 203.640 195.600 205.040 ;
        RECT 0.525 202.320 199.575 203.640 ;
        RECT 0.525 200.920 195.600 202.320 ;
        RECT 0.525 199.600 199.575 200.920 ;
        RECT 4.400 198.200 195.600 199.600 ;
        RECT 0.525 196.880 199.575 198.200 ;
        RECT 0.525 195.480 195.600 196.880 ;
        RECT 0.525 194.160 199.575 195.480 ;
        RECT 4.400 192.760 195.600 194.160 ;
        RECT 0.525 191.440 199.575 192.760 ;
        RECT 0.525 190.040 195.600 191.440 ;
        RECT 0.525 188.720 199.575 190.040 ;
        RECT 4.400 187.320 195.600 188.720 ;
        RECT 0.525 186.000 199.575 187.320 ;
        RECT 0.525 184.600 195.600 186.000 ;
        RECT 0.525 183.280 199.575 184.600 ;
        RECT 4.400 181.880 195.600 183.280 ;
        RECT 0.525 180.560 199.575 181.880 ;
        RECT 0.525 179.160 195.600 180.560 ;
        RECT 0.525 177.840 199.575 179.160 ;
        RECT 4.400 176.440 195.600 177.840 ;
        RECT 0.525 175.120 199.575 176.440 ;
        RECT 0.525 173.720 195.600 175.120 ;
        RECT 0.525 172.400 199.575 173.720 ;
        RECT 4.400 171.000 195.600 172.400 ;
        RECT 0.525 169.680 199.575 171.000 ;
        RECT 0.525 168.280 195.600 169.680 ;
        RECT 0.525 166.960 199.575 168.280 ;
        RECT 4.400 165.560 195.600 166.960 ;
        RECT 0.525 164.240 199.575 165.560 ;
        RECT 0.525 162.840 195.600 164.240 ;
        RECT 0.525 161.520 199.575 162.840 ;
        RECT 4.400 160.120 195.600 161.520 ;
        RECT 0.525 158.800 199.575 160.120 ;
        RECT 0.525 157.400 195.600 158.800 ;
        RECT 0.525 156.080 199.575 157.400 ;
        RECT 4.400 154.680 195.600 156.080 ;
        RECT 0.525 153.360 199.575 154.680 ;
        RECT 0.525 151.960 195.600 153.360 ;
        RECT 0.525 150.640 199.575 151.960 ;
        RECT 4.400 149.240 199.575 150.640 ;
        RECT 0.525 145.200 199.575 149.240 ;
        RECT 4.400 143.800 199.575 145.200 ;
        RECT 0.525 139.760 199.575 143.800 ;
        RECT 4.400 138.360 199.575 139.760 ;
        RECT 0.525 134.320 199.575 138.360 ;
        RECT 4.400 132.920 199.575 134.320 ;
        RECT 0.525 128.880 199.575 132.920 ;
        RECT 4.400 127.480 199.575 128.880 ;
        RECT 0.525 123.440 199.575 127.480 ;
        RECT 4.400 122.040 199.575 123.440 ;
        RECT 0.525 118.000 199.575 122.040 ;
        RECT 4.400 116.600 199.575 118.000 ;
        RECT 0.525 112.560 199.575 116.600 ;
        RECT 4.400 111.160 199.575 112.560 ;
        RECT 0.525 107.120 199.575 111.160 ;
        RECT 4.400 105.720 199.575 107.120 ;
        RECT 0.525 101.680 199.575 105.720 ;
        RECT 4.400 100.280 199.575 101.680 ;
        RECT 0.525 96.240 199.575 100.280 ;
        RECT 4.400 94.840 199.575 96.240 ;
        RECT 0.525 90.800 199.575 94.840 ;
        RECT 4.400 89.400 199.575 90.800 ;
        RECT 0.525 85.360 199.575 89.400 ;
        RECT 4.400 83.960 199.575 85.360 ;
        RECT 0.525 79.920 199.575 83.960 ;
        RECT 4.400 78.520 199.575 79.920 ;
        RECT 0.525 74.480 199.575 78.520 ;
        RECT 4.400 73.080 199.575 74.480 ;
        RECT 0.525 69.040 199.575 73.080 ;
        RECT 4.400 67.640 199.575 69.040 ;
        RECT 0.525 63.600 199.575 67.640 ;
        RECT 4.400 62.200 199.575 63.600 ;
        RECT 0.525 10.715 199.575 62.200 ;
      LAYER met4 ;
        RECT 2.135 72.935 20.640 1072.865 ;
        RECT 23.040 72.935 97.440 1072.865 ;
        RECT 99.840 72.935 174.240 1072.865 ;
        RECT 176.640 72.935 195.665 1072.865 ;
  END
END multiplexer
END LIBRARY

