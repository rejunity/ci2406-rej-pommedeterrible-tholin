// This is the unpowered netlist.
module ci2406_z80 (rst_n,
    wb_clk_i,
    custom_settings,
    io_in,
    io_oeb,
    io_out);
 input rst_n;
 input wb_clk_i;
 input [1:0] custom_settings;
 input [35:0] io_in;
 output [35:0] io_oeb;
 output [35:0] io_out;

 wire net182;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net183;
 wire net201;
 wire net202;
 wire net184;
 wire net211;
 wire net212;
 wire net203;
 wire net204;
 wire net205;
 wire net213;
 wire net185;
 wire net210;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net207;
 wire net208;
 wire net209;
 wire net206;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \z80.early_iorq_n ;
 wire \z80.early_mreq_n ;
 wire \z80.early_rd_n ;
 wire \z80.early_wr_n ;
 wire \z80.normal_iorq_n ;
 wire \z80.normal_mreq_n ;
 wire \z80.normal_rd_n ;
 wire \z80.normal_wr_n ;
 wire \z80.tv80s.di_reg[0] ;
 wire \z80.tv80s.di_reg[1] ;
 wire \z80.tv80s.di_reg[2] ;
 wire \z80.tv80s.di_reg[3] ;
 wire \z80.tv80s.di_reg[4] ;
 wire \z80.tv80s.di_reg[5] ;
 wire \z80.tv80s.di_reg[6] ;
 wire \z80.tv80s.di_reg[7] ;
 wire \z80.tv80s.i_tv80_core.ACC[0] ;
 wire \z80.tv80s.i_tv80_core.ACC[1] ;
 wire \z80.tv80s.i_tv80_core.ACC[2] ;
 wire \z80.tv80s.i_tv80_core.ACC[3] ;
 wire \z80.tv80s.i_tv80_core.ACC[4] ;
 wire \z80.tv80s.i_tv80_core.ACC[5] ;
 wire \z80.tv80s.i_tv80_core.ACC[6] ;
 wire \z80.tv80s.i_tv80_core.ACC[7] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[0] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[1] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[2] ;
 wire \z80.tv80s.i_tv80_core.ALU_Op_r[3] ;
 wire \z80.tv80s.i_tv80_core.Alternate ;
 wire \z80.tv80s.i_tv80_core.Ap[0] ;
 wire \z80.tv80s.i_tv80_core.Ap[1] ;
 wire \z80.tv80s.i_tv80_core.Ap[2] ;
 wire \z80.tv80s.i_tv80_core.Ap[3] ;
 wire \z80.tv80s.i_tv80_core.Ap[4] ;
 wire \z80.tv80s.i_tv80_core.Ap[5] ;
 wire \z80.tv80s.i_tv80_core.Ap[6] ;
 wire \z80.tv80s.i_tv80_core.Ap[7] ;
 wire \z80.tv80s.i_tv80_core.Arith16_r ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t1 ;
 wire \z80.tv80s.i_tv80_core.Auto_Wait_t2 ;
 wire \z80.tv80s.i_tv80_core.BTR_r ;
 wire \z80.tv80s.i_tv80_core.BusA[0] ;
 wire \z80.tv80s.i_tv80_core.BusA[1] ;
 wire \z80.tv80s.i_tv80_core.BusA[2] ;
 wire \z80.tv80s.i_tv80_core.BusA[3] ;
 wire \z80.tv80s.i_tv80_core.BusA[4] ;
 wire \z80.tv80s.i_tv80_core.BusA[5] ;
 wire \z80.tv80s.i_tv80_core.BusA[6] ;
 wire \z80.tv80s.i_tv80_core.BusA[7] ;
 wire \z80.tv80s.i_tv80_core.BusAck ;
 wire \z80.tv80s.i_tv80_core.BusB[0] ;
 wire \z80.tv80s.i_tv80_core.BusB[1] ;
 wire \z80.tv80s.i_tv80_core.BusB[2] ;
 wire \z80.tv80s.i_tv80_core.BusB[3] ;
 wire \z80.tv80s.i_tv80_core.BusB[4] ;
 wire \z80.tv80s.i_tv80_core.BusB[5] ;
 wire \z80.tv80s.i_tv80_core.BusB[6] ;
 wire \z80.tv80s.i_tv80_core.BusB[7] ;
 wire \z80.tv80s.i_tv80_core.BusReq_s ;
 wire \z80.tv80s.i_tv80_core.F[0] ;
 wire \z80.tv80s.i_tv80_core.F[1] ;
 wire \z80.tv80s.i_tv80_core.F[2] ;
 wire \z80.tv80s.i_tv80_core.F[3] ;
 wire \z80.tv80s.i_tv80_core.F[4] ;
 wire \z80.tv80s.i_tv80_core.F[5] ;
 wire \z80.tv80s.i_tv80_core.F[6] ;
 wire \z80.tv80s.i_tv80_core.F[7] ;
 wire \z80.tv80s.i_tv80_core.Fp[0] ;
 wire \z80.tv80s.i_tv80_core.Fp[1] ;
 wire \z80.tv80s.i_tv80_core.Fp[2] ;
 wire \z80.tv80s.i_tv80_core.Fp[3] ;
 wire \z80.tv80s.i_tv80_core.Fp[4] ;
 wire \z80.tv80s.i_tv80_core.Fp[5] ;
 wire \z80.tv80s.i_tv80_core.Fp[6] ;
 wire \z80.tv80s.i_tv80_core.Fp[7] ;
 wire \z80.tv80s.i_tv80_core.Halt_FF ;
 wire \z80.tv80s.i_tv80_core.INT_s ;
 wire \z80.tv80s.i_tv80_core.IR[0] ;
 wire \z80.tv80s.i_tv80_core.IR[1] ;
 wire \z80.tv80s.i_tv80_core.IR[2] ;
 wire \z80.tv80s.i_tv80_core.IR[3] ;
 wire \z80.tv80s.i_tv80_core.IR[4] ;
 wire \z80.tv80s.i_tv80_core.IR[5] ;
 wire \z80.tv80s.i_tv80_core.IR[6] ;
 wire \z80.tv80s.i_tv80_core.IR[7] ;
 wire \z80.tv80s.i_tv80_core.ISet[0] ;
 wire \z80.tv80s.i_tv80_core.ISet[1] ;
 wire \z80.tv80s.i_tv80_core.ISet[2] ;
 wire \z80.tv80s.i_tv80_core.ISet[3] ;
 wire \z80.tv80s.i_tv80_core.IStatus[1] ;
 wire \z80.tv80s.i_tv80_core.IStatus[2] ;
 wire \z80.tv80s.i_tv80_core.I[0] ;
 wire \z80.tv80s.i_tv80_core.I[1] ;
 wire \z80.tv80s.i_tv80_core.I[2] ;
 wire \z80.tv80s.i_tv80_core.I[3] ;
 wire \z80.tv80s.i_tv80_core.I[4] ;
 wire \z80.tv80s.i_tv80_core.I[5] ;
 wire \z80.tv80s.i_tv80_core.I[6] ;
 wire \z80.tv80s.i_tv80_core.I[7] ;
 wire \z80.tv80s.i_tv80_core.IncDecZ ;
 wire \z80.tv80s.i_tv80_core.IntCycle ;
 wire \z80.tv80s.i_tv80_core.IntE ;
 wire \z80.tv80s.i_tv80_core.IntE_FF2 ;
 wire \z80.tv80s.i_tv80_core.NMICycle ;
 wire \z80.tv80s.i_tv80_core.NMI_s ;
 wire \z80.tv80s.i_tv80_core.No_BTR ;
 wire \z80.tv80s.i_tv80_core.Oldnmi_n ;
 wire \z80.tv80s.i_tv80_core.PC[0] ;
 wire \z80.tv80s.i_tv80_core.PC[10] ;
 wire \z80.tv80s.i_tv80_core.PC[11] ;
 wire \z80.tv80s.i_tv80_core.PC[12] ;
 wire \z80.tv80s.i_tv80_core.PC[13] ;
 wire \z80.tv80s.i_tv80_core.PC[14] ;
 wire \z80.tv80s.i_tv80_core.PC[15] ;
 wire \z80.tv80s.i_tv80_core.PC[1] ;
 wire \z80.tv80s.i_tv80_core.PC[2] ;
 wire \z80.tv80s.i_tv80_core.PC[3] ;
 wire \z80.tv80s.i_tv80_core.PC[4] ;
 wire \z80.tv80s.i_tv80_core.PC[5] ;
 wire \z80.tv80s.i_tv80_core.PC[6] ;
 wire \z80.tv80s.i_tv80_core.PC[7] ;
 wire \z80.tv80s.i_tv80_core.PC[8] ;
 wire \z80.tv80s.i_tv80_core.PC[9] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ;
 wire \z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ;
 wire \z80.tv80s.i_tv80_core.PreserveC_r ;
 wire \z80.tv80s.i_tv80_core.R[0] ;
 wire \z80.tv80s.i_tv80_core.R[1] ;
 wire \z80.tv80s.i_tv80_core.R[2] ;
 wire \z80.tv80s.i_tv80_core.R[3] ;
 wire \z80.tv80s.i_tv80_core.R[4] ;
 wire \z80.tv80s.i_tv80_core.R[5] ;
 wire \z80.tv80s.i_tv80_core.R[6] ;
 wire \z80.tv80s.i_tv80_core.R[7] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ;
 wire \z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrB_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[0] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[1] ;
 wire \z80.tv80s.i_tv80_core.RegAddrC[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[0] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[10] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[11] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[12] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[13] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[14] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[15] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[1] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[2] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[3] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[4] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[5] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[6] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[7] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[8] ;
 wire \z80.tv80s.i_tv80_core.RegBusA_r[9] ;
 wire \z80.tv80s.i_tv80_core.SP[0] ;
 wire \z80.tv80s.i_tv80_core.SP[10] ;
 wire \z80.tv80s.i_tv80_core.SP[11] ;
 wire \z80.tv80s.i_tv80_core.SP[12] ;
 wire \z80.tv80s.i_tv80_core.SP[13] ;
 wire \z80.tv80s.i_tv80_core.SP[14] ;
 wire \z80.tv80s.i_tv80_core.SP[15] ;
 wire \z80.tv80s.i_tv80_core.SP[1] ;
 wire \z80.tv80s.i_tv80_core.SP[2] ;
 wire \z80.tv80s.i_tv80_core.SP[3] ;
 wire \z80.tv80s.i_tv80_core.SP[4] ;
 wire \z80.tv80s.i_tv80_core.SP[5] ;
 wire \z80.tv80s.i_tv80_core.SP[6] ;
 wire \z80.tv80s.i_tv80_core.SP[7] ;
 wire \z80.tv80s.i_tv80_core.SP[8] ;
 wire \z80.tv80s.i_tv80_core.SP[9] ;
 wire \z80.tv80s.i_tv80_core.Save_ALU_r ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[0] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[10] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[11] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[12] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[13] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[14] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[15] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[1] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[2] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[3] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[4] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[5] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[6] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[7] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[8] ;
 wire \z80.tv80s.i_tv80_core.TmpAddr[9] ;
 wire \z80.tv80s.i_tv80_core.XY_Ind ;
 wire \z80.tv80s.i_tv80_core.XY_State[0] ;
 wire \z80.tv80s.i_tv80_core.XY_State[1] ;
 wire \z80.tv80s.i_tv80_core.Z16_r ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ;
 wire \z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ;
 wire \z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ;
 wire \z80.tv80s.i_tv80_core.mcycles[1] ;
 wire \z80.tv80s.i_tv80_core.mcycles[2] ;
 wire \z80.tv80s.i_tv80_core.mcycles[4] ;
 wire \z80.tv80s.i_tv80_core.mcycles[5] ;
 wire \z80.tv80s.i_tv80_core.ts[0] ;
 wire \z80.tv80s.i_tv80_core.ts[1] ;
 wire \z80.tv80s.i_tv80_core.ts[2] ;
 wire \z80.tv80s.i_tv80_core.ts[3] ;
 wire \z80.tv80s.i_tv80_core.ts[4] ;
 wire \z80.tv80s.i_tv80_core.ts[5] ;
 wire \z80.tv80s.i_tv80_core.ts[6] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0511_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_1532_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_2170_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\z80.tv80s.i_tv80_core.ISet[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_1296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3045__A (.DIODE(\z80.tv80s.i_tv80_core.ts[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__A (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__A (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__A (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__A (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__C (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__B (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__B (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A_N (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__C (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A_N (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__A (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__B (.DIODE(_2890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__D_N (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__B (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A_N (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A_N (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__B (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__D_N (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__B (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__B (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A2 (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__C (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__B (.DIODE(_2943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__A (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__B (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__B (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__B (.DIODE(_2943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A2 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A2 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A3 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3189__A (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__B (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__B (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__B (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__B (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A1 (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__B (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__D (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A2 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__B (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3220__B (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__B (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__C (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__A (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__B (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A (.DIODE(_2943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__B (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__B (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__C_N (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A1 (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A2 (.DIODE(_2943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__B1 (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__B (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A3 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__B1 (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A3 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A4 (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A3 (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__C (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__C (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__D (.DIODE(_2947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__B (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__B (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3261__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__B (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__B1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__C1 (.DIODE(_2947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__B1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__B2 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__B1 (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__A (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A2 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__B (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__B (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__B (.DIODE(_2943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__D1 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__B (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__C1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__D1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A1 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__B (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__B (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__A2 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__A2 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__B1 (.DIODE(_2943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A1 (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__C (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__B (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__C (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__A0 (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__S (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__B (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A0 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__S (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__B1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__B1 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__B1 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__B1 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__B (.DIODE(_2947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__B (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__B (.DIODE(_2943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__B (.DIODE(_2943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__B (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A1 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__B2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__B (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__B (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__B (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__C_N (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A_N (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__B (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__C (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__C (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__B (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A1 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__B1 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__B (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__D1 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__C1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A2 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__B (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A3 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__C1 (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A1 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A_N (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__B (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__B1 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__B (.DIODE(_2890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__C (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__D_N (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__B (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__B (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__C (.DIODE(_2890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__D (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__B (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A2 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__B (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__B (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A2 (.DIODE(\z80.tv80s.i_tv80_core.ts[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A3 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A2 (.DIODE(\z80.tv80s.i_tv80_core.ts[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A3 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A1 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__B1_N (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__C (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__B (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__C (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__B (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A2 (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__B2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__B2 (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A2 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A3 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A2 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__C1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A2 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__A (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__D (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__C1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__B (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__C (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__B2 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__B2 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__B (.DIODE(\z80.tv80s.i_tv80_core.IR[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__C (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A3 (.DIODE(_2949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A4 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A3 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__A1 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__B1 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__C1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__B1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__A1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A2 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A2 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A1 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__B1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__B (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__B (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A2 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A1 (.DIODE(_2876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A2 (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__B (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A2 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__B (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A1 (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A2 (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__S (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__B (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A2 (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__A1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__B2 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B1 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__B (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__B1 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__C1 (.DIODE(_2833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__B (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__B (.DIODE(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A (.DIODE(_2947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__B (.DIODE(_2947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__D_N (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__C (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__C (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__D (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__B (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A1 (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A2 (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__B (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3655__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__B (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3660__B1 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A1 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3667__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__A1_N (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3671__B2 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3673__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A1 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__B1 (.DIODE(_2996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__B1 (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3678__A2 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3679__A1 (.DIODE(_2946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A2 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3685__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A2 (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__C_N (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__A2 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3696__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__C1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3697__D1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3698__B1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__B1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3701__A1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3703__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3708__C1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3711__B1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__C1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__C (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3717__A (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3718__B (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3721__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__S0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__S1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__3723__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__B (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3730__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3731__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3732__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__C (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A3 (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__C1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__C (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__3752__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A1 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3753__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__D (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__C (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3762__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A2 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__B (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__B (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__A2 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__C1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__C (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__C (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__C (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__C (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__C (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3792__C (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__C (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3806__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3807__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3815__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3816__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__B (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3820__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3821__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3829__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3830__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__S (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3834__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__S (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__S (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3838__S (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3839__S (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A2 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__C1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__B (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3859__A1 (.DIODE(_0805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__S (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3881__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3883__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3901__A (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__B (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__S (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A2 (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3913__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3914__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__S1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3923__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3926__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3927__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3928__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3936__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3961__A2 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3965__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3967__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3978__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__C (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3980__B1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3982__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3984__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3988__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3994__A (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A2 (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3996__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3997__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4005__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4007__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4015__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4016__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__B (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4028__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4031__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A2 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4049__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__A2 (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4052__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4068__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4070__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4076__S (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4080__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__B1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A2 (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4090__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4107__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4126__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4135__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4136__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A1 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A1 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A2 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__A2 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__S1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__A2 (.DIODE(_0880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4151__B1 (.DIODE(_0882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__A2 (.DIODE(_0875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4152__B1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__B1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A2 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__B1 (.DIODE(_0890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4164__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__B (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4169__A3 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4171__A0 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4175__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4181__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4183__A (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A1 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__A2 (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4185__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4188__A (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__A (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4194__A2 (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4196__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__B (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__B (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4198__C (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__4202__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A1 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4204__A1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4211__B (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4213__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__C (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__A2 (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4215__B1 (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A2 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__A3 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4219__A2 (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__A (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4221__A (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__B (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__C (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4225__A1 (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4227__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__4231__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A3 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__B1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__A2 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4233__A3 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A1 (.DIODE(\z80.tv80s.i_tv80_core.IR[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__A2 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4235__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A1 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4237__A2 (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__A3 (.DIODE(_2880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4239__B1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__A (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__B (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__4247__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__A (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A1 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4249__A3 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4251__C1 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4253__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__A2 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4255__B (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__A2 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4257__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__A2 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__B1 (.DIODE(_0442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4259__A1 (.DIODE(_2824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4261__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__4263__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__A (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4265__A2 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__A2 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4267__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A1 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4272__A2 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__B2 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__4278__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__B (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__B (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4284__C (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__C (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__B (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4286__C_N (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__B (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4288__S (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__A3 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__B1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B2 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__S (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A4 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__B (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4300__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__A1 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A2 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__S (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4308__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__4310__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A2 (.DIODE(_1372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__C (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__B (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4321__B (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__B1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__4323__A (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__4325__A0 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__S (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__S (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__S (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__S (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__S (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__S (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__S (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S (.DIODE(_1405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__A (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A1_N (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A2_N (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__S (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4354__S (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4355__S (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4356__S (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__S (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__S (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__S (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__S (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__C_N (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4364__S1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4372__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A1 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A2 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__B (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__B1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A1 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A2 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__A1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4391__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__A1 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__C1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__S0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__C1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__S0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__S1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__S1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__S0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4427__S (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__S (.DIODE(_1415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__S (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4431__S (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__S (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__S (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__S (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__S (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__S (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__S (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__S (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__S (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A1 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__S (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__S (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4443__S (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4444__S (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__S (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__S (.DIODE(_1474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__S (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__S (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__S (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4451__S (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__S (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__S (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__S (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__S (.DIODE(_1475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__S (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__S (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__A0 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__S (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4460__S (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__S (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__S (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__S (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__S (.DIODE(_1476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__S (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__S (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A0 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__S (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__S (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__S (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__S (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__S (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__S (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A0 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__S (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__S (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__S (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A1 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__S (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__S (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4488__S (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4489__S (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__S (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__S (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4492__A (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__S (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__S (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__S (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A1 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__S (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__S (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__S (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__S (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__S (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__S (.DIODE(_1481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A (.DIODE(_0792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S (.DIODE(_1482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__B (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__B (.DIODE(_2960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__B (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__C (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4523__B (.DIODE(_1486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4538__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__B1 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__B (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A2 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A3 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__B (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A2 (.DIODE(_2949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__B2 (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__C1 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A3 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__B (.DIODE(_2949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B (.DIODE(_2949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__B (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__S (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__A (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__C (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__B (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__D (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A_N (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4573__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__B (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A2 (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A1 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__S (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__S (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__S (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__A (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__B (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__A2 (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__B2 (.DIODE(_1540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__B (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A2 (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__S (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusAck ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__B1 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A2 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__B1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A2 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__B1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A2 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A2 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__B1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A2 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__B1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__4627__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A2 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__B1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A2 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__B1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__B (.DIODE(_1551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A2 (.DIODE(_1554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__B1 (.DIODE(_1556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__C (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__B (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__B (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__S (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__B (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__D (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__S (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__S (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__S (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__S (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4664__S (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4667__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4669__S (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4670__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__A (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__S (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4675__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4677__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__A (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__B (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__D (.DIODE(_2950_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__4680__B (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A1_N (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__B (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__A (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__B (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__S (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4687__B1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A2 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4689__A2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4690__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4692__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4693__S (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4696__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__S (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__B1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__S (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__B1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4705__S (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4711__S (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__B1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A0 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__S (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__S (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__B1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__S (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4725__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4726__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__A0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__4727__S (.DIODE(_1370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A1_N (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__B1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4729__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__S (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A0 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__S (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4732__S (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4733__B1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4734__B (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4735__B1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S0 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__S1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S0 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__S1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__A2 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__4749__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__4750__B (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__A1 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4759__B2 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4761__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4762__A0 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4770__A1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4771__B1 (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4773__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__B (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__B1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__C1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4783__A2 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S0 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4784__S1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S0 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__S1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__S (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__B (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__A1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4789__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4790__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4792__A (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__B (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B2 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A1 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A2 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B1 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__C1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A2 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__B (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A0 (.DIODE(_1720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B2 (.DIODE(_1720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A2 (.DIODE(_1720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__B1 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__C1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A2 (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__B1 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4827__B (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__S (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A1 (.DIODE(_0496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__C1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__B2 (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4833__B1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4838__C1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4839__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A2 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__B1 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__B (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A0 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__B2 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4851__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A2 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__C1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__B (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A2 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__B (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A0 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__B2 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A1 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__B (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A2 (.DIODE(_1667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__S (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A0 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__B1_N (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__B2 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__S0 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__S1 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S0 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__S1 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__S (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4900__B (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__S (.DIODE(_0499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A0 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__A2 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__B1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__B (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__C (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__D (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__B (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A1 (.DIODE(_1689_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__C1 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B2 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__S1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__S0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__S1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__B1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A0 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__B (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__B1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A0 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__S (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4952__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__B (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__B1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A0 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__S (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__S (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__B1 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A2 (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__A0 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5011__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__S1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__S (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__S (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5031__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__B1 (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A0 (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A0 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__S (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A0 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__S0 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__S0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5052__S1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__S (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A0 (.DIODE(\z80.tv80s.i_tv80_core.PC[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__S (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__S (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__S (.DIODE(_1685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__B2 (.DIODE(_1678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__C_N (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5071__A (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A2 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A2 (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A2 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A2 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1_N (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__C1 (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__B (.DIODE(_3002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__B (.DIODE(_1994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A2 (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B1_N (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5118__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A2 (.DIODE(_2881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__B2 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__S (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B1_N (.DIODE(_1994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__B (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__B (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__B (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__B (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5166__B2 (.DIODE(_1994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A2 (.DIODE(_3004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B1 (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A1 (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A2 (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__S (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A2 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A2 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__S (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B2 (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__A2 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__S (.DIODE(_1602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__S (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A2 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A0 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A1 (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A2 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__S (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__C1 (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A2 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__B (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__C (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__D (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B2 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A1 (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A0 (.DIODE(_2114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__B (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__C (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5229__D (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__C (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__D (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__B1 (.DIODE(_1994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__A1 (.DIODE(_1994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__S (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A0 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__S (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A0 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__S (.DIODE(_1608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A1 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__S (.DIODE(_1994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A0 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__S (.DIODE(_1969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__B (.DIODE(_0721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A2 (.DIODE(_2138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__B2 (.DIODE(_2114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__C1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__B (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__B1 (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A2 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B1 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__C1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A2 (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__C (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A2 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B1 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A2 (.DIODE(_2823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A2 (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__C (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(\z80.tv80s.i_tv80_core.IR[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A2 (.DIODE(_2949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A2 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A2 (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A2 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__B (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__C1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__A1 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5310__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A2 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A1_N (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5313__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__D (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A3 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A1 (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A1 (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__B1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__C (.DIODE(_1491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A1 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__A3 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A0 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1_N (.DIODE(_2949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A0 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__5361__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__C (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A1 (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A2 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A3 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__B (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__B (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__A (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A3 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__S (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A2 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__B2 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A1 (.DIODE(_1720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A2 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__B2 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__B (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A0 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A1 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A0 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A0 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__B (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A0 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A1 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A1 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A2_N (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__B2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A0 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A1 (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A2 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A2_N (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__S (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__S (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A1 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A2 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__B (.DIODE(_2346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__A2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__A3 (.DIODE(_2346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A1 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A2 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A1 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A1 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A2 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B2 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A2_N (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A1 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__S (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A2_N (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A1 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A2 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__B2 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A1 (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A2_N (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B2 (.DIODE(_2241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A1 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__S (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A2 (.DIODE(_2248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B2 (.DIODE(_2240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__S (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__D (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__B1 (.DIODE(_0692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__B2 (.DIODE(_0383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A2 (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A2 (.DIODE(_2940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__C1 (.DIODE(_2942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B (.DIODE(_2949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A1 (.DIODE(_0395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__C (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__C (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__D (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__B1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5592__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__B1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__C1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A2 (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__C1 (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A2 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__C1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__B (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__B (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5602__A (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__B (.DIODE(_1365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__D (.DIODE(_2440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A3 (.DIODE(_2452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__B2 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A1 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__S (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__S (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__B2 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A1 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__B2 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__S (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__S (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A2 (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__S0 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__S1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B2 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__S0 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__S1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__B2 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__S0 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__S1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__B2 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5672__C1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__C1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__C1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__C1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__S0 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__S1 (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__B2 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A1 (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A1 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__C1 (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A2 (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__S (.DIODE(_1286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__S (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__B2 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A (.DIODE(_2831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__C (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__S (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__S (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__S (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__S (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__S (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A1 (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__S (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__S (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A1 (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__S (.DIODE(_2545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A0 (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A (.DIODE(_1315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__D (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A2 (.DIODE(_2548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A2 (.DIODE(_2548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__B1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A (.DIODE(_2964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__B2 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A2 (.DIODE(_0513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A2 (.DIODE(_2890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__A3 (.DIODE(_0392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__C1 (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__A (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A3 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__C1 (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__B1 (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A2 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A3 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A2 (.DIODE(_1652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__C1 (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B2 (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A2 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A3 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__S (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__B2 (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A2 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A3 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__S (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A2 (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__B2 (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A2 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A3 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A1 (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__B2 (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A2 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A3 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__S (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__S (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A2 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A3 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__S (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A2 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A3 (.DIODE(_0690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__B1 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A (.DIODE(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A (.DIODE(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A1 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A0 (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__S (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A0 (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__S (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A0 (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A1_N (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__B2 (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A2 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A0 (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__B2 (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A0 (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__S (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A2 (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A3 (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A0 (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__S (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A0 (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__B2 (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A0 (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B2 (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A1 (.DIODE(\z80.tv80s.i_tv80_core.PC[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A0 (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__S (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__S (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__S (.DIODE(_2549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__B1 (.DIODE(net845));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A2 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B (.DIODE(_0578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__B1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A2 (.DIODE(_0733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A0 (.DIODE(_1442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A0 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__S (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A0 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__S (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A0 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__S (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A0 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__S (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A0 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__S (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A0 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__S (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A0 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__S (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A0 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__S (.DIODE(_0599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A0 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__S (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A (.DIODE(_0579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A1 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__B2 (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__D_N (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__B1 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__B2 (.DIODE(_1656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__A2 (.DIODE(_1700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__A2 (.DIODE(_1720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__B2 (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__B2 (.DIODE(_1754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__B2 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__B2 (.DIODE(_1790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__B2 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__A (.DIODE(_1281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A2 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B2 (.DIODE(_1826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__B1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__B2 (.DIODE(_1843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__B1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A2 (.DIODE(_1862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__B1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A (.DIODE(_1086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A2_N (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__B1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A (.DIODE(_1140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__B1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A (.DIODE(_1177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__B (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__B (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A3 (.DIODE(_2761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__C (.DIODE(_1934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__B1 (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A1_N (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A2_N (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__S (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A0 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__S (.DIODE(_2790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__S (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__SET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__D (.DIODE(_0018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__SET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__D (.DIODE(_0017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__SET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__D (.DIODE(_0018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__SET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__D (.DIODE(_0017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__SET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__D (.DIODE(_0033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6250__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__RESET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__SET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__SET_B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__RESET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6333__RESET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__RESET_B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__RESET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__RESET_B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__RESET_B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__CLK (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__RESET_B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__RESET_B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__RESET_B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__SET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__SET_B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__SET_B (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__SET_B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_wb_clk_i_A (.DIODE(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_wb_clk_i_A (.DIODE(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_wb_clk_i_A (.DIODE(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_wb_clk_i_A (.DIODE(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(\z80.tv80s.i_tv80_core.BusAck ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(\z80.tv80s.i_tv80_core.BusAck ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(\z80.tv80s.i_tv80_core.IR[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(_1664_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(_0817_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(_1399_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(_1398_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_2884_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(_1668_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold316_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold365_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold375_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold401_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold403_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold409_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold420_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold423_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold425_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold429_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold433_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold439_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold441_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold447_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold457_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold461_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold470_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold474_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold496_A (.DIODE(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold500_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold510_A (.DIODE(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold518_A (.DIODE(\z80.tv80s.i_tv80_core.PC[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold532_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold538_A (.DIODE(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold542_A (.DIODE(\z80.tv80s.i_tv80_core.PC[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold544_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold549_A (.DIODE(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold551_A (.DIODE(\z80.tv80s.i_tv80_core.ts[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold583_A (.DIODE(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold590_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold592_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold595_A (.DIODE(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold599_A (.DIODE(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold600_A (.DIODE(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold601_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold603_A (.DIODE(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold606_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold608_A (.DIODE(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold610_A (.DIODE(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold612_A (.DIODE(\z80.tv80s.i_tv80_core.BusAck ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold613_A (.DIODE(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold616_A (.DIODE(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold617_A (.DIODE(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold619_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold628_A (.DIODE(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold630_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold631_A (.DIODE(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold632_A (.DIODE(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold637_A (.DIODE(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold641_A (.DIODE(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold642_A (.DIODE(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold643_A (.DIODE(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold644_A (.DIODE(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold645_A (.DIODE(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold646_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold647_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold648_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold649_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold652_A (.DIODE(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold653_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold656_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold658_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold661_A (.DIODE(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold662_A (.DIODE(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold663_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold667_A (.DIODE(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold669_A (.DIODE(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold670_A (.DIODE(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold671_A (.DIODE(\z80.tv80s.i_tv80_core.IR[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_output23_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net49));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_8 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_92 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkinv_4 _3032_ (.A(net123),
    .Y(_2819_));
 sky130_fd_sc_hd__inv_2 _3033_ (.A(net156),
    .Y(_2820_));
 sky130_fd_sc_hd__inv_2 _3034_ (.A(net151),
    .Y(_2821_));
 sky130_fd_sc_hd__inv_2 _3035_ (.A(net150),
    .Y(_2822_));
 sky130_fd_sc_hd__clkinv_4 _3036_ (.A(net144),
    .Y(_2823_));
 sky130_fd_sc_hd__inv_2 _3037_ (.A(net139),
    .Y(_2824_));
 sky130_fd_sc_hd__clkinv_4 _3038_ (.A(net125),
    .Y(_2825_));
 sky130_fd_sc_hd__inv_2 _3039_ (.A(net127),
    .Y(_2826_));
 sky130_fd_sc_hd__inv_2 _3040_ (.A(net161),
    .Y(_2827_));
 sky130_fd_sc_hd__inv_2 _3041_ (.A(\z80.tv80s.i_tv80_core.F[6] ),
    .Y(_2828_));
 sky130_fd_sc_hd__clkinv_4 _3042_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .Y(_2829_));
 sky130_fd_sc_hd__inv_2 _3043_ (.A(net761),
    .Y(_2830_));
 sky130_fd_sc_hd__inv_4 _3044_ (.A(net116),
    .Y(_2831_));
 sky130_fd_sc_hd__inv_2 _3045_ (.A(\z80.tv80s.i_tv80_core.ts[1] ),
    .Y(_2832_));
 sky130_fd_sc_hd__inv_2 _3046_ (.A(net118),
    .Y(net23));
 sky130_fd_sc_hd__inv_2 _3047_ (.A(net635),
    .Y(_2833_));
 sky130_fd_sc_hd__inv_2 _3048_ (.A(net773),
    .Y(net46));
 sky130_fd_sc_hd__inv_2 _3049_ (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .Y(_2834_));
 sky130_fd_sc_hd__inv_2 _3050_ (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .Y(_2835_));
 sky130_fd_sc_hd__inv_2 _3051_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .Y(_2836_));
 sky130_fd_sc_hd__inv_2 _3052_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .Y(_2837_));
 sky130_fd_sc_hd__inv_2 _3053_ (.A(net136),
    .Y(_2838_));
 sky130_fd_sc_hd__inv_2 _3054_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .Y(_2839_));
 sky130_fd_sc_hd__inv_2 _3055_ (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .Y(_2840_));
 sky130_fd_sc_hd__inv_2 _3056_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .Y(_2841_));
 sky130_fd_sc_hd__inv_2 _3057_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .Y(_2842_));
 sky130_fd_sc_hd__inv_2 _3058_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .Y(_2843_));
 sky130_fd_sc_hd__inv_2 _3059_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .Y(_2844_));
 sky130_fd_sc_hd__inv_2 _3060_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .Y(_2845_));
 sky130_fd_sc_hd__inv_2 _3061_ (.A(net582),
    .Y(_2846_));
 sky130_fd_sc_hd__inv_2 _3062_ (.A(net691),
    .Y(_2847_));
 sky130_fd_sc_hd__inv_2 _3063_ (.A(net642),
    .Y(_2848_));
 sky130_fd_sc_hd__inv_2 _3064_ (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .Y(_2849_));
 sky130_fd_sc_hd__inv_2 _3065_ (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .Y(_2850_));
 sky130_fd_sc_hd__inv_2 _3066_ (.A(net798),
    .Y(_2851_));
 sky130_fd_sc_hd__inv_2 _3067_ (.A(\z80.tv80s.di_reg[0] ),
    .Y(_2852_));
 sky130_fd_sc_hd__inv_2 _3068_ (.A(\z80.tv80s.di_reg[2] ),
    .Y(_2853_));
 sky130_fd_sc_hd__inv_2 _3069_ (.A(net630),
    .Y(_2854_));
 sky130_fd_sc_hd__inv_2 _3070_ (.A(net531),
    .Y(_2855_));
 sky130_fd_sc_hd__inv_2 _3071_ (.A(net535),
    .Y(_2856_));
 sky130_fd_sc_hd__inv_2 _3072_ (.A(net866),
    .Y(_2857_));
 sky130_fd_sc_hd__inv_2 _3073_ (.A(net624),
    .Y(_2858_));
 sky130_fd_sc_hd__inv_2 _3074_ (.A(\z80.tv80s.i_tv80_core.ACC[3] ),
    .Y(_2859_));
 sky130_fd_sc_hd__inv_2 _3075_ (.A(\z80.tv80s.i_tv80_core.ACC[5] ),
    .Y(_2860_));
 sky130_fd_sc_hd__inv_2 _3076_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .Y(_2861_));
 sky130_fd_sc_hd__inv_2 _3077_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .Y(_2862_));
 sky130_fd_sc_hd__inv_2 _3078_ (.A(net559),
    .Y(_2863_));
 sky130_fd_sc_hd__inv_2 _3079_ (.A(net560),
    .Y(_2864_));
 sky130_fd_sc_hd__inv_2 _3080_ (.A(net570),
    .Y(_2865_));
 sky130_fd_sc_hd__inv_2 _3081_ (.A(net781),
    .Y(_2866_));
 sky130_fd_sc_hd__inv_2 _3082_ (.A(net11),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _3083_ (.A(net12),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _3084__1 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net214));
 sky130_fd_sc_hd__o31a_2 _3085_ (.A1(net159),
    .A2(net680),
    .A3(net473),
    .B1(net123),
    .X(_2867_));
 sky130_fd_sc_hd__and2_4 _3086_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2868_));
 sky130_fd_sc_hd__nand2_8 _3087_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2869_));
 sky130_fd_sc_hd__nor2_2 _3088_ (.A(net144),
    .B(net141),
    .Y(_2870_));
 sky130_fd_sc_hd__or2_4 _3089_ (.A(net143),
    .B(net140),
    .X(_2871_));
 sky130_fd_sc_hd__nor2_1 _3090_ (.A(_2869_),
    .B(_2871_),
    .Y(_2872_));
 sky130_fd_sc_hd__or4bb_2 _3091_ (.A(net143),
    .B(net140),
    .C_N(\z80.tv80s.i_tv80_core.IR[7] ),
    .D_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2873_));
 sky130_fd_sc_hd__nand2_1 _3092_ (.A(net155),
    .B(net156),
    .Y(_2874_));
 sky130_fd_sc_hd__nor2_1 _3093_ (.A(net152),
    .B(_2874_),
    .Y(_2875_));
 sky130_fd_sc_hd__nand3b_4 _3094_ (.A_N(net151),
    .B(net156),
    .C(net154),
    .Y(_2876_));
 sky130_fd_sc_hd__nor2_2 _3095_ (.A(net114),
    .B(_2876_),
    .Y(_2877_));
 sky130_fd_sc_hd__and2_1 _3096_ (.A(_2872_),
    .B(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__nor2_2 _3097_ (.A(net148),
    .B(_2823_),
    .Y(_2879_));
 sky130_fd_sc_hd__nand2_2 _3098_ (.A(net114),
    .B(net143),
    .Y(_2880_));
 sky130_fd_sc_hd__and3b_4 _3099_ (.A_N(net150),
    .B(net144),
    .C(net141),
    .X(_2881_));
 sky130_fd_sc_hd__nand2_4 _3100_ (.A(net139),
    .B(_2879_),
    .Y(_2882_));
 sky130_fd_sc_hd__nand2b_4 _3101_ (.A_N(net156),
    .B(net154),
    .Y(_2883_));
 sky130_fd_sc_hd__nor2_1 _3102_ (.A(_2821_),
    .B(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__or2_4 _3103_ (.A(_2821_),
    .B(_2883_),
    .X(_2885_));
 sky130_fd_sc_hd__nor2_2 _3104_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2886_));
 sky130_fd_sc_hd__or2_4 _3105_ (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2887_));
 sky130_fd_sc_hd__nor2_2 _3106_ (.A(_2885_),
    .B(_2887_),
    .Y(_2888_));
 sky130_fd_sc_hd__nand2_2 _3107_ (.A(net88),
    .B(_2886_),
    .Y(_2889_));
 sky130_fd_sc_hd__nor2_2 _3108_ (.A(_2882_),
    .B(_2889_),
    .Y(_2890_));
 sky130_fd_sc_hd__nand2_1 _3109_ (.A(_2881_),
    .B(_2888_),
    .Y(_2891_));
 sky130_fd_sc_hd__or2_1 _3110_ (.A(_2878_),
    .B(_2890_),
    .X(_2892_));
 sky130_fd_sc_hd__or3_4 _3111_ (.A(net155),
    .B(_2821_),
    .C(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(_2893_));
 sky130_fd_sc_hd__or3_2 _3112_ (.A(net154),
    .B(_2820_),
    .C(net151),
    .X(_2894_));
 sky130_fd_sc_hd__or4b_4 _3113_ (.A(net155),
    .B(net151),
    .C(\z80.tv80s.i_tv80_core.IR[3] ),
    .D_N(net156),
    .X(_2895_));
 sky130_fd_sc_hd__nor2_1 _3114_ (.A(net152),
    .B(\z80.tv80s.i_tv80_core.IR[3] ),
    .Y(_2896_));
 sky130_fd_sc_hd__or3_2 _3115_ (.A(net151),
    .B(\z80.tv80s.i_tv80_core.IR[3] ),
    .C(_2883_),
    .X(_2897_));
 sky130_fd_sc_hd__and3_1 _3116_ (.A(_2893_),
    .B(_2895_),
    .C(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__nor2_1 _3117_ (.A(net154),
    .B(net156),
    .Y(_2899_));
 sky130_fd_sc_hd__or3_4 _3118_ (.A(net155),
    .B(net156),
    .C(net152),
    .X(_2900_));
 sky130_fd_sc_hd__or2_2 _3119_ (.A(_2822_),
    .B(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__nand2_1 _3120_ (.A(net151),
    .B(net146),
    .Y(_2902_));
 sky130_fd_sc_hd__nand2_1 _3121_ (.A(_2821_),
    .B(net146),
    .Y(_2903_));
 sky130_fd_sc_hd__o22a_1 _3122_ (.A1(net154),
    .A2(_2902_),
    .B1(_2903_),
    .B2(_2820_),
    .X(_2904_));
 sky130_fd_sc_hd__nand2_1 _3123_ (.A(net140),
    .B(_2886_),
    .Y(_2905_));
 sky130_fd_sc_hd__or2_2 _3124_ (.A(net143),
    .B(_2905_),
    .X(_2906_));
 sky130_fd_sc_hd__a31o_1 _3125_ (.A1(_2893_),
    .A2(_2901_),
    .A3(_2904_),
    .B1(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__o211a_1 _3126_ (.A1(net156),
    .A2(_2893_),
    .B1(_2895_),
    .C1(_2897_),
    .X(_2908_));
 sky130_fd_sc_hd__and3_1 _3127_ (.A(net142),
    .B(_2824_),
    .C(_2868_),
    .X(_2909_));
 sky130_fd_sc_hd__or3_2 _3128_ (.A(_2823_),
    .B(net140),
    .C(_2869_),
    .X(_2910_));
 sky130_fd_sc_hd__and2b_2 _3129_ (.A_N(net142),
    .B(net139),
    .X(_2911_));
 sky130_fd_sc_hd__nand2b_4 _3130_ (.A_N(net144),
    .B(net141),
    .Y(_2912_));
 sky130_fd_sc_hd__nor2_4 _3131_ (.A(_2869_),
    .B(_2912_),
    .Y(_2913_));
 sky130_fd_sc_hd__nand2_1 _3132_ (.A(_2868_),
    .B(_2911_),
    .Y(_2914_));
 sky130_fd_sc_hd__a21o_1 _3133_ (.A1(_2910_),
    .A2(_2914_),
    .B1(_2908_),
    .X(_2915_));
 sky130_fd_sc_hd__o211ai_1 _3134_ (.A1(_2873_),
    .A2(_2898_),
    .B1(_2907_),
    .C1(_2915_),
    .Y(_2916_));
 sky130_fd_sc_hd__or3_1 _3135_ (.A(net151),
    .B(net114),
    .C(_2883_),
    .X(_2917_));
 sky130_fd_sc_hd__or3_4 _3136_ (.A(net154),
    .B(_2820_),
    .C(_2821_),
    .X(_2918_));
 sky130_fd_sc_hd__o21ai_1 _3137_ (.A1(net146),
    .A2(_2918_),
    .B1(_2917_),
    .Y(_2919_));
 sky130_fd_sc_hd__or4bb_4 _3138_ (.A(net154),
    .B(net151),
    .C_N(net146),
    .D_N(net156),
    .X(_2920_));
 sky130_fd_sc_hd__and2b_2 _3139_ (.A_N(net139),
    .B(net142),
    .X(_2921_));
 sky130_fd_sc_hd__nand2_2 _3140_ (.A(_2886_),
    .B(_2921_),
    .Y(_2922_));
 sky130_fd_sc_hd__nor3_4 _3141_ (.A(net146),
    .B(_2900_),
    .C(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__o21bai_2 _3142_ (.A1(_2873_),
    .A2(_2920_),
    .B1_N(_2923_),
    .Y(_2924_));
 sky130_fd_sc_hd__and3_1 _3143_ (.A(net151),
    .B(\z80.tv80s.i_tv80_core.IR[3] ),
    .C(_2899_),
    .X(_2925_));
 sky130_fd_sc_hd__o21ba_1 _3144_ (.A1(_2883_),
    .A2(_2903_),
    .B1_N(_2925_),
    .X(_2926_));
 sky130_fd_sc_hd__a21oi_1 _3145_ (.A1(_2893_),
    .A2(_2926_),
    .B1(_2910_),
    .Y(_2927_));
 sky130_fd_sc_hd__nor2_1 _3146_ (.A(net147),
    .B(_2876_),
    .Y(_2928_));
 sky130_fd_sc_hd__inv_2 _3147_ (.A(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__o21a_1 _3148_ (.A1(net148),
    .A2(_2876_),
    .B1(_2893_),
    .X(_2930_));
 sky130_fd_sc_hd__and2b_2 _3149_ (.A_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(_2931_));
 sky130_fd_sc_hd__nand2b_2 _3150_ (.A_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .Y(_2932_));
 sky130_fd_sc_hd__and2_1 _3151_ (.A(_2921_),
    .B(_2931_),
    .X(_2933_));
 sky130_fd_sc_hd__nand2_1 _3152_ (.A(_2921_),
    .B(_2931_),
    .Y(_2934_));
 sky130_fd_sc_hd__and2_2 _3153_ (.A(_2913_),
    .B(_2928_),
    .X(_2935_));
 sky130_fd_sc_hd__nand2_2 _3154_ (.A(_2913_),
    .B(_2928_),
    .Y(_2936_));
 sky130_fd_sc_hd__or2_1 _3155_ (.A(_2910_),
    .B(_2920_),
    .X(_2937_));
 sky130_fd_sc_hd__nand2_1 _3156_ (.A(_2936_),
    .B(_2937_),
    .Y(_2938_));
 sky130_fd_sc_hd__nor2_2 _3157_ (.A(_2869_),
    .B(_2900_),
    .Y(_2939_));
 sky130_fd_sc_hd__and2b_4 _3158_ (.A_N(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(_2940_));
 sky130_fd_sc_hd__nand2b_1 _3159_ (.A_N(\z80.tv80s.i_tv80_core.IR[7] ),
    .B(\z80.tv80s.i_tv80_core.IR[6] ),
    .Y(_2941_));
 sky130_fd_sc_hd__and3_2 _3160_ (.A(net151),
    .B(_2899_),
    .C(_2940_),
    .X(_2942_));
 sky130_fd_sc_hd__or2_4 _3161_ (.A(net151),
    .B(_2883_),
    .X(_2943_));
 sky130_fd_sc_hd__nor2_4 _3162_ (.A(net102),
    .B(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__and2_1 _3163_ (.A(net114),
    .B(_2944_),
    .X(_2945_));
 sky130_fd_sc_hd__nor2_2 _3164_ (.A(_2918_),
    .B(net102),
    .Y(_2946_));
 sky130_fd_sc_hd__or2_2 _3165_ (.A(_2918_),
    .B(net102),
    .X(_2947_));
 sky130_fd_sc_hd__nor2_2 _3166_ (.A(_2823_),
    .B(_2824_),
    .Y(_2948_));
 sky130_fd_sc_hd__nand2_4 _3167_ (.A(net145),
    .B(net139),
    .Y(_2949_));
 sky130_fd_sc_hd__or2_4 _3168_ (.A(_2821_),
    .B(_2874_),
    .X(_2950_));
 sky130_fd_sc_hd__nor2_2 _3169_ (.A(_2887_),
    .B(_2943_),
    .Y(_2951_));
 sky130_fd_sc_hd__a211o_1 _3170_ (.A1(_2885_),
    .A2(_2940_),
    .B1(_2951_),
    .C1(_2939_),
    .X(_2952_));
 sky130_fd_sc_hd__o21ai_1 _3171_ (.A1(net148),
    .A2(_2900_),
    .B1(_2920_),
    .Y(_2953_));
 sky130_fd_sc_hd__nor2_2 _3172_ (.A(net123),
    .B(net127),
    .Y(_2954_));
 sky130_fd_sc_hd__o31a_1 _3173_ (.A1(_2825_),
    .A2(_2885_),
    .A3(_2940_),
    .B1(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__a2bb2o_1 _3174_ (.A1_N(_2930_),
    .A2_N(_2934_),
    .B1(_2913_),
    .B2(_2919_),
    .X(_2956_));
 sky130_fd_sc_hd__or3_1 _3175_ (.A(_2924_),
    .B(_2938_),
    .C(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__a31o_1 _3176_ (.A1(_2870_),
    .A2(_2931_),
    .A3(_2953_),
    .B1(_2952_),
    .X(_2958_));
 sky130_fd_sc_hd__or4_1 _3177_ (.A(_2927_),
    .B(_2955_),
    .C(_2957_),
    .D(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__nor3_4 _3178_ (.A(_2871_),
    .B(_2887_),
    .C(_2901_),
    .Y(_2960_));
 sky130_fd_sc_hd__nor2_1 _3179_ (.A(_2900_),
    .B(_2905_),
    .Y(_2961_));
 sky130_fd_sc_hd__or2_1 _3180_ (.A(_2900_),
    .B(_2905_),
    .X(_2962_));
 sky130_fd_sc_hd__a2bb2o_1 _3181_ (.A1_N(_2873_),
    .A2_N(_2926_),
    .B1(_2961_),
    .B2(_2879_),
    .X(_2963_));
 sky130_fd_sc_hd__nor2_4 _3182_ (.A(_2887_),
    .B(_2895_),
    .Y(_2964_));
 sky130_fd_sc_hd__and4b_1 _3183_ (.A_N(net155),
    .B(net156),
    .C(net152),
    .D(net148),
    .X(_2965_));
 sky130_fd_sc_hd__and3_1 _3184_ (.A(_2868_),
    .B(_2870_),
    .C(_2965_),
    .X(_2966_));
 sky130_fd_sc_hd__nand2_1 _3185_ (.A(_2872_),
    .B(_2965_),
    .Y(_2967_));
 sky130_fd_sc_hd__nor2_1 _3186_ (.A(_2901_),
    .B(_2922_),
    .Y(_2968_));
 sky130_fd_sc_hd__and2_1 _3187_ (.A(_2877_),
    .B(_2913_),
    .X(_2969_));
 sky130_fd_sc_hd__or4_1 _3188_ (.A(_2964_),
    .B(_2966_),
    .C(_2968_),
    .D(_2969_),
    .X(_2970_));
 sky130_fd_sc_hd__or3_1 _3189_ (.A(_2960_),
    .B(_2963_),
    .C(_2970_),
    .X(_2971_));
 sky130_fd_sc_hd__or3_2 _3190_ (.A(_2823_),
    .B(_2824_),
    .C(_2869_),
    .X(_2972_));
 sky130_fd_sc_hd__o21ba_1 _3191_ (.A1(_2919_),
    .A2(_2925_),
    .B1_N(_2972_),
    .X(_2973_));
 sky130_fd_sc_hd__nor4_4 _3192_ (.A(net148),
    .B(_2871_),
    .C(_2887_),
    .D(_2900_),
    .Y(_2974_));
 sky130_fd_sc_hd__nor2_2 _3193_ (.A(_2876_),
    .B(_2910_),
    .Y(_2975_));
 sky130_fd_sc_hd__nand2_1 _3194_ (.A(_2875_),
    .B(_2909_),
    .Y(_2976_));
 sky130_fd_sc_hd__nor2_2 _3195_ (.A(net146),
    .B(_2976_),
    .Y(_2977_));
 sky130_fd_sc_hd__or4_1 _3196_ (.A(_2971_),
    .B(_2973_),
    .C(_2974_),
    .D(_2977_),
    .X(_2978_));
 sky130_fd_sc_hd__or3_1 _3197_ (.A(_2916_),
    .B(_2959_),
    .C(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__nor2_2 _3198_ (.A(_2905_),
    .B(_2950_),
    .Y(_2980_));
 sky130_fd_sc_hd__nor2_2 _3199_ (.A(_2920_),
    .B(_2972_),
    .Y(_2981_));
 sky130_fd_sc_hd__or2_1 _3200_ (.A(_2878_),
    .B(_2981_),
    .X(_2982_));
 sky130_fd_sc_hd__nor2_1 _3201_ (.A(_2876_),
    .B(_2972_),
    .Y(_2983_));
 sky130_fd_sc_hd__or2_1 _3202_ (.A(_2982_),
    .B(_2983_),
    .X(_2984_));
 sky130_fd_sc_hd__or2_1 _3203_ (.A(_2980_),
    .B(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__nor2_1 _3204_ (.A(_2869_),
    .B(_2950_),
    .Y(_2986_));
 sky130_fd_sc_hd__or2_1 _3205_ (.A(_2869_),
    .B(_2950_),
    .X(_2987_));
 sky130_fd_sc_hd__and2_1 _3206_ (.A(_2872_),
    .B(_2928_),
    .X(_2988_));
 sky130_fd_sc_hd__a211o_1 _3207_ (.A1(net146),
    .A2(_2975_),
    .B1(_2986_),
    .C1(_2988_),
    .X(_2989_));
 sky130_fd_sc_hd__a211o_1 _3208_ (.A1(_2876_),
    .A2(_2900_),
    .B1(_2906_),
    .C1(net148),
    .X(_2990_));
 sky130_fd_sc_hd__nand2_1 _3209_ (.A(_2824_),
    .B(_2886_),
    .Y(_2991_));
 sky130_fd_sc_hd__or2_4 _3210_ (.A(net150),
    .B(net144),
    .X(_2992_));
 sky130_fd_sc_hd__or2_1 _3211_ (.A(_2962_),
    .B(_2992_),
    .X(_2993_));
 sky130_fd_sc_hd__a32o_1 _3212_ (.A1(_2904_),
    .A2(_2930_),
    .A3(_2993_),
    .B1(_2991_),
    .B2(_2990_),
    .X(_2994_));
 sky130_fd_sc_hd__nand2_1 _3213_ (.A(net142),
    .B(_2883_),
    .Y(_2995_));
 sky130_fd_sc_hd__nand3b_4 _3214_ (.A_N(\z80.tv80s.i_tv80_core.IR[6] ),
    .B(\z80.tv80s.i_tv80_core.IR[7] ),
    .C(net140),
    .Y(_2996_));
 sky130_fd_sc_hd__or4_1 _3215_ (.A(_2821_),
    .B(net147),
    .C(_2995_),
    .D(_2996_),
    .X(_2997_));
 sky130_fd_sc_hd__and3_1 _3216_ (.A(_2870_),
    .B(_2896_),
    .C(_2931_),
    .X(_2998_));
 sky130_fd_sc_hd__a31o_1 _3217_ (.A1(net146),
    .A2(_2885_),
    .A3(_2933_),
    .B1(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__o22a_1 _3218_ (.A1(net156),
    .A2(_2893_),
    .B1(_2902_),
    .B2(_2874_),
    .X(_3000_));
 sky130_fd_sc_hd__or3_1 _3219_ (.A(net142),
    .B(_2996_),
    .C(_3000_),
    .X(_3001_));
 sky130_fd_sc_hd__or2_4 _3220_ (.A(_2900_),
    .B(_2996_),
    .X(_3002_));
 sky130_fd_sc_hd__or2_2 _3221_ (.A(_2894_),
    .B(_2996_),
    .X(_3003_));
 sky130_fd_sc_hd__or3_4 _3222_ (.A(net154),
    .B(net153),
    .C(_2996_),
    .X(_3004_));
 sky130_fd_sc_hd__nor2_1 _3223_ (.A(_2876_),
    .B(_2996_),
    .Y(_3005_));
 sky130_fd_sc_hd__or2_2 _3224_ (.A(_2943_),
    .B(_2996_),
    .X(_3006_));
 sky130_fd_sc_hd__or3b_4 _3225_ (.A(net153),
    .B(_2996_),
    .C_N(net154),
    .X(_3007_));
 sky130_fd_sc_hd__a21oi_2 _3226_ (.A1(_2876_),
    .A2(_2943_),
    .B1(_2996_),
    .Y(_3008_));
 sky130_fd_sc_hd__nor2_1 _3227_ (.A(net151),
    .B(_2996_),
    .Y(_3009_));
 sky130_fd_sc_hd__or4bb_1 _3228_ (.A(_2999_),
    .B(_3009_),
    .C_N(_3001_),
    .D_N(_2997_),
    .X(_3010_));
 sky130_fd_sc_hd__or4b_1 _3229_ (.A(_2985_),
    .B(_2989_),
    .C(_3010_),
    .D_N(_2994_),
    .X(_3011_));
 sky130_fd_sc_hd__o32a_1 _3230_ (.A1(net146),
    .A2(_2934_),
    .A3(_2950_),
    .B1(_2996_),
    .B2(net143),
    .X(_3012_));
 sky130_fd_sc_hd__a31oi_1 _3231_ (.A1(net156),
    .A2(net152),
    .A3(net114),
    .B1(_2925_),
    .Y(_3013_));
 sky130_fd_sc_hd__nand3_1 _3232_ (.A(_2874_),
    .B(_2896_),
    .C(_2933_),
    .Y(_3014_));
 sky130_fd_sc_hd__or4_1 _3233_ (.A(_2871_),
    .B(net88),
    .C(_2896_),
    .D(_2932_),
    .X(_3015_));
 sky130_fd_sc_hd__o41a_1 _3234_ (.A1(net114),
    .A2(net142),
    .A3(_2918_),
    .A4(_2996_),
    .B1(_3015_),
    .X(_3016_));
 sky130_fd_sc_hd__o311a_1 _3235_ (.A1(_2902_),
    .A2(_2995_),
    .A3(_2996_),
    .B1(_3014_),
    .C1(_3016_),
    .X(_3017_));
 sky130_fd_sc_hd__o21ai_1 _3236_ (.A1(_3012_),
    .A2(_3013_),
    .B1(_3017_),
    .Y(_3018_));
 sky130_fd_sc_hd__nor2_2 _3237_ (.A(_2914_),
    .B(_2920_),
    .Y(_3019_));
 sky130_fd_sc_hd__and3_2 _3238_ (.A(net143),
    .B(_2868_),
    .C(_2965_),
    .X(_3020_));
 sky130_fd_sc_hd__a21o_1 _3239_ (.A1(_2913_),
    .A2(_2965_),
    .B1(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__or2_1 _3240_ (.A(_3019_),
    .B(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__nor2_1 _3241_ (.A(_2950_),
    .B(_2991_),
    .Y(_3023_));
 sky130_fd_sc_hd__or2_1 _3242_ (.A(_3022_),
    .B(_3023_),
    .X(_3024_));
 sky130_fd_sc_hd__or2_2 _3243_ (.A(_2823_),
    .B(_2905_),
    .X(_3025_));
 sky130_fd_sc_hd__a41o_1 _3244_ (.A1(_2893_),
    .A2(_2901_),
    .A3(_2904_),
    .A4(_2929_),
    .B1(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__a2bb2o_1 _3245_ (.A1_N(_2908_),
    .A2_N(_2972_),
    .B1(_2925_),
    .B2(_2913_),
    .X(_3027_));
 sky130_fd_sc_hd__or4b_1 _3246_ (.A(_3018_),
    .B(_3024_),
    .C(_3027_),
    .D_N(_3026_),
    .X(_3028_));
 sky130_fd_sc_hd__or3_1 _3247_ (.A(_2979_),
    .B(_3011_),
    .C(_3028_),
    .X(_3029_));
 sky130_fd_sc_hd__a22oi_1 _3248_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .A2(_2892_),
    .B1(_3029_),
    .B2(net158),
    .Y(_3030_));
 sky130_fd_sc_hd__nor2_1 _3249_ (.A(net158),
    .B(net159),
    .Y(_3031_));
 sky130_fd_sc_hd__or2_4 _3250_ (.A(net158),
    .B(net159),
    .X(_0383_));
 sky130_fd_sc_hd__nor3_4 _3251_ (.A(_2912_),
    .B(net103),
    .C(_2950_),
    .Y(_0384_));
 sky130_fd_sc_hd__or3_2 _3252_ (.A(_2912_),
    .B(net103),
    .C(_2950_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _3253_ (.A(_3009_),
    .B(_0384_),
    .X(_0386_));
 sky130_fd_sc_hd__or3_2 _3254_ (.A(net154),
    .B(net153),
    .C(net102),
    .X(_0387_));
 sky130_fd_sc_hd__nor2_2 _3255_ (.A(_2876_),
    .B(net102),
    .Y(_0388_));
 sky130_fd_sc_hd__or2_1 _3256_ (.A(_2876_),
    .B(net102),
    .X(_0389_));
 sky130_fd_sc_hd__and4b_1 _3257_ (.A_N(_0386_),
    .B(_0387_),
    .C(_0389_),
    .D(_2947_),
    .X(_0390_));
 sky130_fd_sc_hd__nor2_4 _3258_ (.A(net124),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .Y(_0391_));
 sky130_fd_sc_hd__or2_4 _3259_ (.A(net124),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .X(_0392_));
 sky130_fd_sc_hd__a21oi_1 _3260_ (.A1(_0384_),
    .A2(_0391_),
    .B1(_0390_),
    .Y(_0393_));
 sky130_fd_sc_hd__nor2_2 _3261_ (.A(net124),
    .B(net127),
    .Y(_0394_));
 sky130_fd_sc_hd__or2_4 _3262_ (.A(net125),
    .B(net129),
    .X(_0395_));
 sky130_fd_sc_hd__nor2_1 _3263_ (.A(_3007_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__o221a_1 _3264_ (.A1(net128),
    .A2(_0387_),
    .B1(_0395_),
    .B2(_3007_),
    .C1(_2947_),
    .X(_0397_));
 sky130_fd_sc_hd__o221a_1 _3265_ (.A1(net128),
    .A2(_3003_),
    .B1(_0395_),
    .B2(_3002_),
    .C1(_0389_),
    .X(_0398_));
 sky130_fd_sc_hd__a31o_1 _3266_ (.A1(_0393_),
    .A2(_0397_),
    .A3(_0398_),
    .B1(_0383_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _3267_ (.A(_2881_),
    .B(net88),
    .Y(_0400_));
 sky130_fd_sc_hd__or2_1 _3268_ (.A(_2881_),
    .B(net88),
    .X(_0401_));
 sky130_fd_sc_hd__a41o_1 _3269_ (.A1(net131),
    .A2(_2940_),
    .A3(_0400_),
    .A4(_0401_),
    .B1(net111),
    .X(_0402_));
 sky130_fd_sc_hd__a21bo_1 _3270_ (.A1(_2877_),
    .A2(_2913_),
    .B1_N(_2937_),
    .X(_0403_));
 sky130_fd_sc_hd__nor2_1 _3271_ (.A(_2869_),
    .B(_2885_),
    .Y(_0404_));
 sky130_fd_sc_hd__nor2_1 _3272_ (.A(_2887_),
    .B(_2894_),
    .Y(_0405_));
 sky130_fd_sc_hd__or3_1 _3273_ (.A(_3020_),
    .B(_0404_),
    .C(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__or4_1 _3274_ (.A(_2923_),
    .B(_2960_),
    .C(_0403_),
    .D(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__nor2_1 _3275_ (.A(_2869_),
    .B(_2943_),
    .Y(_0408_));
 sky130_fd_sc_hd__or2_2 _3276_ (.A(_2988_),
    .B(_0408_),
    .X(_0409_));
 sky130_fd_sc_hd__or2_2 _3277_ (.A(_2961_),
    .B(_2968_),
    .X(_0410_));
 sky130_fd_sc_hd__nor2_4 _3278_ (.A(_2876_),
    .B(_2887_),
    .Y(_0411_));
 sky130_fd_sc_hd__a2111o_1 _3279_ (.A1(_2913_),
    .A2(_2965_),
    .B1(_3019_),
    .C1(_3023_),
    .D1(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__or4_1 _3280_ (.A(_0407_),
    .B(_0409_),
    .C(_0410_),
    .D(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__nor2_1 _3281_ (.A(_2985_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__and3b_2 _3282_ (.A_N(_2918_),
    .B(net114),
    .C(_2868_),
    .X(_0415_));
 sky130_fd_sc_hd__o2111ai_4 _3283_ (.A1(net154),
    .A2(net114),
    .B1(_2868_),
    .C1(net156),
    .D1(net153),
    .Y(_0416_));
 sky130_fd_sc_hd__nor2_2 _3284_ (.A(_2869_),
    .B(_2895_),
    .Y(_0417_));
 sky130_fd_sc_hd__or2_1 _3285_ (.A(_2869_),
    .B(_2895_),
    .X(_0418_));
 sky130_fd_sc_hd__o22a_2 _3286_ (.A1(_2869_),
    .A2(_2900_),
    .B1(_2920_),
    .B2(_2873_),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_1 _3287_ (.A(_0418_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__and3_1 _3288_ (.A(_0416_),
    .B(_0418_),
    .C(_0419_),
    .X(_0421_));
 sky130_fd_sc_hd__and3_2 _3289_ (.A(net151),
    .B(_2868_),
    .C(_2899_),
    .X(_0422_));
 sky130_fd_sc_hd__or3b_2 _3290_ (.A(_2821_),
    .B(_2869_),
    .C_N(_2899_),
    .X(_0423_));
 sky130_fd_sc_hd__nor2_1 _3291_ (.A(_2966_),
    .B(_0422_),
    .Y(_0424_));
 sky130_fd_sc_hd__and3b_2 _3292_ (.A_N(net155),
    .B(net152),
    .C(_2886_),
    .X(_0425_));
 sky130_fd_sc_hd__or3_4 _3293_ (.A(net155),
    .B(_2821_),
    .C(_2887_),
    .X(_0426_));
 sky130_fd_sc_hd__a21o_1 _3294_ (.A1(_2881_),
    .A2(_0395_),
    .B1(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__and4b_1 _3295_ (.A_N(net87),
    .B(_0421_),
    .C(_0424_),
    .D(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__a21o_1 _3296_ (.A1(net129),
    .A2(net88),
    .B1(_2932_),
    .X(_0429_));
 sky130_fd_sc_hd__and3_2 _3297_ (.A(net114),
    .B(net125),
    .C(_2948_),
    .X(_0430_));
 sky130_fd_sc_hd__o21a_1 _3298_ (.A1(_2889_),
    .A2(_0430_),
    .B1(_0429_),
    .X(_0431_));
 sky130_fd_sc_hd__and3_1 _3299_ (.A(_2936_),
    .B(net102),
    .C(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__nand2_2 _3300_ (.A(net139),
    .B(_2951_),
    .Y(_0433_));
 sky130_fd_sc_hd__nand2_2 _3301_ (.A(_2824_),
    .B(_2951_),
    .Y(_0434_));
 sky130_fd_sc_hd__o2111a_1 _3302_ (.A1(net130),
    .A2(_0434_),
    .B1(_0433_),
    .C1(_0432_),
    .D1(_2976_),
    .X(_0435_));
 sky130_fd_sc_hd__a31o_1 _3303_ (.A1(_0414_),
    .A2(_0428_),
    .A3(_0435_),
    .B1(_0402_),
    .X(_0436_));
 sky130_fd_sc_hd__and3_2 _3304_ (.A(_3030_),
    .B(_0399_),
    .C(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__inv_2 _3305_ (.A(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__or2_1 _3306_ (.A(_2867_),
    .B(_0437_),
    .X(_0439_));
 sky130_fd_sc_hd__nor2_1 _3307_ (.A(net129),
    .B(_3004_),
    .Y(_0440_));
 sky130_fd_sc_hd__or2_1 _3308_ (.A(net128),
    .B(_3004_),
    .X(_0441_));
 sky130_fd_sc_hd__a21oi_4 _3309_ (.A1(_2829_),
    .A2(_2830_),
    .B1(net125),
    .Y(_0442_));
 sky130_fd_sc_hd__a21o_1 _3310_ (.A1(_2829_),
    .A2(_2830_),
    .B1(net124),
    .X(_0443_));
 sky130_fd_sc_hd__o2111a_1 _3311_ (.A1(_0389_),
    .A2(_0442_),
    .B1(_0441_),
    .C1(_0397_),
    .D1(_0393_),
    .X(_0444_));
 sky130_fd_sc_hd__o21ai_1 _3312_ (.A1(net126),
    .A2(_2976_),
    .B1(_0414_),
    .Y(_0445_));
 sky130_fd_sc_hd__or2_1 _3313_ (.A(net142),
    .B(net129),
    .X(_0446_));
 sky130_fd_sc_hd__o21a_1 _3314_ (.A1(_0434_),
    .A2(_0446_),
    .B1(_0432_),
    .X(_0447_));
 sky130_fd_sc_hd__a21oi_1 _3315_ (.A1(net114),
    .A2(net126),
    .B1(_2829_),
    .Y(_0448_));
 sky130_fd_sc_hd__o22a_1 _3316_ (.A1(_2906_),
    .A2(_0442_),
    .B1(_0448_),
    .B2(_3025_),
    .X(_0449_));
 sky130_fd_sc_hd__a21o_1 _3317_ (.A1(_2922_),
    .A2(_0449_),
    .B1(_2943_),
    .X(_0450_));
 sky130_fd_sc_hd__and4b_1 _3318_ (.A_N(_0445_),
    .B(_0450_),
    .C(_0447_),
    .D(_0428_),
    .X(_0451_));
 sky130_fd_sc_hd__o221a_2 _3319_ (.A1(_0383_),
    .A2(_0444_),
    .B1(_0451_),
    .B2(_0402_),
    .C1(_3030_),
    .X(_0452_));
 sky130_fd_sc_hd__nor2_1 _3320_ (.A(_2867_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__nand2_1 _3321_ (.A(net148),
    .B(net143),
    .Y(_0454_));
 sky130_fd_sc_hd__nor2_1 _3322_ (.A(net140),
    .B(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__and4b_1 _3323_ (.A_N(net140),
    .B(net138),
    .C(net148),
    .D(net143),
    .X(_0456_));
 sky130_fd_sc_hd__nor4b_1 _3324_ (.A(net148),
    .B(net140),
    .C(net138),
    .D_N(net143),
    .Y(_0457_));
 sky130_fd_sc_hd__nand2_1 _3325_ (.A(net148),
    .B(_2823_),
    .Y(_0458_));
 sky130_fd_sc_hd__and3b_2 _3326_ (.A_N(net143),
    .B(net140),
    .C(net148),
    .X(_0459_));
 sky130_fd_sc_hd__nor2_1 _3327_ (.A(net148),
    .B(_2912_),
    .Y(_0460_));
 sky130_fd_sc_hd__nor4b_1 _3328_ (.A(net148),
    .B(net143),
    .C(\z80.tv80s.i_tv80_core.F[2] ),
    .D_N(net140),
    .Y(_0461_));
 sky130_fd_sc_hd__a2111o_1 _3329_ (.A1(\z80.tv80s.i_tv80_core.F[2] ),
    .A2(_0459_),
    .B1(_0461_),
    .C1(_0456_),
    .D1(_0457_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _3330_ (.A0(_2992_),
    .A1(_0458_),
    .S(\z80.tv80s.i_tv80_core.F[6] ),
    .X(_0463_));
 sky130_fd_sc_hd__nor3b_2 _3331_ (.A(net143),
    .B(net140),
    .C_N(net149),
    .Y(_0464_));
 sky130_fd_sc_hd__nor3_1 _3332_ (.A(net148),
    .B(net143),
    .C(net140),
    .Y(_0465_));
 sky130_fd_sc_hd__mux2_1 _3333_ (.A0(_0464_),
    .A1(_0465_),
    .S(_2828_),
    .X(_0466_));
 sky130_fd_sc_hd__and3_2 _3334_ (.A(net150),
    .B(net144),
    .C(net140),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _3335_ (.A0(_2881_),
    .A1(_0467_),
    .S(\z80.tv80s.i_tv80_core.F[7] ),
    .X(_0468_));
 sky130_fd_sc_hd__nor3_2 _3336_ (.A(_0462_),
    .B(_0466_),
    .C(_0468_),
    .Y(_0469_));
 sky130_fd_sc_hd__nand2_1 _3337_ (.A(net130),
    .B(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__o31a_1 _3338_ (.A1(_2869_),
    .A2(_2900_),
    .A3(_0470_),
    .B1(_0395_),
    .X(_0471_));
 sky130_fd_sc_hd__nor2_1 _3339_ (.A(_0421_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__or2_4 _3340_ (.A(net648),
    .B(\z80.tv80s.i_tv80_core.NMICycle ),
    .X(_0473_));
 sky130_fd_sc_hd__a21bo_1 _3341_ (.A1(_0395_),
    .A2(_0473_),
    .B1_N(_2974_),
    .X(_0474_));
 sky130_fd_sc_hd__o221a_1 _3342_ (.A1(net130),
    .A2(_0434_),
    .B1(_0442_),
    .B2(_2967_),
    .C1(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_2 _3343_ (.A(net127),
    .B(_2936_),
    .Y(_0476_));
 sky130_fd_sc_hd__nand2_2 _3344_ (.A(_2889_),
    .B(net102),
    .Y(_0477_));
 sky130_fd_sc_hd__or4b_1 _3345_ (.A(net111),
    .B(_2931_),
    .C(_0425_),
    .D_N(_0433_),
    .X(_0478_));
 sky130_fd_sc_hd__a311oi_1 _3346_ (.A1(_2830_),
    .A2(_0391_),
    .A3(_0476_),
    .B1(_0477_),
    .C1(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__o41a_2 _3347_ (.A1(_2829_),
    .A2(_0462_),
    .A3(_0466_),
    .A4(_0468_),
    .B1(_0442_),
    .X(_0480_));
 sky130_fd_sc_hd__o211a_1 _3348_ (.A1(_0423_),
    .A2(_0480_),
    .B1(_0479_),
    .C1(_0475_),
    .X(_0481_));
 sky130_fd_sc_hd__or3b_1 _3349_ (.A(_0445_),
    .B(_0472_),
    .C_N(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__nor2_2 _3350_ (.A(_2825_),
    .B(net129),
    .Y(_0483_));
 sky130_fd_sc_hd__nand2_4 _3351_ (.A(net124),
    .B(net113),
    .Y(_0484_));
 sky130_fd_sc_hd__a21oi_1 _3352_ (.A1(_3003_),
    .A2(_0483_),
    .B1(_3004_),
    .Y(_0485_));
 sky130_fd_sc_hd__or2_1 _3353_ (.A(_0384_),
    .B(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__nor2_1 _3354_ (.A(net128),
    .B(_2947_),
    .Y(_0487_));
 sky130_fd_sc_hd__o21a_1 _3355_ (.A1(_3005_),
    .A2(_0487_),
    .B1(_0484_),
    .X(_0488_));
 sky130_fd_sc_hd__a21oi_1 _3356_ (.A1(_3006_),
    .A2(_0387_),
    .B1(net128),
    .Y(_0489_));
 sky130_fd_sc_hd__or4_1 _3357_ (.A(net159),
    .B(_0388_),
    .C(_0486_),
    .D(_0488_),
    .X(_0490_));
 sky130_fd_sc_hd__o31a_1 _3358_ (.A1(_0390_),
    .A2(_0489_),
    .A3(_0490_),
    .B1(_0482_),
    .X(_0491_));
 sky130_fd_sc_hd__or3_4 _3359_ (.A(net158),
    .B(_2867_),
    .C(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__and2b_1 _3360_ (.A_N(_0453_),
    .B(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _3361_ (.A(_0439_),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__and2_1 _3362_ (.A(net128),
    .B(_2892_),
    .X(_0495_));
 sky130_fd_sc_hd__nor2_4 _3363_ (.A(net785),
    .B(net666),
    .Y(_0496_));
 sky130_fd_sc_hd__or2_1 _3364_ (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .B(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .X(_0497_));
 sky130_fd_sc_hd__nor2_2 _3365_ (.A(net878),
    .B(_0496_),
    .Y(_0498_));
 sky130_fd_sc_hd__o21ai_4 _3366_ (.A1(net57),
    .A2(_0495_),
    .B1(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__nand2_1 _3367_ (.A(_0416_),
    .B(_0419_),
    .Y(_0500_));
 sky130_fd_sc_hd__nor2_2 _3368_ (.A(_2906_),
    .B(_2943_),
    .Y(_0501_));
 sky130_fd_sc_hd__or2_1 _3369_ (.A(_2906_),
    .B(_2943_),
    .X(_0502_));
 sky130_fd_sc_hd__a31o_1 _3370_ (.A1(net142),
    .A2(_2868_),
    .A3(_2875_),
    .B1(_2980_),
    .X(_0503_));
 sky130_fd_sc_hd__or4_1 _3371_ (.A(_2878_),
    .B(_0409_),
    .C(_0501_),
    .D(_0503_),
    .X(_0504_));
 sky130_fd_sc_hd__or3_1 _3372_ (.A(_2960_),
    .B(_0403_),
    .C(_0417_),
    .X(_0505_));
 sky130_fd_sc_hd__or2_1 _3373_ (.A(_2931_),
    .B(_0404_),
    .X(_0506_));
 sky130_fd_sc_hd__and2_1 _3374_ (.A(_2912_),
    .B(_2951_),
    .X(_0507_));
 sky130_fd_sc_hd__or4_1 _3375_ (.A(_2964_),
    .B(_0477_),
    .C(_0506_),
    .D(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__or4_1 _3376_ (.A(_3024_),
    .B(_0504_),
    .C(_0505_),
    .D(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__nor2_1 _3377_ (.A(_0500_),
    .B(_0509_),
    .Y(_0510_));
 sky130_fd_sc_hd__nor2_4 _3378_ (.A(_2887_),
    .B(_2920_),
    .Y(_0511_));
 sky130_fd_sc_hd__or2_2 _3379_ (.A(_2887_),
    .B(_2920_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_8 _3380_ (.A(net126),
    .B(_2829_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_2 _3381_ (.A(_2825_),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .Y(_0514_));
 sky130_fd_sc_hd__o21a_1 _3382_ (.A1(_0469_),
    .A2(_0514_),
    .B1(net113),
    .X(_0515_));
 sky130_fd_sc_hd__and2_1 _3383_ (.A(_0422_),
    .B(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__nor2_1 _3384_ (.A(net128),
    .B(_0513_),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_1 _3385_ (.A(net113),
    .B(_0514_),
    .Y(_0518_));
 sky130_fd_sc_hd__or2_1 _3386_ (.A(_2966_),
    .B(_0410_),
    .X(_0519_));
 sky130_fd_sc_hd__or2_1 _3387_ (.A(_2923_),
    .B(_0519_),
    .X(_0520_));
 sky130_fd_sc_hd__a21oi_2 _3388_ (.A1(_2830_),
    .A2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .B1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .Y(_0521_));
 sky130_fd_sc_hd__o21ai_1 _3389_ (.A1(net124),
    .A2(_0521_),
    .B1(_0476_),
    .Y(_0522_));
 sky130_fd_sc_hd__a21oi_2 _3390_ (.A1(_0392_),
    .A2(_0473_),
    .B1(net128),
    .Y(_0523_));
 sky130_fd_sc_hd__inv_2 _3391_ (.A(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__o32ai_4 _3392_ (.A1(net130),
    .A2(_0426_),
    .A3(_0430_),
    .B1(_0512_),
    .B2(_0395_),
    .Y(_0525_));
 sky130_fd_sc_hd__a221o_1 _3393_ (.A1(_0517_),
    .A2(_0520_),
    .B1(_0523_),
    .B2(net87),
    .C1(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__or4_1 _3394_ (.A(_2981_),
    .B(_0411_),
    .C(_0516_),
    .D(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__o21ai_1 _3395_ (.A1(net127),
    .A2(_0510_),
    .B1(_0522_),
    .Y(_0528_));
 sky130_fd_sc_hd__o21ai_1 _3396_ (.A1(_0527_),
    .A2(_0528_),
    .B1(net159),
    .Y(_0529_));
 sky130_fd_sc_hd__and2_1 _3397_ (.A(net124),
    .B(_2954_),
    .X(_0530_));
 sky130_fd_sc_hd__and2_2 _3398_ (.A(net88),
    .B(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__or2_1 _3399_ (.A(net127),
    .B(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__or3b_1 _3400_ (.A(net127),
    .B(_0531_),
    .C_N(net158),
    .X(_0533_));
 sky130_fd_sc_hd__inv_2 _3401_ (.A(_0533_),
    .Y(_0534_));
 sky130_fd_sc_hd__and3b_2 _3402_ (.A_N(_2950_),
    .B(_2824_),
    .C(_2940_),
    .X(_0535_));
 sky130_fd_sc_hd__or2_1 _3403_ (.A(_2944_),
    .B(_0386_),
    .X(_0536_));
 sky130_fd_sc_hd__inv_2 _3404_ (.A(_0536_),
    .Y(_0537_));
 sky130_fd_sc_hd__nor2_1 _3405_ (.A(_0535_),
    .B(_0536_),
    .Y(_0538_));
 sky130_fd_sc_hd__a221oi_1 _3406_ (.A1(_2944_),
    .A2(_0394_),
    .B1(_0517_),
    .B2(_0384_),
    .C1(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__nor2_1 _3407_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .B(_2830_),
    .Y(_0540_));
 sky130_fd_sc_hd__and3_2 _3408_ (.A(_2825_),
    .B(_2829_),
    .C(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(_0541_));
 sky130_fd_sc_hd__nand2_4 _3409_ (.A(_2825_),
    .B(_0540_),
    .Y(_0542_));
 sky130_fd_sc_hd__nand2_1 _3410_ (.A(net113),
    .B(_0542_),
    .Y(_0543_));
 sky130_fd_sc_hd__a21oi_1 _3411_ (.A1(_3004_),
    .A2(_3006_),
    .B1(_0443_),
    .Y(_0544_));
 sky130_fd_sc_hd__nor2_2 _3412_ (.A(_0385_),
    .B(_0514_),
    .Y(_0545_));
 sky130_fd_sc_hd__a221o_1 _3413_ (.A1(_2944_),
    .A2(_0395_),
    .B1(_0541_),
    .B2(_3005_),
    .C1(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__or4_1 _3414_ (.A(net127),
    .B(_0535_),
    .C(_0544_),
    .D(_0546_),
    .X(_0547_));
 sky130_fd_sc_hd__or2_1 _3415_ (.A(_0383_),
    .B(_0547_),
    .X(_0548_));
 sky130_fd_sc_hd__a31o_1 _3416_ (.A1(_0529_),
    .A2(_0533_),
    .A3(_0548_),
    .B1(net123),
    .X(_0549_));
 sky130_fd_sc_hd__a21oi_1 _3417_ (.A1(_0426_),
    .A2(_0510_),
    .B1(net113),
    .Y(_0550_));
 sky130_fd_sc_hd__nor2_1 _3418_ (.A(_0423_),
    .B(_0515_),
    .Y(_0551_));
 sky130_fd_sc_hd__a2111o_1 _3419_ (.A1(_0425_),
    .A2(_0430_),
    .B1(_2935_),
    .C1(_2981_),
    .D1(_0411_),
    .X(_0552_));
 sky130_fd_sc_hd__a221o_1 _3420_ (.A1(_0395_),
    .A2(_0511_),
    .B1(_0524_),
    .B2(net87),
    .C1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__a2111o_1 _3421_ (.A1(_0518_),
    .A2(_0520_),
    .B1(_0550_),
    .C1(_0551_),
    .D1(_0553_),
    .X(_0554_));
 sky130_fd_sc_hd__a221o_1 _3422_ (.A1(net158),
    .A2(_0532_),
    .B1(_0547_),
    .B2(net99),
    .C1(net123),
    .X(_0555_));
 sky130_fd_sc_hd__a31oi_2 _3423_ (.A1(net159),
    .A2(_0522_),
    .A3(_0554_),
    .B1(_0555_),
    .Y(_0556_));
 sky130_fd_sc_hd__and2_1 _3424_ (.A(net131),
    .B(_0473_),
    .X(_0557_));
 sky130_fd_sc_hd__o21a_1 _3425_ (.A1(_0523_),
    .A2(_0557_),
    .B1(net87),
    .X(_0558_));
 sky130_fd_sc_hd__or3_1 _3426_ (.A(_2923_),
    .B(_0500_),
    .C(_0558_),
    .X(_0559_));
 sky130_fd_sc_hd__nand2_1 _3427_ (.A(_2936_),
    .B(_2967_),
    .Y(_0560_));
 sky130_fd_sc_hd__a221o_1 _3428_ (.A1(_0410_),
    .A2(_0513_),
    .B1(_0517_),
    .B2(_0560_),
    .C1(_0559_),
    .X(_0561_));
 sky130_fd_sc_hd__o21a_1 _3429_ (.A1(_0410_),
    .A2(_0509_),
    .B1(net113),
    .X(_0562_));
 sky130_fd_sc_hd__o41a_1 _3430_ (.A1(_0516_),
    .A2(_0525_),
    .A3(_0561_),
    .A4(_0562_),
    .B1(net159),
    .X(_0563_));
 sky130_fd_sc_hd__nor2_1 _3431_ (.A(_3005_),
    .B(_0535_),
    .Y(_0564_));
 sky130_fd_sc_hd__o311a_1 _3432_ (.A1(net127),
    .A2(_3006_),
    .A3(_0513_),
    .B1(_0564_),
    .C1(_0441_),
    .X(_0565_));
 sky130_fd_sc_hd__a221o_1 _3433_ (.A1(net127),
    .A2(_0538_),
    .B1(_0539_),
    .B2(_0565_),
    .C1(_0383_),
    .X(_0566_));
 sky130_fd_sc_hd__or4b_2 _3434_ (.A(net123),
    .B(_0534_),
    .C(_0563_),
    .D_N(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__inv_2 _3435_ (.A(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__and3_1 _3436_ (.A(net115),
    .B(_0556_),
    .C(_0567_),
    .X(_0569_));
 sky130_fd_sc_hd__a21o_1 _3437_ (.A1(net523),
    .A2(_0568_),
    .B1(_0569_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_1 _3438_ (.A0(net486),
    .A1(net481),
    .S(_0567_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_1 _3439_ (.A0(_0570_),
    .A1(_0571_),
    .S(_0549_),
    .X(_0572_));
 sky130_fd_sc_hd__inv_2 _3440_ (.A(_0572_),
    .Y(_0573_));
 sky130_fd_sc_hd__o41a_4 _3441_ (.A1(_2833_),
    .A2(_0549_),
    .A3(_0556_),
    .A4(_0568_),
    .B1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__inv_2 _3442_ (.A(net56),
    .Y(_0575_));
 sky130_fd_sc_hd__or2_1 _3443_ (.A(net567),
    .B(net56),
    .X(_0576_));
 sky130_fd_sc_hd__or2_1 _3444_ (.A(_0499_),
    .B(_0576_),
    .X(_0577_));
 sky130_fd_sc_hd__and2b_2 _3445_ (.A_N(net13),
    .B(net117),
    .X(_0578_));
 sky130_fd_sc_hd__a21o_2 _3446_ (.A1(net122),
    .A2(net567),
    .B1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__or4b_1 _3447_ (.A(net123),
    .B(_2890_),
    .C(_0579_),
    .D_N(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .X(_0580_));
 sky130_fd_sc_hd__nor2_1 _3448_ (.A(_0577_),
    .B(_0580_),
    .Y(_0581_));
 sky130_fd_sc_hd__or2_4 _3449_ (.A(_0577_),
    .B(_0578_),
    .X(_0582_));
 sky130_fd_sc_hd__a21o_1 _3450_ (.A1(net286),
    .A2(_0582_),
    .B1(_0581_),
    .X(_0008_));
 sky130_fd_sc_hd__or4_1 _3451_ (.A(net123),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .C(_2890_),
    .D(_0579_),
    .X(_0583_));
 sky130_fd_sc_hd__nor2_1 _3452_ (.A(_0577_),
    .B(_0583_),
    .Y(_0584_));
 sky130_fd_sc_hd__and2b_1 _3453_ (.A_N(net542),
    .B(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__and3_1 _3454_ (.A(_2830_),
    .B(_0391_),
    .C(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__a21o_1 _3455_ (.A1(net248),
    .A2(_0582_),
    .B1(_0586_),
    .X(_0009_));
 sky130_fd_sc_hd__a22o_1 _3456_ (.A1(net388),
    .A2(_0582_),
    .B1(_0584_),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(_0010_));
 sky130_fd_sc_hd__and3_1 _3457_ (.A(net640),
    .B(_2830_),
    .C(_0585_),
    .X(_0587_));
 sky130_fd_sc_hd__a21o_1 _3458_ (.A1(net264),
    .A2(_0582_),
    .B1(_0587_),
    .X(_0011_));
 sky130_fd_sc_hd__nand2_1 _3459_ (.A(net123),
    .B(_2891_),
    .Y(_0588_));
 sky130_fd_sc_hd__a211oi_2 _3460_ (.A1(net122),
    .A2(net567),
    .B1(_0582_),
    .C1(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__a21o_1 _3461_ (.A1(net408),
    .A2(_0582_),
    .B1(_0589_),
    .X(_0012_));
 sky130_fd_sc_hd__or4_1 _3462_ (.A(net248),
    .B(net388),
    .C(net264),
    .D(net408),
    .X(_0590_));
 sky130_fd_sc_hd__a221o_1 _3463_ (.A1(net542),
    .A2(_0584_),
    .B1(_0590_),
    .B2(_0582_),
    .C1(_0589_),
    .X(_0591_));
 sky130_fd_sc_hd__or3_1 _3464_ (.A(_0586_),
    .B(net641),
    .C(_0591_),
    .X(_0029_));
 sky130_fd_sc_hd__or2_1 _3465_ (.A(_0581_),
    .B(_0589_),
    .X(_0592_));
 sky130_fd_sc_hd__or2_1 _3466_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(net542),
    .X(_0593_));
 sky130_fd_sc_hd__or2_1 _3467_ (.A(net123),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .X(_0594_));
 sky130_fd_sc_hd__o41a_1 _3468_ (.A1(_2825_),
    .A2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .A3(_0593_),
    .A4(_0594_),
    .B1(_2891_),
    .X(_0595_));
 sky130_fd_sc_hd__nor3_1 _3469_ (.A(_0577_),
    .B(_0579_),
    .C(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__o41a_1 _3470_ (.A1(net286),
    .A2(net264),
    .A3(net408),
    .A4(net250),
    .B1(_0582_),
    .X(_0597_));
 sky130_fd_sc_hd__or4_1 _3471_ (.A(net641),
    .B(_0592_),
    .C(_0596_),
    .D(_0597_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_2 _3472_ (.A(net117),
    .B(net13),
    .X(_0598_));
 sky130_fd_sc_hd__nand2_8 _3473_ (.A(net117),
    .B(net13),
    .Y(_0599_));
 sky130_fd_sc_hd__nor2_1 _3474_ (.A(net122),
    .B(_0599_),
    .Y(_0600_));
 sky130_fd_sc_hd__o31a_1 _3475_ (.A1(net116),
    .A2(\z80.tv80s.i_tv80_core.ts[1] ),
    .A3(net117),
    .B1(net131),
    .X(_0601_));
 sky130_fd_sc_hd__o31ai_1 _3476_ (.A1(net116),
    .A2(\z80.tv80s.i_tv80_core.ts[1] ),
    .A3(net117),
    .B1(net131),
    .Y(_0602_));
 sky130_fd_sc_hd__a21o_2 _3477_ (.A1(_0599_),
    .A2(net96),
    .B1(net119),
    .X(_0603_));
 sky130_fd_sc_hd__o21bai_1 _3478_ (.A1(net845),
    .A2(net96),
    .B1_N(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__and2_1 _3479_ (.A(net161),
    .B(_3021_),
    .X(_0605_));
 sky130_fd_sc_hd__o211a_1 _3480_ (.A1(_2878_),
    .A2(_3020_),
    .B1(_2912_),
    .C1(net161),
    .X(_0606_));
 sky130_fd_sc_hd__or2_2 _3481_ (.A(_0605_),
    .B(_0606_),
    .X(_0607_));
 sky130_fd_sc_hd__and3_1 _3482_ (.A(net145),
    .B(net96),
    .C(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__and4_1 _3483_ (.A(_2878_),
    .B(_0600_),
    .C(net97),
    .D(_0607_),
    .X(_0609_));
 sky130_fd_sc_hd__or3_1 _3484_ (.A(net96),
    .B(_0604_),
    .C(_0609_),
    .X(_0610_));
 sky130_fd_sc_hd__inv_2 _3485_ (.A(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__and2b_1 _3486_ (.A_N(_3021_),
    .B(_0606_),
    .X(_0612_));
 sky130_fd_sc_hd__o21bai_1 _3487_ (.A1(_0610_),
    .A2(_0612_),
    .B1_N(_0604_),
    .Y(_0613_));
 sky130_fd_sc_hd__nor2_4 _3488_ (.A(net113),
    .B(_0599_),
    .Y(_0614_));
 sky130_fd_sc_hd__and3_1 _3489_ (.A(net128),
    .B(net107),
    .C(_0598_),
    .X(_0615_));
 sky130_fd_sc_hd__nand2_1 _3490_ (.A(net107),
    .B(_0614_),
    .Y(_0616_));
 sky130_fd_sc_hd__or4b_1 _3491_ (.A(net158),
    .B(net680),
    .C(net473),
    .D_N(_0607_),
    .X(_0617_));
 sky130_fd_sc_hd__a22o_1 _3492_ (.A1(net161),
    .A2(_0613_),
    .B1(_0615_),
    .B2(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__a31o_1 _3493_ (.A1(net161),
    .A2(_2912_),
    .A3(_3020_),
    .B1(_0618_),
    .X(_0000_));
 sky130_fd_sc_hd__or2_1 _3494_ (.A(\z80.tv80s.i_tv80_core.F[6] ),
    .B(_0458_),
    .X(_0619_));
 sky130_fd_sc_hd__o221a_1 _3495_ (.A1(_2828_),
    .A2(_2992_),
    .B1(_0454_),
    .B2(net138),
    .C1(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__nor2_1 _3496_ (.A(_2962_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__a31o_1 _3497_ (.A1(net138),
    .A2(_2879_),
    .A3(_2961_),
    .B1(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__o21ai_1 _3498_ (.A1(\z80.tv80s.i_tv80_core.IR[7] ),
    .A2(_2882_),
    .B1(net88),
    .Y(_0623_));
 sky130_fd_sc_hd__o311a_1 _3499_ (.A1(_2882_),
    .A2(net88),
    .A3(net102),
    .B1(_0434_),
    .C1(_0623_),
    .X(_0624_));
 sky130_fd_sc_hd__a21bo_1 _3500_ (.A1(net126),
    .A2(_0622_),
    .B1_N(_0624_),
    .X(_0625_));
 sky130_fd_sc_hd__nor2_1 _3501_ (.A(_0383_),
    .B(_0387_),
    .Y(_0626_));
 sky130_fd_sc_hd__nor2_1 _3502_ (.A(_2885_),
    .B(net103),
    .Y(_0627_));
 sky130_fd_sc_hd__a221o_1 _3503_ (.A1(net160),
    .A2(_0625_),
    .B1(_0627_),
    .B2(\z80.tv80s.i_tv80_core.ISet[2] ),
    .C1(_0626_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_1 _3504_ (.A0(net466),
    .A1(_0628_),
    .S(net107),
    .X(_0014_));
 sky130_fd_sc_hd__nand2_1 _3505_ (.A(_0605_),
    .B(_0615_),
    .Y(_0629_));
 sky130_fd_sc_hd__a2bb2o_1 _3506_ (.A1_N(_0606_),
    .A2_N(_0629_),
    .B1(_0616_),
    .B2(net680),
    .X(_0001_));
 sky130_fd_sc_hd__or4_1 _3507_ (.A(net286),
    .B(net388),
    .C(net408),
    .D(net254),
    .X(_0630_));
 sky130_fd_sc_hd__a221o_1 _3508_ (.A1(_0584_),
    .A2(net543),
    .B1(_0630_),
    .B2(_0582_),
    .C1(_0592_),
    .X(_0031_));
 sky130_fd_sc_hd__a21oi_1 _3509_ (.A1(_0469_),
    .A2(_0513_),
    .B1(_0423_),
    .Y(_0631_));
 sky130_fd_sc_hd__and3b_1 _3510_ (.A_N(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(_2974_),
    .C(\z80.tv80s.i_tv80_core.IntCycle ),
    .X(_0632_));
 sky130_fd_sc_hd__or4_1 _3511_ (.A(_0501_),
    .B(_0560_),
    .C(_0631_),
    .D(_0632_),
    .X(_0633_));
 sky130_fd_sc_hd__nand2_2 _3512_ (.A(net101),
    .B(_0388_),
    .Y(_0634_));
 sky130_fd_sc_hd__a21bo_1 _3513_ (.A1(net161),
    .A2(_0633_),
    .B1_N(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__mux2_1 _3514_ (.A0(net335),
    .A1(_0635_),
    .S(net107),
    .X(_0015_));
 sky130_fd_sc_hd__a32o_1 _3515_ (.A1(_0422_),
    .A2(_0469_),
    .A3(_0513_),
    .B1(_0470_),
    .B2(_2939_),
    .X(_0636_));
 sky130_fd_sc_hd__a21oi_1 _3516_ (.A1(_2889_),
    .A2(_0426_),
    .B1(_2882_),
    .Y(_0637_));
 sky130_fd_sc_hd__o211a_1 _3517_ (.A1(net138),
    .A2(_2880_),
    .B1(_0463_),
    .C1(net126),
    .X(_0638_));
 sky130_fd_sc_hd__a2bb2o_1 _3518_ (.A1_N(_2962_),
    .A2_N(_0638_),
    .B1(_2974_),
    .B2(\z80.tv80s.i_tv80_core.NMICycle ),
    .X(_0639_));
 sky130_fd_sc_hd__or4_1 _3519_ (.A(_2964_),
    .B(_0415_),
    .C(_0637_),
    .D(_0639_),
    .X(_0640_));
 sky130_fd_sc_hd__or4_1 _3520_ (.A(_2968_),
    .B(_0408_),
    .C(_0417_),
    .D(_0511_),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _3521_ (.A(_2924_),
    .B(_2977_),
    .C(_0640_),
    .D(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__o31a_1 _3522_ (.A1(_2989_),
    .A2(_0636_),
    .A3(_0642_),
    .B1(net160),
    .X(_0643_));
 sky130_fd_sc_hd__o21a_1 _3523_ (.A1(_2944_),
    .A2(_2946_),
    .B1(net100),
    .X(_0644_));
 sky130_fd_sc_hd__and3_1 _3524_ (.A(\z80.tv80s.i_tv80_core.ISet[2] ),
    .B(net88),
    .C(net102),
    .X(_0645_));
 sky130_fd_sc_hd__and4_1 _3525_ (.A(net148),
    .B(net143),
    .C(net162),
    .D(net138),
    .X(_0646_));
 sky130_fd_sc_hd__a311o_1 _3526_ (.A1(net125),
    .A2(_2961_),
    .A3(_0646_),
    .B1(_0645_),
    .C1(net122),
    .X(_0647_));
 sky130_fd_sc_hd__o32a_1 _3527_ (.A1(_0643_),
    .A2(_0644_),
    .A3(_0647_),
    .B1(net318),
    .B2(net107),
    .X(_0016_));
 sky130_fd_sc_hd__nor2_1 _3528_ (.A(net122),
    .B(_0383_),
    .Y(_0648_));
 sky130_fd_sc_hd__nand2_1 _3529_ (.A(net109),
    .B(net101),
    .Y(_0649_));
 sky130_fd_sc_hd__and4bb_1 _3530_ (.A_N(net122),
    .B_N(_0433_),
    .C(net142),
    .D(net160),
    .X(_0650_));
 sky130_fd_sc_hd__a221o_1 _3531_ (.A1(net122),
    .A2(net506),
    .B1(_0386_),
    .B2(_0648_),
    .C1(_0650_),
    .X(_0013_));
 sky130_fd_sc_hd__a21o_1 _3532_ (.A1(net250),
    .A2(_0582_),
    .B1(_0596_),
    .X(_0007_));
 sky130_fd_sc_hd__a22o_1 _3533_ (.A1(net254),
    .A2(_0582_),
    .B1(_0585_),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(_0006_));
 sky130_fd_sc_hd__or2_1 _3534_ (.A(_2883_),
    .B(_2902_),
    .X(_0651_));
 sky130_fd_sc_hd__or4_1 _3535_ (.A(_2823_),
    .B(\z80.tv80s.i_tv80_core.IR[5] ),
    .C(net103),
    .D(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__o41a_1 _3536_ (.A1(net147),
    .A2(net103),
    .A3(_2949_),
    .A4(_2950_),
    .B1(_0652_),
    .X(_0653_));
 sky130_fd_sc_hd__nand2_1 _3537_ (.A(_0454_),
    .B(_0627_),
    .Y(_0654_));
 sky130_fd_sc_hd__a21o_1 _3538_ (.A1(_0653_),
    .A2(_0654_),
    .B1(_0649_),
    .X(_0655_));
 sky130_fd_sc_hd__a32o_1 _3539_ (.A1(_2879_),
    .A2(_0627_),
    .A3(_0648_),
    .B1(_0655_),
    .B2(net412),
    .X(_0005_));
 sky130_fd_sc_hd__a2bb2o_1 _3540_ (.A1_N(_0649_),
    .A2_N(_0653_),
    .B1(_0655_),
    .B2(net576),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _3541_ (.A(net473),
    .B(_0616_),
    .X(_0003_));
 sky130_fd_sc_hd__a221o_1 _3542_ (.A1(_0611_),
    .A2(_0612_),
    .B1(_0616_),
    .B2(net158),
    .C1(_0609_),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_2 _3543_ (.A(net113),
    .B(_0513_),
    .Y(_0656_));
 sky130_fd_sc_hd__a21o_1 _3544_ (.A1(_3002_),
    .A2(_3007_),
    .B1(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__and2_1 _3545_ (.A(_0391_),
    .B(_0593_),
    .X(_0658_));
 sky130_fd_sc_hd__nor2_1 _3546_ (.A(net147),
    .B(_0389_),
    .Y(_0659_));
 sky130_fd_sc_hd__o31ai_1 _3547_ (.A1(_2894_),
    .A2(net102),
    .A3(_0484_),
    .B1(net99),
    .Y(_0660_));
 sky130_fd_sc_hd__a221oi_2 _3548_ (.A1(_0384_),
    .A2(_0541_),
    .B1(_0658_),
    .B2(_0659_),
    .C1(_0660_),
    .Y(_0661_));
 sky130_fd_sc_hd__nor2_1 _3549_ (.A(net146),
    .B(_0434_),
    .Y(_0662_));
 sky130_fd_sc_hd__a32o_1 _3550_ (.A1(_2823_),
    .A2(net124),
    .A3(_0662_),
    .B1(_0513_),
    .B2(_2977_),
    .X(_0663_));
 sky130_fd_sc_hd__or4_1 _3551_ (.A(net124),
    .B(net129),
    .C(_2936_),
    .D(_0521_),
    .X(_0664_));
 sky130_fd_sc_hd__o211a_1 _3552_ (.A1(_0394_),
    .A2(_0426_),
    .B1(_0637_),
    .C1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .X(_0665_));
 sky130_fd_sc_hd__nor2_4 _3553_ (.A(net129),
    .B(_0391_),
    .Y(_0666_));
 sky130_fd_sc_hd__a21bo_1 _3554_ (.A1(net87),
    .A2(_0473_),
    .B1_N(_0416_),
    .X(_0667_));
 sky130_fd_sc_hd__o21ai_1 _3555_ (.A1(net147),
    .A2(_0502_),
    .B1(_0424_),
    .Y(_0668_));
 sky130_fd_sc_hd__o22a_1 _3556_ (.A1(_2922_),
    .A2(_0484_),
    .B1(_0542_),
    .B2(_3025_),
    .X(_0669_));
 sky130_fd_sc_hd__o21ai_1 _3557_ (.A1(_2897_),
    .A2(_0669_),
    .B1(net102),
    .Y(_0670_));
 sky130_fd_sc_hd__a221o_1 _3558_ (.A1(_0666_),
    .A2(_0667_),
    .B1(_0668_),
    .B2(_0658_),
    .C1(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__or4b_1 _3559_ (.A(_0663_),
    .B(_0671_),
    .C(_0665_),
    .D_N(_0664_),
    .X(_0672_));
 sky130_fd_sc_hd__a21o_1 _3560_ (.A1(_2885_),
    .A2(_0430_),
    .B1(net102),
    .X(_0673_));
 sky130_fd_sc_hd__and3_1 _3561_ (.A(net159),
    .B(_0672_),
    .C(_0673_),
    .X(_0674_));
 sky130_fd_sc_hd__a31o_1 _3562_ (.A1(_2954_),
    .A2(_0513_),
    .A3(_0645_),
    .B1(net99),
    .X(_0675_));
 sky130_fd_sc_hd__a2bb2o_4 _3563_ (.A1_N(_0675_),
    .A2_N(_0674_),
    .B1(_0661_),
    .B2(_0657_),
    .X(net22));
 sky130_fd_sc_hd__inv_2 _3564_ (.A(net22),
    .Y(_0676_));
 sky130_fd_sc_hd__or2_2 _3565_ (.A(_0383_),
    .B(_0656_),
    .X(_0677_));
 sky130_fd_sc_hd__or3_1 _3566_ (.A(net153),
    .B(_2996_),
    .C(_0677_),
    .X(_0678_));
 sky130_fd_sc_hd__o21a_1 _3567_ (.A1(\z80.tv80s.i_tv80_core.F[2] ),
    .A2(_3004_),
    .B1(_2828_),
    .X(_0679_));
 sky130_fd_sc_hd__a31o_1 _3568_ (.A1(\z80.tv80s.i_tv80_core.F[2] ),
    .A2(_3003_),
    .A3(_3007_),
    .B1(_0679_),
    .X(_0680_));
 sky130_fd_sc_hd__a21oi_1 _3569_ (.A1(net145),
    .A2(_0680_),
    .B1(_0678_),
    .Y(_0028_));
 sky130_fd_sc_hd__a211o_1 _3570_ (.A1(_3002_),
    .A2(_3007_),
    .B1(_0542_),
    .C1(net127),
    .X(_0681_));
 sky130_fd_sc_hd__or3_1 _3571_ (.A(net127),
    .B(_3003_),
    .C(_0443_),
    .X(_0682_));
 sky130_fd_sc_hd__nand2_1 _3572_ (.A(_2944_),
    .B(_0392_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor2_1 _3573_ (.A(net114),
    .B(_0385_),
    .Y(_0684_));
 sky130_fd_sc_hd__nand2_1 _3574_ (.A(net124),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__a41o_1 _3575_ (.A1(_0681_),
    .A2(_0682_),
    .A3(_0683_),
    .A4(_0685_),
    .B1(net159),
    .X(_0686_));
 sky130_fd_sc_hd__a21oi_2 _3576_ (.A1(_0588_),
    .A2(_0686_),
    .B1(net158),
    .Y(_0687_));
 sky130_fd_sc_hd__nor2_1 _3577_ (.A(net768),
    .B(_0578_),
    .Y(_0688_));
 sky130_fd_sc_hd__a21o_2 _3578_ (.A1(net113),
    .A2(_2923_),
    .B1(_0410_),
    .X(_0689_));
 sky130_fd_sc_hd__nand2_4 _3579_ (.A(_0513_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__inv_2 _3580_ (.A(_0690_),
    .Y(_0691_));
 sky130_fd_sc_hd__nor2_4 _3581_ (.A(_0391_),
    .B(_0512_),
    .Y(_0692_));
 sky130_fd_sc_hd__o21a_1 _3582_ (.A1(_0691_),
    .A2(_0692_),
    .B1(net161),
    .X(_0693_));
 sky130_fd_sc_hd__or4_1 _3583_ (.A(_0676_),
    .B(_0687_),
    .C(_0688_),
    .D(_0693_),
    .X(_0694_));
 sky130_fd_sc_hd__or2_1 _3584_ (.A(net648),
    .B(_0688_),
    .X(_0695_));
 sky130_fd_sc_hd__mux2_1 _3585_ (.A0(_0694_),
    .A1(_0695_),
    .S(net131),
    .X(_0019_));
 sky130_fd_sc_hd__a21o_1 _3586_ (.A1(_3006_),
    .A2(_0387_),
    .B1(_0484_),
    .X(_0696_));
 sky130_fd_sc_hd__o31a_1 _3587_ (.A1(_2876_),
    .A2(_2996_),
    .A3(_0656_),
    .B1(_0696_),
    .X(_0697_));
 sky130_fd_sc_hd__nor2_1 _3588_ (.A(_2906_),
    .B(_2950_),
    .Y(_0698_));
 sky130_fd_sc_hd__a2111o_1 _3589_ (.A1(net140),
    .A2(_2964_),
    .B1(_2982_),
    .C1(_0507_),
    .D1(_0698_),
    .X(_0699_));
 sky130_fd_sc_hd__nor2_1 _3590_ (.A(_2950_),
    .B(_3025_),
    .Y(_0700_));
 sky130_fd_sc_hd__or4_1 _3591_ (.A(_2983_),
    .B(_3020_),
    .C(_0477_),
    .D(_0700_),
    .X(_0701_));
 sky130_fd_sc_hd__nor2_1 _3592_ (.A(_0412_),
    .B(_0701_),
    .Y(_0702_));
 sky130_fd_sc_hd__or4_1 _3593_ (.A(_2960_),
    .B(_2969_),
    .C(_0415_),
    .D(_0417_),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_1 _3594_ (.A(_2824_),
    .B(_2964_),
    .Y(_0704_));
 sky130_fd_sc_hd__and4bb_1 _3595_ (.A_N(_0699_),
    .B_N(_0703_),
    .C(_0704_),
    .D(_0502_),
    .X(_0705_));
 sky130_fd_sc_hd__and2_1 _3596_ (.A(_0702_),
    .B(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__inv_2 _3597_ (.A(_0706_),
    .Y(_0707_));
 sky130_fd_sc_hd__a21o_1 _3598_ (.A1(_2871_),
    .A2(_2939_),
    .B1(_0409_),
    .X(_0708_));
 sky130_fd_sc_hd__or3_1 _3599_ (.A(_2986_),
    .B(_0422_),
    .C(_0519_),
    .X(_0709_));
 sky130_fd_sc_hd__or4_1 _3600_ (.A(_2924_),
    .B(_2939_),
    .C(_0409_),
    .D(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__or2_1 _3601_ (.A(_2938_),
    .B(_0506_),
    .X(_0711_));
 sky130_fd_sc_hd__or4_1 _3602_ (.A(net111),
    .B(net87),
    .C(_0425_),
    .D(_0514_),
    .X(_0712_));
 sky130_fd_sc_hd__or4_1 _3603_ (.A(_0511_),
    .B(_0710_),
    .C(_0711_),
    .D(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__o22a_1 _3604_ (.A1(_0383_),
    .A2(_0697_),
    .B1(_0707_),
    .B2(_0713_),
    .X(_0714_));
 sky130_fd_sc_hd__or2_1 _3605_ (.A(net22),
    .B(_0688_),
    .X(_0715_));
 sky130_fd_sc_hd__nand2_1 _3606_ (.A(_0694_),
    .B(_0715_),
    .Y(_0716_));
 sky130_fd_sc_hd__a21o_1 _3607_ (.A1(_0694_),
    .A2(_0715_),
    .B1(_0714_),
    .X(_0717_));
 sky130_fd_sc_hd__o21ai_1 _3608_ (.A1(net768),
    .A2(_0578_),
    .B1(net648),
    .Y(_0718_));
 sky130_fd_sc_hd__mux2_2 _3609_ (.A0(_0717_),
    .A1(_0718_),
    .S(net131),
    .X(_0017_));
 sky130_fd_sc_hd__a21oi_1 _3610_ (.A1(_0714_),
    .A2(_0716_),
    .B1(net131),
    .Y(_0719_));
 sky130_fd_sc_hd__nand2_1 _3611_ (.A(net128),
    .B(_2831_),
    .Y(_0720_));
 sky130_fd_sc_hd__a31o_1 _3612_ (.A1(net131),
    .A2(_2831_),
    .A3(_0695_),
    .B1(_0719_),
    .X(_0018_));
 sky130_fd_sc_hd__or3b_4 _3613_ (.A(net111),
    .B(_0394_),
    .C_N(_2923_),
    .X(_0721_));
 sky130_fd_sc_hd__or4_1 _3614_ (.A(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .B(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .C(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .D(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .X(_0722_));
 sky130_fd_sc_hd__nor2_1 _3615_ (.A(net113),
    .B(_0722_),
    .Y(_0723_));
 sky130_fd_sc_hd__a221o_1 _3616_ (.A1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .A2(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .B1(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .C1(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__a221o_2 _3617_ (.A1(net125),
    .A2(net466),
    .B1(net335),
    .B2(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .C1(_0724_),
    .X(_0725_));
 sky130_fd_sc_hd__a41o_1 _3618_ (.A1(net126),
    .A2(net159),
    .A3(net574),
    .A4(_2923_),
    .B1(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__nor2_1 _3619_ (.A(net882),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__or2_2 _3620_ (.A(net123),
    .B(_0727_),
    .X(_0728_));
 sky130_fd_sc_hd__inv_2 _3621_ (.A(_0728_),
    .Y(_0729_));
 sky130_fd_sc_hd__or2_2 _3622_ (.A(_0576_),
    .B(_0578_),
    .X(_0730_));
 sky130_fd_sc_hd__inv_2 _3623_ (.A(_0730_),
    .Y(_0731_));
 sky130_fd_sc_hd__and2_2 _3624_ (.A(_0499_),
    .B(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__nand2_2 _3625_ (.A(_0729_),
    .B(_0732_),
    .Y(_0733_));
 sky130_fd_sc_hd__o211a_1 _3626_ (.A1(net34),
    .A2(_0614_),
    .B1(_0733_),
    .C1(_2833_),
    .X(_0032_));
 sky130_fd_sc_hd__nor2_1 _3627_ (.A(_0607_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__nor2_1 _3628_ (.A(net111),
    .B(_2972_),
    .Y(_0735_));
 sky130_fd_sc_hd__nand2_1 _3629_ (.A(_2877_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__and3_1 _3630_ (.A(net787),
    .B(\z80.tv80s.i_tv80_core.INT_s ),
    .C(_0736_),
    .X(_0737_));
 sky130_fd_sc_hd__nor2_1 _3631_ (.A(_2947_),
    .B(_0677_),
    .Y(_0738_));
 sky130_fd_sc_hd__or4b_1 _3632_ (.A(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .B(_2947_),
    .C(_0677_),
    .D_N(net117),
    .X(_0739_));
 sky130_fd_sc_hd__or3b_1 _3633_ (.A(_2831_),
    .B(_2929_),
    .C_N(_0735_),
    .X(_0740_));
 sky130_fd_sc_hd__nor2_1 _3634_ (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(_0736_),
    .Y(_0741_));
 sky130_fd_sc_hd__o21a_1 _3635_ (.A1(_0738_),
    .A2(_0741_),
    .B1(net639),
    .X(_0742_));
 sky130_fd_sc_hd__o21a_1 _3636_ (.A1(net484),
    .A2(_0737_),
    .B1(_0734_),
    .X(_0743_));
 sky130_fd_sc_hd__o21ba_1 _3637_ (.A1(net787),
    .A2(_0742_),
    .B1_N(_0743_),
    .X(_0744_));
 sky130_fd_sc_hd__and3_1 _3638_ (.A(_0739_),
    .B(_0740_),
    .C(net788),
    .X(_0026_));
 sky130_fd_sc_hd__or4b_1 _3639_ (.A(net484),
    .B(_0607_),
    .C(_0733_),
    .D_N(_0737_),
    .X(_0745_));
 sky130_fd_sc_hd__a31o_1 _3640_ (.A1(net639),
    .A2(_2877_),
    .A3(_0735_),
    .B1(net805),
    .X(_0746_));
 sky130_fd_sc_hd__and3_1 _3641_ (.A(_0740_),
    .B(_0745_),
    .C(_0746_),
    .X(_0027_));
 sky130_fd_sc_hd__and4_1 _3642_ (.A(net162),
    .B(_2881_),
    .C(_2884_),
    .D(_2940_),
    .X(_0747_));
 sky130_fd_sc_hd__or3b_1 _3643_ (.A(net56),
    .B(_0579_),
    .C_N(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__o21ai_1 _3644_ (.A1(net46),
    .A2(_0473_),
    .B1(_0748_),
    .Y(_0024_));
 sky130_fd_sc_hd__nor2_1 _3645_ (.A(net733),
    .B(_0714_),
    .Y(_0749_));
 sky130_fd_sc_hd__o21a_1 _3646_ (.A1(_0557_),
    .A2(_0749_),
    .B1(net56),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_2 _3647_ (.A0(\z80.normal_wr_n ),
    .A1(\z80.early_wr_n ),
    .S(net1),
    .X(net49));
 sky130_fd_sc_hd__mux2_2 _3648_ (.A0(\z80.normal_rd_n ),
    .A1(\z80.early_rd_n ),
    .S(net1),
    .X(net45));
 sky130_fd_sc_hd__mux2_1 _3649_ (.A0(\z80.normal_iorq_n ),
    .A1(\z80.early_iorq_n ),
    .S(net1),
    .X(net48));
 sky130_fd_sc_hd__mux2_1 _3650_ (.A0(\z80.normal_mreq_n ),
    .A1(\z80.early_mreq_n ),
    .S(net1),
    .X(net47));
 sky130_fd_sc_hd__a21o_2 _3651_ (.A1(_2831_),
    .A2(_0599_),
    .B1(net113),
    .X(_0033_));
 sky130_fd_sc_hd__or2_1 _3652_ (.A(net131),
    .B(_0715_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _3653_ (.A(net334),
    .B(net56),
    .X(_0022_));
 sky130_fd_sc_hd__or2_1 _3654_ (.A(_0395_),
    .B(_0521_),
    .X(_0750_));
 sky130_fd_sc_hd__a21oi_2 _3655_ (.A1(_2935_),
    .A2(_0750_),
    .B1(net111),
    .Y(_0751_));
 sky130_fd_sc_hd__and2_1 _3656_ (.A(net139),
    .B(_0411_),
    .X(_0752_));
 sky130_fd_sc_hd__and2_1 _3657_ (.A(_0422_),
    .B(_0480_),
    .X(_0753_));
 sky130_fd_sc_hd__nor2_1 _3658_ (.A(_0394_),
    .B(_0416_),
    .Y(_0754_));
 sky130_fd_sc_hd__a21o_1 _3659_ (.A1(_0422_),
    .A2(_0480_),
    .B1(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__a32o_2 _3660_ (.A1(_2974_),
    .A2(_0395_),
    .A3(_0473_),
    .B1(_0442_),
    .B2(_2966_),
    .X(_0756_));
 sky130_fd_sc_hd__or2_1 _3661_ (.A(_2935_),
    .B(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__a221o_1 _3662_ (.A1(_0422_),
    .A2(_0480_),
    .B1(_0666_),
    .B2(_0420_),
    .C1(_0754_),
    .X(_0758_));
 sky130_fd_sc_hd__o31a_1 _3663_ (.A1(_0752_),
    .A2(_0757_),
    .A3(_0758_),
    .B1(_0751_),
    .X(_0759_));
 sky130_fd_sc_hd__o21a_1 _3664_ (.A1(_2946_),
    .A2(_3005_),
    .B1(_0666_),
    .X(_0760_));
 sky130_fd_sc_hd__or2_1 _3665_ (.A(_3004_),
    .B(_0484_),
    .X(_0761_));
 sky130_fd_sc_hd__inv_2 _3666_ (.A(_0761_),
    .Y(_0762_));
 sky130_fd_sc_hd__o21ai_1 _3667_ (.A1(_3006_),
    .A2(_0656_),
    .B1(net99),
    .Y(_0763_));
 sky130_fd_sc_hd__or3_2 _3668_ (.A(_0760_),
    .B(_0762_),
    .C(_0763_),
    .X(_0764_));
 sky130_fd_sc_hd__o21a_1 _3669_ (.A1(net99),
    .A2(_0759_),
    .B1(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__o21ai_4 _3670_ (.A1(net99),
    .A2(_0759_),
    .B1(_0764_),
    .Y(_0766_));
 sky130_fd_sc_hd__a2bb2o_1 _3671_ (.A1_N(_3002_),
    .A2_N(_0656_),
    .B1(_0666_),
    .B2(_2946_),
    .X(_0767_));
 sky130_fd_sc_hd__a211o_1 _3672_ (.A1(net145),
    .A2(_0411_),
    .B1(_0757_),
    .C1(_0758_),
    .X(_0768_));
 sky130_fd_sc_hd__a22oi_4 _3673_ (.A1(net99),
    .A2(_0767_),
    .B1(_0768_),
    .B2(_0751_),
    .Y(_0769_));
 sky130_fd_sc_hd__nor2_1 _3674_ (.A(_0766_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__o31a_1 _3675_ (.A1(_0411_),
    .A2(_0757_),
    .A3(_0758_),
    .B1(_0751_),
    .X(_0771_));
 sky130_fd_sc_hd__a2111o_1 _3676_ (.A1(net154),
    .A2(net129),
    .B1(_2996_),
    .C1(_2820_),
    .D1(net151),
    .X(_0772_));
 sky130_fd_sc_hd__o21ai_1 _3677_ (.A1(_0394_),
    .A2(_0772_),
    .B1(_3002_),
    .Y(_0773_));
 sky130_fd_sc_hd__o21a_1 _3678_ (.A1(net127),
    .A2(_0392_),
    .B1(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__a211o_1 _3679_ (.A1(_2946_),
    .A2(_0666_),
    .B1(_0763_),
    .C1(_0774_),
    .X(_0775_));
 sky130_fd_sc_hd__o21a_1 _3680_ (.A1(net99),
    .A2(_0771_),
    .B1(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__o21ai_1 _3681_ (.A1(net128),
    .A2(_0598_),
    .B1(_0720_),
    .Y(_0777_));
 sky130_fd_sc_hd__or3b_2 _3682_ (.A(_0777_),
    .B(_0770_),
    .C_N(_0776_),
    .X(_0778_));
 sky130_fd_sc_hd__and3_2 _3683_ (.A(net161),
    .B(_2877_),
    .C(_2913_),
    .X(_0779_));
 sky130_fd_sc_hd__and3_1 _3684_ (.A(net159),
    .B(net115),
    .C(_2969_),
    .X(_0780_));
 sky130_fd_sc_hd__nand2_8 _3685_ (.A(net115),
    .B(_0779_),
    .Y(_0781_));
 sky130_fd_sc_hd__and3_2 _3686_ (.A(net159),
    .B(\z80.tv80s.i_tv80_core.ts[4] ),
    .C(_2969_),
    .X(_0782_));
 sky130_fd_sc_hd__nand2_1 _3687_ (.A(\z80.tv80s.i_tv80_core.ts[4] ),
    .B(_0779_),
    .Y(_0783_));
 sky130_fd_sc_hd__nand2_1 _3688_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net136),
    .Y(_0784_));
 sky130_fd_sc_hd__nand3_4 _3689_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(net136),
    .Y(_0785_));
 sky130_fd_sc_hd__or2_4 _3690_ (.A(_2832_),
    .B(net334),
    .X(_0786_));
 sky130_fd_sc_hd__nand2_1 _3691_ (.A(_2835_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__o31a_2 _3692_ (.A1(_2835_),
    .A2(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .A3(_0785_),
    .B1(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__and2_1 _3693_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .B(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .X(_0789_));
 sky130_fd_sc_hd__or3_1 _3694_ (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .B(_2856_),
    .C(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__or3b_1 _3695_ (.A(net892),
    .B(_0790_),
    .C_N(_0788_),
    .X(_0791_));
 sky130_fd_sc_hd__a41o_4 _3696_ (.A1(_0778_),
    .A2(_0781_),
    .A3(net83),
    .A4(_0791_),
    .B1(net119),
    .X(_0792_));
 sky130_fd_sc_hd__o2111a_4 _3697_ (.A1(net99),
    .A2(_0771_),
    .B1(_0775_),
    .C1(net115),
    .D1(net128),
    .X(_0793_));
 sky130_fd_sc_hd__o21a_1 _3698_ (.A1(net117),
    .A2(_0793_),
    .B1(_0496_),
    .X(_0794_));
 sky130_fd_sc_hd__o21ai_4 _3699_ (.A1(net117),
    .A2(_0793_),
    .B1(_0496_),
    .Y(_0795_));
 sky130_fd_sc_hd__or3_2 _3700_ (.A(net85),
    .B(_0782_),
    .C(_0794_),
    .X(_0796_));
 sky130_fd_sc_hd__a31o_1 _3701_ (.A1(_0781_),
    .A2(net83),
    .A3(_0795_),
    .B1(\z80.tv80s.i_tv80_core.Alternate ),
    .X(_0797_));
 sky130_fd_sc_hd__o211a_1 _3702_ (.A1(net117),
    .A2(_0793_),
    .B1(_0769_),
    .C1(_0765_),
    .X(_0798_));
 sky130_fd_sc_hd__o211ai_4 _3703_ (.A1(net117),
    .A2(_0793_),
    .B1(_0769_),
    .C1(_0765_),
    .Y(_0799_));
 sky130_fd_sc_hd__mux2_2 _3704_ (.A0(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .A1(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ),
    .S(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__o21a_4 _3705_ (.A1(_0796_),
    .A2(_0800_),
    .B1(_0797_),
    .X(_0801_));
 sky130_fd_sc_hd__o21ai_4 _3706_ (.A1(_0796_),
    .A2(_0800_),
    .B1(_0797_),
    .Y(_0802_));
 sky130_fd_sc_hd__a21o_1 _3707_ (.A1(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .A2(net83),
    .B1(net86),
    .X(_0803_));
 sky130_fd_sc_hd__o211ai_4 _3708_ (.A1(net117),
    .A2(_0793_),
    .B1(_0766_),
    .C1(_0496_),
    .Y(_0804_));
 sky130_fd_sc_hd__o31ai_4 _3709_ (.A1(_0794_),
    .A2(_0798_),
    .A3(_0803_),
    .B1(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__o31a_4 _3710_ (.A1(_0794_),
    .A2(_0798_),
    .A3(_0803_),
    .B1(_0804_),
    .X(_0806_));
 sky130_fd_sc_hd__o21ai_2 _3711_ (.A1(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .A2(_0782_),
    .B1(_0781_),
    .Y(_0807_));
 sky130_fd_sc_hd__o211a_2 _3712_ (.A1(net117),
    .A2(_0793_),
    .B1(_0769_),
    .C1(_0496_),
    .X(_0808_));
 sky130_fd_sc_hd__a31o_4 _3713_ (.A1(_0795_),
    .A2(_0799_),
    .A3(_0807_),
    .B1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__a31oi_4 _3714_ (.A1(_0795_),
    .A2(_0799_),
    .A3(_0807_),
    .B1(_0808_),
    .Y(_0810_));
 sky130_fd_sc_hd__and3_4 _3715_ (.A(_0802_),
    .B(_0806_),
    .C(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__or3_1 _3716_ (.A(_0801_),
    .B(_0805_),
    .C(_0809_),
    .X(_0812_));
 sky130_fd_sc_hd__or2_4 _3717_ (.A(_0792_),
    .B(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__nor2_4 _3718_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B(net86),
    .Y(_0814_));
 sky130_fd_sc_hd__or2_1 _3719_ (.A(\z80.tv80s.i_tv80_core.Alternate ),
    .B(net84),
    .X(_0815_));
 sky130_fd_sc_hd__o21a_1 _3720_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .A2(net86),
    .B1(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__o21ai_4 _3721_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .A2(net86),
    .B1(_0815_),
    .Y(_0817_));
 sky130_fd_sc_hd__mux4_1 _3722_ (.A0(net450),
    .A1(net396),
    .A2(net314),
    .A3(net355),
    .S0(net75),
    .S1(net72),
    .X(_0818_));
 sky130_fd_sc_hd__o211a_2 _3723_ (.A1(net128),
    .A2(net117),
    .B1(_0720_),
    .C1(_0776_),
    .X(_0819_));
 sky130_fd_sc_hd__inv_2 _3724_ (.A(net69),
    .Y(_0820_));
 sky130_fd_sc_hd__nor3_4 _3725_ (.A(net111),
    .B(net103),
    .C(_0401_),
    .Y(_0821_));
 sky130_fd_sc_hd__inv_4 _3726_ (.A(_0821_),
    .Y(_0822_));
 sky130_fd_sc_hd__and2_1 _3727_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0785_),
    .X(_0823_));
 sky130_fd_sc_hd__nand2_4 _3728_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_0785_),
    .Y(_0824_));
 sky130_fd_sc_hd__and2_2 _3729_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_2837_),
    .X(_0825_));
 sky130_fd_sc_hd__xnor2_1 _3730_ (.A(net137),
    .B(\z80.tv80s.i_tv80_core.BusB[0] ),
    .Y(_0826_));
 sky130_fd_sc_hd__a21o_1 _3731_ (.A1(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A2(\z80.tv80s.i_tv80_core.BusB[0] ),
    .B1(net137),
    .X(_0827_));
 sky130_fd_sc_hd__xnor2_1 _3732_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_0826_),
    .Y(_0828_));
 sky130_fd_sc_hd__and2b_1 _3733_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(net138),
    .X(_0829_));
 sky130_fd_sc_hd__nor2_1 _3734_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net136),
    .Y(_0830_));
 sky130_fd_sc_hd__xor2_1 _3735_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(net137),
    .X(_0831_));
 sky130_fd_sc_hd__mux2_1 _3736_ (.A0(net137),
    .A1(_0831_),
    .S(_0829_),
    .X(_0832_));
 sky130_fd_sc_hd__or2_1 _3737_ (.A(_0828_),
    .B(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__nand2_1 _3738_ (.A(_0828_),
    .B(_0832_),
    .Y(_0834_));
 sky130_fd_sc_hd__and2_1 _3739_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0784_),
    .X(_0835_));
 sky130_fd_sc_hd__nand2_4 _3740_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0784_),
    .Y(_0836_));
 sky130_fd_sc_hd__and3_2 _3741_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(_2838_),
    .X(_0837_));
 sky130_fd_sc_hd__a22o_1 _3742_ (.A1(_0825_),
    .A2(_0827_),
    .B1(_0828_),
    .B2(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__a31o_1 _3743_ (.A1(_0833_),
    .A2(_0834_),
    .A3(_0836_),
    .B1(_0838_),
    .X(_0839_));
 sky130_fd_sc_hd__o41a_2 _3744_ (.A1(_2838_),
    .A2(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A4(_0836_),
    .B1(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__and3b_1 _3745_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(net137),
    .C(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0841_));
 sky130_fd_sc_hd__and2_4 _3746_ (.A(_2837_),
    .B(_0841_),
    .X(_0842_));
 sky130_fd_sc_hd__nand2_1 _3747_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(_0841_),
    .Y(_0843_));
 sky130_fd_sc_hd__inv_2 _3748_ (.A(_0843_),
    .Y(_0844_));
 sky130_fd_sc_hd__o311a_1 _3749_ (.A1(net141),
    .A2(_2837_),
    .A3(_2992_),
    .B1(_0841_),
    .C1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_0845_));
 sky130_fd_sc_hd__and3b_4 _3750_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0830_),
    .C(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0846_));
 sky130_fd_sc_hd__or2_1 _3751_ (.A(net141),
    .B(net138),
    .X(_0847_));
 sky130_fd_sc_hd__a221o_1 _3752_ (.A1(net157),
    .A2(_2870_),
    .B1(_0847_),
    .B2(net143),
    .C1(net149),
    .X(_0848_));
 sky130_fd_sc_hd__o21a_1 _3753_ (.A1(_2822_),
    .A2(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B1(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__and4b_4 _3754_ (.A_N(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .C(_2838_),
    .D(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0850_));
 sky130_fd_sc_hd__or4_1 _3755_ (.A(_2836_),
    .B(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .C(_2837_),
    .D(net137),
    .X(_0851_));
 sky130_fd_sc_hd__a21o_1 _3756_ (.A1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A2(_0850_),
    .B1(_0842_),
    .X(_0852_));
 sky130_fd_sc_hd__nand2_2 _3757_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(_0830_),
    .Y(_0853_));
 sky130_fd_sc_hd__nor2_4 _3758_ (.A(_2836_),
    .B(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__or2_1 _3759_ (.A(_2836_),
    .B(_0853_),
    .X(_0855_));
 sky130_fd_sc_hd__and3b_4 _3760_ (.A_N(_0830_),
    .B(_0835_),
    .C(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_0856_));
 sky130_fd_sc_hd__inv_2 _3761_ (.A(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__mux2_1 _3762_ (.A0(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_0858_));
 sky130_fd_sc_hd__a22o_1 _3763_ (.A1(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A2(_0854_),
    .B1(_0856_),
    .B2(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__a221o_1 _3764_ (.A1(_0846_),
    .A2(_0849_),
    .B1(_0852_),
    .B2(_0465_),
    .C1(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__a2111o_1 _3765_ (.A1(_0824_),
    .A2(_0840_),
    .B1(_0845_),
    .C1(_0860_),
    .D1(_2835_),
    .X(_0861_));
 sky130_fd_sc_hd__o211a_1 _3766_ (.A1(net840),
    .A2(net854),
    .B1(_0822_),
    .C1(_0861_),
    .X(_0862_));
 sky130_fd_sc_hd__a21oi_4 _3767_ (.A1(net713),
    .A2(_0821_),
    .B1(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__o21ai_2 _3768_ (.A1(_0819_),
    .A2(_0863_),
    .B1(net83),
    .Y(_0864_));
 sky130_fd_sc_hd__and2_1 _3769_ (.A(net147),
    .B(_0411_),
    .X(_0865_));
 sky130_fd_sc_hd__or3b_2 _3770_ (.A(_0392_),
    .B(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .C_N(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(_0866_));
 sky130_fd_sc_hd__inv_2 _3771_ (.A(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__nor2_1 _3772_ (.A(net131),
    .B(_0866_),
    .Y(_0868_));
 sky130_fd_sc_hd__or2_1 _3773_ (.A(_2936_),
    .B(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__o311a_2 _3774_ (.A1(_0755_),
    .A2(_0757_),
    .A3(_0865_),
    .B1(_0869_),
    .C1(net159),
    .X(_0870_));
 sky130_fd_sc_hd__a21o_1 _3775_ (.A1(net147),
    .A2(_0392_),
    .B1(net127),
    .X(_0871_));
 sky130_fd_sc_hd__o211a_2 _3776_ (.A1(_0396_),
    .A2(_0773_),
    .B1(_0871_),
    .C1(net99),
    .X(_0872_));
 sky130_fd_sc_hd__nor2_8 _3777_ (.A(_0870_),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__inv_2 _3778_ (.A(_0873_),
    .Y(_0874_));
 sky130_fd_sc_hd__and3_4 _3779_ (.A(_0801_),
    .B(_0805_),
    .C(_0809_),
    .X(_0875_));
 sky130_fd_sc_hd__or3_4 _3780_ (.A(_0802_),
    .B(_0806_),
    .C(_0810_),
    .X(_0876_));
 sky130_fd_sc_hd__and3_4 _3781_ (.A(_0801_),
    .B(_0805_),
    .C(_0810_),
    .X(_0877_));
 sky130_fd_sc_hd__or3_4 _3782_ (.A(_0802_),
    .B(_0806_),
    .C(_0809_),
    .X(_0878_));
 sky130_fd_sc_hd__o22a_1 _3783_ (.A1(net355),
    .A2(_0876_),
    .B1(_0878_),
    .B2(net314),
    .X(_0879_));
 sky130_fd_sc_hd__and3_4 _3784_ (.A(_0802_),
    .B(_0805_),
    .C(_0809_),
    .X(_0880_));
 sky130_fd_sc_hd__or3_1 _3785_ (.A(_0801_),
    .B(_0806_),
    .C(_0810_),
    .X(_0881_));
 sky130_fd_sc_hd__and3_4 _3786_ (.A(_0802_),
    .B(_0805_),
    .C(_0810_),
    .X(_0882_));
 sky130_fd_sc_hd__or3_1 _3787_ (.A(_0801_),
    .B(_0806_),
    .C(_0809_),
    .X(_0883_));
 sky130_fd_sc_hd__o221a_1 _3788_ (.A1(net396),
    .A2(_0881_),
    .B1(_0883_),
    .B2(net450),
    .C1(_0879_),
    .X(_0884_));
 sky130_fd_sc_hd__and3_4 _3789_ (.A(_0801_),
    .B(_0806_),
    .C(_0809_),
    .X(_0885_));
 sky130_fd_sc_hd__or3_4 _3790_ (.A(_0802_),
    .B(_0805_),
    .C(_0810_),
    .X(_0886_));
 sky130_fd_sc_hd__and3_4 _3791_ (.A(_0802_),
    .B(_0806_),
    .C(_0809_),
    .X(_0887_));
 sky130_fd_sc_hd__or3_1 _3792_ (.A(_0801_),
    .B(_0805_),
    .C(_0810_),
    .X(_0888_));
 sky130_fd_sc_hd__o22a_1 _3793_ (.A1(net424),
    .A2(_0886_),
    .B1(_0888_),
    .B2(net509),
    .X(_0889_));
 sky130_fd_sc_hd__and3_4 _3794_ (.A(_0801_),
    .B(_0806_),
    .C(_0810_),
    .X(_0890_));
 sky130_fd_sc_hd__or3_4 _3795_ (.A(_0802_),
    .B(_0805_),
    .C(_0809_),
    .X(_0891_));
 sky130_fd_sc_hd__o221a_1 _3796_ (.A1(net515),
    .A2(_0812_),
    .B1(_0891_),
    .B2(net495),
    .C1(_0889_),
    .X(_0892_));
 sky130_fd_sc_hd__nand2_2 _3797_ (.A(_0884_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__xnor2_1 _3798_ (.A(net68),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__inv_2 _3799_ (.A(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__a22o_1 _3800_ (.A1(net288),
    .A2(_0875_),
    .B1(_0877_),
    .B2(net282),
    .X(_0896_));
 sky130_fd_sc_hd__a22o_1 _3801_ (.A1(net500),
    .A2(_0880_),
    .B1(_0882_),
    .B2(net458),
    .X(_0897_));
 sky130_fd_sc_hd__a22o_1 _3802_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .X(_0898_));
 sky130_fd_sc_hd__a221o_1 _3803_ (.A1(net493),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .C1(_0898_),
    .X(_0899_));
 sky130_fd_sc_hd__or3_2 _3804_ (.A(_0896_),
    .B(_0897_),
    .C(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__xnor2_1 _3805_ (.A(net68),
    .B(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__a22o_1 _3806_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .X(_0902_));
 sky130_fd_sc_hd__a221o_1 _3807_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(net353),
    .C1(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__a22o_1 _3808_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .X(_0904_));
 sky130_fd_sc_hd__a221o_1 _3809_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .C1(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__nor2_2 _3810_ (.A(_0903_),
    .B(_0905_),
    .Y(_0906_));
 sky130_fd_sc_hd__inv_2 _3811_ (.A(_0906_),
    .Y(_0907_));
 sky130_fd_sc_hd__xnor2_2 _3812_ (.A(_0873_),
    .B(_0906_),
    .Y(_0908_));
 sky130_fd_sc_hd__a22o_1 _3813_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .X(_0909_));
 sky130_fd_sc_hd__a221o_1 _3814_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .C1(_0909_),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _3815_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .X(_0911_));
 sky130_fd_sc_hd__a221o_1 _3816_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .C1(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__nor2_2 _3817_ (.A(_0910_),
    .B(_0912_),
    .Y(_0913_));
 sky130_fd_sc_hd__inv_2 _3818_ (.A(_0913_),
    .Y(_0914_));
 sky130_fd_sc_hd__xnor2_1 _3819_ (.A(_0873_),
    .B(_0913_),
    .Y(_0915_));
 sky130_fd_sc_hd__a22o_1 _3820_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .X(_0916_));
 sky130_fd_sc_hd__a221o_1 _3821_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .C1(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__a22o_1 _3822_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .X(_0918_));
 sky130_fd_sc_hd__a221o_1 _3823_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .C1(_0918_),
    .X(_0919_));
 sky130_fd_sc_hd__or2_2 _3824_ (.A(_0917_),
    .B(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__and2_1 _3825_ (.A(net68),
    .B(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__xnor2_1 _3826_ (.A(net68),
    .B(_0920_),
    .Y(_0922_));
 sky130_fd_sc_hd__a22o_1 _3827_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .X(_0923_));
 sky130_fd_sc_hd__a22o_1 _3828_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ),
    .X(_0924_));
 sky130_fd_sc_hd__a22o_1 _3829_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .X(_0925_));
 sky130_fd_sc_hd__a221o_1 _3830_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .C1(_0925_),
    .X(_0926_));
 sky130_fd_sc_hd__or3_4 _3831_ (.A(_0923_),
    .B(_0924_),
    .C(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__nand2_1 _3832_ (.A(net68),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__mux2_1 _3833_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .S(_0810_),
    .X(_0929_));
 sky130_fd_sc_hd__nor2_1 _3834_ (.A(_0806_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__mux2_1 _3835_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .S(_0810_),
    .X(_0931_));
 sky130_fd_sc_hd__o21ai_1 _3836_ (.A1(_0805_),
    .A2(_0931_),
    .B1(_0801_),
    .Y(_0932_));
 sky130_fd_sc_hd__mux2_1 _3837_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .S(_0810_),
    .X(_0933_));
 sky130_fd_sc_hd__mux2_1 _3838_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .S(_0810_),
    .X(_0934_));
 sky130_fd_sc_hd__mux2_1 _3839_ (.A0(_0933_),
    .A1(_0934_),
    .S(_0806_),
    .X(_0935_));
 sky130_fd_sc_hd__o2bb2a_2 _3840_ (.A1_N(_0802_),
    .A2_N(_0935_),
    .B1(_0932_),
    .B2(_0930_),
    .X(_0936_));
 sky130_fd_sc_hd__inv_2 _3841_ (.A(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__or2_1 _3842_ (.A(_0873_),
    .B(_0936_),
    .X(_0938_));
 sky130_fd_sc_hd__a311o_1 _3843_ (.A1(_0795_),
    .A2(_0799_),
    .A3(_0807_),
    .B1(_0808_),
    .C1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .X(_0939_));
 sky130_fd_sc_hd__mux2_1 _3844_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .S(_0809_),
    .X(_0940_));
 sky130_fd_sc_hd__o211a_1 _3845_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .A2(_0810_),
    .B1(_0939_),
    .C1(_0805_),
    .X(_0941_));
 sky130_fd_sc_hd__a211o_1 _3846_ (.A1(_0806_),
    .A2(_0940_),
    .B1(_0941_),
    .C1(_0802_),
    .X(_0942_));
 sky130_fd_sc_hd__mux2_1 _3847_ (.A0(net284),
    .A1(net384),
    .S(_0809_),
    .X(_0943_));
 sky130_fd_sc_hd__or3_1 _3848_ (.A(_0801_),
    .B(_0806_),
    .C(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__mux2_1 _3849_ (.A0(net332),
    .A1(net456),
    .S(_0809_),
    .X(_0945_));
 sky130_fd_sc_hd__or3_1 _3850_ (.A(_0801_),
    .B(_0805_),
    .C(_0945_),
    .X(_0946_));
 sky130_fd_sc_hd__nand3_2 _3851_ (.A(_0942_),
    .B(_0944_),
    .C(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__nand4_1 _3852_ (.A(net68),
    .B(_0942_),
    .C(_0944_),
    .D(_0946_),
    .Y(_0948_));
 sky130_fd_sc_hd__a31oi_1 _3853_ (.A1(_0942_),
    .A2(_0944_),
    .A3(_0946_),
    .B1(net68),
    .Y(_0949_));
 sky130_fd_sc_hd__nand2_1 _3854_ (.A(_0873_),
    .B(_0947_),
    .Y(_0950_));
 sky130_fd_sc_hd__nand2_1 _3855_ (.A(_0948_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__mux2_1 _3856_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .S(_0809_),
    .X(_0952_));
 sky130_fd_sc_hd__mux2_1 _3857_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .S(_0809_),
    .X(_0953_));
 sky130_fd_sc_hd__a21o_1 _3858_ (.A1(_0806_),
    .A2(_0953_),
    .B1(_0801_),
    .X(_0954_));
 sky130_fd_sc_hd__a21oi_1 _3859_ (.A1(_0805_),
    .A2(_0952_),
    .B1(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__mux2_1 _3860_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .S(_0809_),
    .X(_0956_));
 sky130_fd_sc_hd__mux2_1 _3861_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .S(_0809_),
    .X(_0957_));
 sky130_fd_sc_hd__mux2_1 _3862_ (.A0(_0956_),
    .A1(_0957_),
    .S(_0806_),
    .X(_0958_));
 sky130_fd_sc_hd__nor2_1 _3863_ (.A(_0802_),
    .B(_0958_),
    .Y(_0959_));
 sky130_fd_sc_hd__or2_2 _3864_ (.A(_0955_),
    .B(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__o31a_1 _3865_ (.A1(_0949_),
    .A2(_0955_),
    .A3(_0959_),
    .B1(_0948_),
    .X(_0961_));
 sky130_fd_sc_hd__xnor2_1 _3866_ (.A(_0873_),
    .B(_0936_),
    .Y(_0962_));
 sky130_fd_sc_hd__or2_1 _3867_ (.A(_0961_),
    .B(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__nand2_1 _3868_ (.A(_0938_),
    .B(_0963_),
    .Y(_0964_));
 sky130_fd_sc_hd__o21bai_1 _3869_ (.A1(net68),
    .A2(_0927_),
    .B1_N(_0963_),
    .Y(_0965_));
 sky130_fd_sc_hd__nand3_1 _3870_ (.A(_0928_),
    .B(_0938_),
    .C(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__a31o_1 _3871_ (.A1(_0928_),
    .A2(_0938_),
    .A3(_0965_),
    .B1(_0922_),
    .X(_0967_));
 sky130_fd_sc_hd__nor2_1 _3872_ (.A(_0915_),
    .B(_0967_),
    .Y(_0968_));
 sky130_fd_sc_hd__or4_1 _3873_ (.A(_0901_),
    .B(_0908_),
    .C(_0915_),
    .D(_0967_),
    .X(_0969_));
 sky130_fd_sc_hd__o41ai_2 _3874_ (.A1(_0900_),
    .A2(_0907_),
    .A3(_0914_),
    .A4(_0920_),
    .B1(net68),
    .Y(_0970_));
 sky130_fd_sc_hd__a21oi_1 _3875_ (.A1(_0969_),
    .A2(_0970_),
    .B1(_0895_),
    .Y(_0971_));
 sky130_fd_sc_hd__a21o_1 _3876_ (.A1(_0969_),
    .A2(_0970_),
    .B1(_0895_),
    .X(_0972_));
 sky130_fd_sc_hd__and3_1 _3877_ (.A(_0895_),
    .B(_0969_),
    .C(_0970_),
    .X(_0973_));
 sky130_fd_sc_hd__nor2_1 _3878_ (.A(_0971_),
    .B(_0973_),
    .Y(_0974_));
 sky130_fd_sc_hd__a21o_1 _3879_ (.A1(net69),
    .A2(_0974_),
    .B1(_0864_),
    .X(_0975_));
 sky130_fd_sc_hd__a21oi_1 _3880_ (.A1(_2863_),
    .A2(_0782_),
    .B1(net86),
    .Y(_0976_));
 sky130_fd_sc_hd__a22o_2 _3881_ (.A1(net85),
    .A2(_0818_),
    .B1(_0975_),
    .B2(_0976_),
    .X(_0977_));
 sky130_fd_sc_hd__mux2_1 _3882_ (.A0(_0977_),
    .A1(net515),
    .S(_0813_),
    .X(_0041_));
 sky130_fd_sc_hd__xnor2_1 _3883_ (.A(net136),
    .B(\z80.tv80s.i_tv80_core.BusB[1] ),
    .Y(_0978_));
 sky130_fd_sc_hd__nor2_1 _3884_ (.A(_2839_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__or2_1 _3885_ (.A(net136),
    .B(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__nand2_1 _3886_ (.A(_2839_),
    .B(_0978_),
    .Y(_0981_));
 sky130_fd_sc_hd__and2b_1 _3887_ (.A_N(_0979_),
    .B(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__o21ai_1 _3888_ (.A1(_2841_),
    .A2(_0826_),
    .B1(_0834_),
    .Y(_0983_));
 sky130_fd_sc_hd__xor2_1 _3889_ (.A(_0982_),
    .B(_0983_),
    .X(_0984_));
 sky130_fd_sc_hd__a22o_1 _3890_ (.A1(_0825_),
    .A2(_0980_),
    .B1(_0982_),
    .B2(_0837_),
    .X(_0985_));
 sky130_fd_sc_hd__a21o_1 _3891_ (.A1(_0836_),
    .A2(_0984_),
    .B1(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__o41a_1 _3892_ (.A1(_2838_),
    .A2(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A4(_0836_),
    .B1(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__mux2_1 _3893_ (.A0(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_0988_));
 sky130_fd_sc_hd__mux2_1 _3894_ (.A0(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[2] ),
    .S(net149),
    .X(_0989_));
 sky130_fd_sc_hd__a22o_1 _3895_ (.A1(_0856_),
    .A2(_0988_),
    .B1(_0989_),
    .B2(_0846_),
    .X(_0990_));
 sky130_fd_sc_hd__mux2_1 _3896_ (.A0(_0844_),
    .A1(_0850_),
    .S(_0464_),
    .X(_0991_));
 sky130_fd_sc_hd__o21a_1 _3897_ (.A1(_0842_),
    .A2(_0991_),
    .B1(net592),
    .X(_0992_));
 sky130_fd_sc_hd__a211o_1 _3898_ (.A1(_0464_),
    .A2(_0842_),
    .B1(_0990_),
    .C1(_0992_),
    .X(_0993_));
 sky130_fd_sc_hd__o21a_1 _3899_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_0994_));
 sky130_fd_sc_hd__o21ai_2 _3900_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .Y(_0995_));
 sky130_fd_sc_hd__nor2_1 _3901_ (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .B(_0994_),
    .Y(_0996_));
 sky130_fd_sc_hd__or2_1 _3902_ (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B(\z80.tv80s.i_tv80_core.F[4] ),
    .X(_0997_));
 sky130_fd_sc_hd__mux2_1 _3903_ (.A0(_0996_),
    .A1(_0997_),
    .S(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(_0998_));
 sky130_fd_sc_hd__inv_2 _3904_ (.A(_0998_),
    .Y(_0999_));
 sky130_fd_sc_hd__a221o_1 _3905_ (.A1(_0824_),
    .A2(_0987_),
    .B1(_0999_),
    .B2(_0854_),
    .C1(_0993_),
    .X(_1000_));
 sky130_fd_sc_hd__mux2_1 _3906_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_1000_),
    .S(net896),
    .X(_1001_));
 sky130_fd_sc_hd__and2_1 _3907_ (.A(net592),
    .B(_0821_),
    .X(_1002_));
 sky130_fd_sc_hd__a21oi_4 _3908_ (.A1(_0822_),
    .A2(_1001_),
    .B1(_1002_),
    .Y(_1003_));
 sky130_fd_sc_hd__inv_2 _3909_ (.A(_1003_),
    .Y(_1004_));
 sky130_fd_sc_hd__o21ai_2 _3910_ (.A1(net69),
    .A2(_1003_),
    .B1(net83),
    .Y(_1005_));
 sky130_fd_sc_hd__a22o_1 _3911_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .X(_1006_));
 sky130_fd_sc_hd__a221o_1 _3912_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .C1(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__a22o_1 _3913_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .X(_1008_));
 sky130_fd_sc_hd__a221o_1 _3914_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .C1(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nor2_2 _3915_ (.A(_1007_),
    .B(_1009_),
    .Y(_1010_));
 sky130_fd_sc_hd__inv_2 _3916_ (.A(_1010_),
    .Y(_1011_));
 sky130_fd_sc_hd__xnor2_2 _3917_ (.A(_0873_),
    .B(_1010_),
    .Y(_1012_));
 sky130_fd_sc_hd__o21ai_1 _3918_ (.A1(_0873_),
    .A2(_0893_),
    .B1(_0972_),
    .Y(_1013_));
 sky130_fd_sc_hd__xnor2_1 _3919_ (.A(_1012_),
    .B(_1013_),
    .Y(_1014_));
 sky130_fd_sc_hd__a21o_1 _3920_ (.A1(net69),
    .A2(_1014_),
    .B1(_1005_),
    .X(_1015_));
 sky130_fd_sc_hd__o21a_1 _3921_ (.A1(net230),
    .A2(net82),
    .B1(net84),
    .X(_1016_));
 sky130_fd_sc_hd__mux4_1 _3922_ (.A0(net420),
    .A1(net268),
    .A2(net426),
    .A3(net343),
    .S0(net72),
    .S1(net75),
    .X(_1017_));
 sky130_fd_sc_hd__a22o_2 _3923_ (.A1(_1015_),
    .A2(_1016_),
    .B1(_1017_),
    .B2(net85),
    .X(_1018_));
 sky130_fd_sc_hd__mux2_1 _3924_ (.A0(_1018_),
    .A1(net422),
    .S(_0813_),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_1 _3925_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .X(_1019_));
 sky130_fd_sc_hd__a221o_1 _3926_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .C1(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__a22o_1 _3927_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .X(_1021_));
 sky130_fd_sc_hd__a221o_1 _3928_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .C1(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__or2_2 _3929_ (.A(_1020_),
    .B(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__xnor2_1 _3930_ (.A(net68),
    .B(_1023_),
    .Y(_1024_));
 sky130_fd_sc_hd__a21o_1 _3931_ (.A1(_0893_),
    .A2(_1010_),
    .B1(_0873_),
    .X(_1025_));
 sky130_fd_sc_hd__a21o_1 _3932_ (.A1(_0873_),
    .A2(_1010_),
    .B1(_0972_),
    .X(_1026_));
 sky130_fd_sc_hd__a21oi_1 _3933_ (.A1(_1025_),
    .A2(_1026_),
    .B1(_1024_),
    .Y(_1027_));
 sky130_fd_sc_hd__and3_1 _3934_ (.A(_1024_),
    .B(_1025_),
    .C(_1026_),
    .X(_1028_));
 sky130_fd_sc_hd__nor2_1 _3935_ (.A(_1027_),
    .B(_1028_),
    .Y(_1029_));
 sky130_fd_sc_hd__xnor2_1 _3936_ (.A(net137),
    .B(\z80.tv80s.i_tv80_core.BusB[2] ),
    .Y(_1030_));
 sky130_fd_sc_hd__nor2_1 _3937_ (.A(_2840_),
    .B(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__or2_1 _3938_ (.A(net137),
    .B(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__nand2_1 _3939_ (.A(_2840_),
    .B(_1030_),
    .Y(_1033_));
 sky130_fd_sc_hd__and2b_1 _3940_ (.A_N(_1031_),
    .B(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__a21o_1 _3941_ (.A1(_0982_),
    .A2(_0983_),
    .B1(_0979_),
    .X(_1035_));
 sky130_fd_sc_hd__xor2_1 _3942_ (.A(_1034_),
    .B(_1035_),
    .X(_1036_));
 sky130_fd_sc_hd__a22o_1 _3943_ (.A1(_0825_),
    .A2(_1032_),
    .B1(_1034_),
    .B2(_0837_),
    .X(_1037_));
 sky130_fd_sc_hd__a21oi_1 _3944_ (.A1(_0836_),
    .A2(_1036_),
    .B1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__a41o_1 _3945_ (.A1(net137),
    .A2(_2840_),
    .A3(_2846_),
    .A4(_0835_),
    .B1(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__mux2_1 _3946_ (.A0(\z80.tv80s.i_tv80_core.F[1] ),
    .A1(_2839_),
    .S(_0996_),
    .X(_1040_));
 sky130_fd_sc_hd__xor2_1 _3947_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(\z80.tv80s.i_tv80_core.BusA[2] ),
    .X(_1041_));
 sky130_fd_sc_hd__xnor2_2 _3948_ (.A(_1040_),
    .B(_1041_),
    .Y(_1042_));
 sky130_fd_sc_hd__mux2_1 _3949_ (.A0(\z80.tv80s.i_tv80_core.BusB[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[6] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_1043_));
 sky130_fd_sc_hd__mux2_1 _3950_ (.A0(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .S(net149),
    .X(_1044_));
 sky130_fd_sc_hd__a221o_1 _3951_ (.A1(_0856_),
    .A2(_1043_),
    .B1(_1044_),
    .B2(_0846_),
    .C1(_0824_),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_1 _3952_ (.A(net141),
    .B(_2880_),
    .Y(_1046_));
 sky130_fd_sc_hd__nor2_1 _3953_ (.A(_0843_),
    .B(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__a211o_1 _3954_ (.A1(_0850_),
    .A2(_1046_),
    .B1(_1047_),
    .C1(_0842_),
    .X(_1048_));
 sky130_fd_sc_hd__a22o_1 _3955_ (.A1(_0854_),
    .A2(_1042_),
    .B1(_1048_),
    .B2(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(_1049_));
 sky130_fd_sc_hd__a211o_1 _3956_ (.A1(_0842_),
    .A2(_1046_),
    .B1(_1049_),
    .C1(_1045_),
    .X(_1050_));
 sky130_fd_sc_hd__a21bo_1 _3957_ (.A1(_0824_),
    .A2(_1039_),
    .B1_N(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__mux2_1 _3958_ (.A0(_2853_),
    .A1(_1051_),
    .S(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1052_));
 sky130_fd_sc_hd__mux2_8 _3959_ (.A0(_2846_),
    .A1(_1052_),
    .S(_0822_),
    .X(_1053_));
 sky130_fd_sc_hd__inv_2 _3960_ (.A(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__o21ai_2 _3961_ (.A1(_0819_),
    .A2(_1053_),
    .B1(net83),
    .Y(_1055_));
 sky130_fd_sc_hd__a21o_1 _3962_ (.A1(net69),
    .A2(_1029_),
    .B1(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__o21a_1 _3963_ (.A1(net236),
    .A2(net82),
    .B1(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__mux4_1 _3964_ (.A0(net400),
    .A1(net280),
    .A2(net505),
    .A3(net326),
    .S0(net72),
    .S1(net76),
    .X(_1058_));
 sky130_fd_sc_hd__mux2_2 _3965_ (.A0(_1057_),
    .A1(_1058_),
    .S(net85),
    .X(_1059_));
 sky130_fd_sc_hd__mux2_1 _3966_ (.A0(_1059_),
    .A1(net392),
    .S(_0813_),
    .X(_0043_));
 sky130_fd_sc_hd__xnor2_1 _3967_ (.A(net136),
    .B(\z80.tv80s.i_tv80_core.BusB[3] ),
    .Y(_1060_));
 sky130_fd_sc_hd__nor2_1 _3968_ (.A(_2842_),
    .B(_1060_),
    .Y(_1061_));
 sky130_fd_sc_hd__or2_1 _3969_ (.A(net136),
    .B(_1061_),
    .X(_1062_));
 sky130_fd_sc_hd__nand2_1 _3970_ (.A(_2842_),
    .B(_1060_),
    .Y(_1063_));
 sky130_fd_sc_hd__and2b_1 _3971_ (.A_N(_1061_),
    .B(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__a21o_1 _3972_ (.A1(_1034_),
    .A2(_1035_),
    .B1(_1031_),
    .X(_1065_));
 sky130_fd_sc_hd__xor2_1 _3973_ (.A(_1064_),
    .B(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__a22o_1 _3974_ (.A1(_0825_),
    .A2(_1062_),
    .B1(_1064_),
    .B2(_0837_),
    .X(_1067_));
 sky130_fd_sc_hd__a21o_1 _3975_ (.A1(_0836_),
    .A2(_1066_),
    .B1(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__o41a_2 _3976_ (.A1(_2838_),
    .A2(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A4(_0836_),
    .B1(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__a21o_1 _3977_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .B1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_1070_));
 sky130_fd_sc_hd__a31oi_1 _3978_ (.A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A3(\z80.tv80s.i_tv80_core.BusA[3] ),
    .B1(_0996_),
    .Y(_1071_));
 sky130_fd_sc_hd__or3_1 _3979_ (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .B(\z80.tv80s.i_tv80_core.BusA[2] ),
    .C(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(_1072_));
 sky130_fd_sc_hd__a21o_1 _3980_ (.A1(_0995_),
    .A2(_1072_),
    .B1(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1073_));
 sky130_fd_sc_hd__nand2_1 _3981_ (.A(_0997_),
    .B(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__a31o_1 _3982_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1070_),
    .A3(_1071_),
    .B1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_1 _3983_ (.A0(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[7] ),
    .S(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(_1076_));
 sky130_fd_sc_hd__mux2_1 _3984_ (.A0(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .S(net149),
    .X(_1077_));
 sky130_fd_sc_hd__and2_1 _3985_ (.A(_0846_),
    .B(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__a2bb2o_1 _3986_ (.A1_N(_0855_),
    .A2_N(_1075_),
    .B1(_1076_),
    .B2(_0856_),
    .X(_1079_));
 sky130_fd_sc_hd__mux2_1 _3987_ (.A0(_0844_),
    .A1(_0850_),
    .S(_0455_),
    .X(_1080_));
 sky130_fd_sc_hd__or2_1 _3988_ (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .B(_0455_),
    .X(_1081_));
 sky130_fd_sc_hd__a221o_1 _3989_ (.A1(net656),
    .A2(_1080_),
    .B1(_1081_),
    .B2(_0842_),
    .C1(_1078_),
    .X(_1082_));
 sky130_fd_sc_hd__a211o_1 _3990_ (.A1(_0824_),
    .A2(_1069_),
    .B1(_1079_),
    .C1(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__mux2_1 _3991_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_1083_),
    .S(net895),
    .X(_1084_));
 sky130_fd_sc_hd__and2_1 _3992_ (.A(net656),
    .B(_0821_),
    .X(_1085_));
 sky130_fd_sc_hd__a21oi_4 _3993_ (.A1(_0822_),
    .A2(_1084_),
    .B1(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__inv_2 _3994_ (.A(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__o21ai_1 _3995_ (.A1(net69),
    .A2(_1086_),
    .B1(net82),
    .Y(_1088_));
 sky130_fd_sc_hd__a22o_1 _3996_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .X(_1089_));
 sky130_fd_sc_hd__a221o_1 _3997_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .C1(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__a22o_1 _3998_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .X(_1091_));
 sky130_fd_sc_hd__a221o_1 _3999_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .C1(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__or2_2 _4000_ (.A(_1090_),
    .B(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__xnor2_1 _4001_ (.A(net68),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__a21o_1 _4002_ (.A1(net68),
    .A2(_1023_),
    .B1(_1027_),
    .X(_1095_));
 sky130_fd_sc_hd__xnor2_1 _4003_ (.A(_1094_),
    .B(_1095_),
    .Y(_1096_));
 sky130_fd_sc_hd__a21o_1 _4004_ (.A1(net69),
    .A2(_1096_),
    .B1(_1088_),
    .X(_1097_));
 sky130_fd_sc_hd__o21a_1 _4005_ (.A1(net226),
    .A2(net82),
    .B1(net84),
    .X(_1098_));
 sky130_fd_sc_hd__mux4_2 _4006_ (.A0(net488),
    .A1(net324),
    .A2(net448),
    .A3(net380),
    .S0(net72),
    .S1(net76),
    .X(_1099_));
 sky130_fd_sc_hd__a22o_2 _4007_ (.A1(_1097_),
    .A2(_1098_),
    .B1(_1099_),
    .B2(net85),
    .X(_1100_));
 sky130_fd_sc_hd__mux2_1 _4008_ (.A0(_1100_),
    .A1(net497),
    .S(_0813_),
    .X(_0044_));
 sky130_fd_sc_hd__or2_1 _4009_ (.A(_1024_),
    .B(_1094_),
    .X(_1101_));
 sky130_fd_sc_hd__o21ai_1 _4010_ (.A1(_1023_),
    .A2(_1093_),
    .B1(net68),
    .Y(_1102_));
 sky130_fd_sc_hd__o21a_1 _4011_ (.A1(_1025_),
    .A2(_1101_),
    .B1(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__o31ai_4 _4012_ (.A1(_0972_),
    .A2(_1012_),
    .A3(_1101_),
    .B1(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__a22o_1 _4013_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .X(_1105_));
 sky130_fd_sc_hd__a221o_1 _4014_ (.A1(net429),
    .A2(_0880_),
    .B1(_0882_),
    .B2(net452),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__a22o_1 _4015_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .X(_1107_));
 sky130_fd_sc_hd__a221o_1 _4016_ (.A1(net441),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .C1(_1107_),
    .X(_1108_));
 sky130_fd_sc_hd__nor2_1 _4017_ (.A(_1106_),
    .B(_1108_),
    .Y(_1109_));
 sky130_fd_sc_hd__inv_2 _4018_ (.A(_1109_),
    .Y(_1110_));
 sky130_fd_sc_hd__nor2_1 _4019_ (.A(_0873_),
    .B(_1109_),
    .Y(_1111_));
 sky130_fd_sc_hd__nor2_1 _4020_ (.A(net68),
    .B(_1110_),
    .Y(_1112_));
 sky130_fd_sc_hd__nor2_1 _4021_ (.A(_1111_),
    .B(_1112_),
    .Y(_1113_));
 sky130_fd_sc_hd__xnor2_1 _4022_ (.A(_1104_),
    .B(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__nand2_1 _4023_ (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .B(\z80.tv80s.i_tv80_core.F[4] ),
    .Y(_1115_));
 sky130_fd_sc_hd__o22a_1 _4024_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_0995_),
    .B1(_1070_),
    .B2(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__xnor2_2 _4025_ (.A(_2843_),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__inv_2 _4026_ (.A(_1117_),
    .Y(_1118_));
 sky130_fd_sc_hd__mux2_1 _4027_ (.A0(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .S(net149),
    .X(_1119_));
 sky130_fd_sc_hd__nor2_1 _4028_ (.A(_2838_),
    .B(\z80.tv80s.i_tv80_core.BusB[4] ),
    .Y(_1120_));
 sky130_fd_sc_hd__nor2_1 _4029_ (.A(net136),
    .B(_2847_),
    .Y(_1121_));
 sky130_fd_sc_hd__o21ai_2 _4030_ (.A1(_1120_),
    .A2(_1121_),
    .B1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .Y(_1122_));
 sky130_fd_sc_hd__or3_1 _4031_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_1120_),
    .C(_1121_),
    .X(_1123_));
 sky130_fd_sc_hd__and2_1 _4032_ (.A(_1122_),
    .B(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__a21o_1 _4033_ (.A1(_1064_),
    .A2(_1065_),
    .B1(_1061_),
    .X(_1125_));
 sky130_fd_sc_hd__or2_1 _4034_ (.A(_1124_),
    .B(_1125_),
    .X(_1126_));
 sky130_fd_sc_hd__nand2_1 _4035_ (.A(_1124_),
    .B(_1125_),
    .Y(_1127_));
 sky130_fd_sc_hd__nand2_1 _4036_ (.A(_2838_),
    .B(_1122_),
    .Y(_1128_));
 sky130_fd_sc_hd__a22o_1 _4037_ (.A1(_0837_),
    .A2(_1124_),
    .B1(_1128_),
    .B2(_0825_),
    .X(_1129_));
 sky130_fd_sc_hd__a31oi_1 _4038_ (.A1(_0836_),
    .A2(_1126_),
    .A3(_1127_),
    .B1(_1129_),
    .Y(_1130_));
 sky130_fd_sc_hd__a31o_1 _4039_ (.A1(_2843_),
    .A2(_0835_),
    .A3(_1120_),
    .B1(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__nand2_1 _4040_ (.A(_0824_),
    .B(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__a221o_1 _4041_ (.A1(_0460_),
    .A2(_0842_),
    .B1(_0846_),
    .B2(_1119_),
    .C1(_0824_),
    .X(_1133_));
 sky130_fd_sc_hd__nor2_1 _4042_ (.A(_0460_),
    .B(_0843_),
    .Y(_1134_));
 sky130_fd_sc_hd__a211o_1 _4043_ (.A1(_0460_),
    .A2(_0850_),
    .B1(_1134_),
    .C1(_0842_),
    .X(_1135_));
 sky130_fd_sc_hd__a221o_1 _4044_ (.A1(\z80.tv80s.i_tv80_core.BusA[4] ),
    .A2(_0856_),
    .B1(_1135_),
    .B2(\z80.tv80s.i_tv80_core.BusB[4] ),
    .C1(_1133_),
    .X(_1136_));
 sky130_fd_sc_hd__a21o_1 _4045_ (.A1(_0854_),
    .A2(_1118_),
    .B1(_1136_),
    .X(_1137_));
 sky130_fd_sc_hd__and3_1 _4046_ (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .B(_1132_),
    .C(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__a21oi_1 _4047_ (.A1(_2835_),
    .A2(\z80.tv80s.di_reg[4] ),
    .B1(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__mux2_4 _4048_ (.A0(_2847_),
    .A1(_1139_),
    .S(_0822_),
    .X(_1140_));
 sky130_fd_sc_hd__inv_2 _4049_ (.A(_1140_),
    .Y(_1141_));
 sky130_fd_sc_hd__o21a_1 _4050_ (.A1(net69),
    .A2(_1140_),
    .B1(net82),
    .X(_1142_));
 sky130_fd_sc_hd__o21ai_1 _4051_ (.A1(_0820_),
    .A2(_1114_),
    .B1(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__o21a_1 _4052_ (.A1(net234),
    .A2(net82),
    .B1(net84),
    .X(_1144_));
 sky130_fd_sc_hd__mux4_2 _4053_ (.A0(net452),
    .A1(net294),
    .A2(net429),
    .A3(net337),
    .S0(net72),
    .S1(net76),
    .X(_1145_));
 sky130_fd_sc_hd__a22o_2 _4054_ (.A1(_1143_),
    .A2(_1144_),
    .B1(_1145_),
    .B2(net85),
    .X(_1146_));
 sky130_fd_sc_hd__mux2_1 _4055_ (.A0(_1146_),
    .A1(net441),
    .S(_0813_),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _4056_ (.A(net674),
    .B(_0821_),
    .X(_1147_));
 sky130_fd_sc_hd__xnor2_1 _4057_ (.A(net136),
    .B(\z80.tv80s.i_tv80_core.BusB[5] ),
    .Y(_1148_));
 sky130_fd_sc_hd__xnor2_1 _4058_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _4059_ (.A(_1122_),
    .B(_1127_),
    .Y(_1150_));
 sky130_fd_sc_hd__a21bo_1 _4060_ (.A1(_1122_),
    .A2(_1127_),
    .B1_N(_1149_),
    .X(_1151_));
 sky130_fd_sc_hd__or2_1 _4061_ (.A(_1149_),
    .B(_1150_),
    .X(_1152_));
 sky130_fd_sc_hd__a21o_1 _4062_ (.A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A2(\z80.tv80s.i_tv80_core.BusB[5] ),
    .B1(net136),
    .X(_1153_));
 sky130_fd_sc_hd__a22o_1 _4063_ (.A1(_0837_),
    .A2(_1149_),
    .B1(_1153_),
    .B2(_0825_),
    .X(_1154_));
 sky130_fd_sc_hd__a31o_1 _4064_ (.A1(_0836_),
    .A2(_1151_),
    .A3(_1152_),
    .B1(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__o41a_2 _4065_ (.A1(_2838_),
    .A2(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A4(_0836_),
    .B1(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__nor2_1 _4066_ (.A(_2843_),
    .B(_0995_),
    .Y(_1157_));
 sky130_fd_sc_hd__nor2_1 _4067_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1157_),
    .Y(_1158_));
 sky130_fd_sc_hd__o31a_1 _4068_ (.A1(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A3(_1157_),
    .B1(net157),
    .X(_1159_));
 sky130_fd_sc_hd__nor2_1 _4069_ (.A(net138),
    .B(_1159_),
    .Y(_1160_));
 sky130_fd_sc_hd__or2_2 _4070_ (.A(net138),
    .B(_1159_),
    .X(_1161_));
 sky130_fd_sc_hd__and3_1 _4071_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(\z80.tv80s.i_tv80_core.BusA[5] ),
    .C(_0994_),
    .X(_1162_));
 sky130_fd_sc_hd__or2_1 _4072_ (.A(_1158_),
    .B(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__or3_1 _4073_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(_0996_),
    .C(_1070_),
    .X(_1164_));
 sky130_fd_sc_hd__or2_1 _4074_ (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .B(_1164_),
    .X(_1165_));
 sky130_fd_sc_hd__xnor2_1 _4075_ (.A(_2844_),
    .B(_1164_),
    .Y(_1166_));
 sky130_fd_sc_hd__mux2_1 _4076_ (.A0(_1163_),
    .A1(_1166_),
    .S(\z80.tv80s.i_tv80_core.F[1] ),
    .X(_1167_));
 sky130_fd_sc_hd__xnor2_1 _4077_ (.A(_1161_),
    .B(_1167_),
    .Y(_1168_));
 sky130_fd_sc_hd__o2bb2a_1 _4078_ (.A1_N(_0854_),
    .A2_N(_1168_),
    .B1(_0857_),
    .B2(_2844_),
    .X(_1169_));
 sky130_fd_sc_hd__inv_2 _4079_ (.A(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__mux2_2 _4080_ (.A0(\z80.tv80s.i_tv80_core.BusA[4] ),
    .A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .S(net149),
    .X(_1171_));
 sky130_fd_sc_hd__mux2_1 _4081_ (.A0(_0844_),
    .A1(_0850_),
    .S(_0459_),
    .X(_1172_));
 sky130_fd_sc_hd__o21a_1 _4082_ (.A1(_0842_),
    .A2(_1172_),
    .B1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(_1173_));
 sky130_fd_sc_hd__a221o_1 _4083_ (.A1(_0459_),
    .A2(_0842_),
    .B1(_0846_),
    .B2(_1171_),
    .C1(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__a211o_1 _4084_ (.A1(_0824_),
    .A2(_1156_),
    .B1(_1170_),
    .C1(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_1 _4085_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1175_),
    .S(net895),
    .X(_1176_));
 sky130_fd_sc_hd__a21oi_4 _4086_ (.A1(_0822_),
    .A2(_1176_),
    .B1(_1147_),
    .Y(_1177_));
 sky130_fd_sc_hd__inv_2 _4087_ (.A(_1177_),
    .Y(_1178_));
 sky130_fd_sc_hd__o21ai_1 _4088_ (.A1(net69),
    .A2(_1177_),
    .B1(net82),
    .Y(_1179_));
 sky130_fd_sc_hd__a22o_1 _4089_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .X(_1180_));
 sky130_fd_sc_hd__a221o_1 _4090_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .C1(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__a22o_1 _4091_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .X(_1182_));
 sky130_fd_sc_hd__a221o_1 _4092_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .C1(_1182_),
    .X(_1183_));
 sky130_fd_sc_hd__nor2_2 _4093_ (.A(_1181_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__inv_2 _4094_ (.A(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__xnor2_1 _4095_ (.A(_0873_),
    .B(_1184_),
    .Y(_1186_));
 sky130_fd_sc_hd__inv_2 _4096_ (.A(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__a21oi_1 _4097_ (.A1(_1104_),
    .A2(_1113_),
    .B1(_1111_),
    .Y(_1188_));
 sky130_fd_sc_hd__xnor2_1 _4098_ (.A(_1187_),
    .B(_1188_),
    .Y(_1189_));
 sky130_fd_sc_hd__a21o_1 _4099_ (.A1(net69),
    .A2(_1189_),
    .B1(_1179_),
    .X(_1190_));
 sky130_fd_sc_hd__o21a_1 _4100_ (.A1(net244),
    .A2(net82),
    .B1(net84),
    .X(_1191_));
 sky130_fd_sc_hd__mux4_1 _4101_ (.A0(net302),
    .A1(net360),
    .A2(net320),
    .A3(net463),
    .S0(net72),
    .S1(net76),
    .X(_1192_));
 sky130_fd_sc_hd__a22o_2 _4102_ (.A1(_1190_),
    .A2(_1191_),
    .B1(_1192_),
    .B2(net85),
    .X(_1193_));
 sky130_fd_sc_hd__mux2_1 _4103_ (.A0(_1193_),
    .A1(net513),
    .S(_0813_),
    .X(_0046_));
 sky130_fd_sc_hd__a22o_1 _4104_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .X(_1194_));
 sky130_fd_sc_hd__a221o_1 _4105_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .C1(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__a22o_1 _4106_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .X(_1196_));
 sky130_fd_sc_hd__a221o_1 _4107_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .A2(_0811_),
    .B1(_0890_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .C1(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__nor2_1 _4108_ (.A(_1195_),
    .B(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__inv_2 _4109_ (.A(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__nor2_1 _4110_ (.A(_0873_),
    .B(_1198_),
    .Y(_1200_));
 sky130_fd_sc_hd__nor2_1 _4111_ (.A(net68),
    .B(_1199_),
    .Y(_1201_));
 sky130_fd_sc_hd__nor2_1 _4112_ (.A(_1200_),
    .B(_1201_),
    .Y(_1202_));
 sky130_fd_sc_hd__a21oi_1 _4113_ (.A1(_1109_),
    .A2(_1184_),
    .B1(_0873_),
    .Y(_1203_));
 sky130_fd_sc_hd__a31o_1 _4114_ (.A1(_1104_),
    .A2(_1113_),
    .A3(_1187_),
    .B1(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__xor2_1 _4115_ (.A(_1202_),
    .B(_1204_),
    .X(_1205_));
 sky130_fd_sc_hd__xnor2_1 _4116_ (.A(net136),
    .B(\z80.tv80s.i_tv80_core.BusB[6] ),
    .Y(_1206_));
 sky130_fd_sc_hd__nor2_1 _4117_ (.A(_2845_),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__nand2_1 _4118_ (.A(_2845_),
    .B(_1206_),
    .Y(_1208_));
 sky130_fd_sc_hd__and2b_1 _4119_ (.A_N(_1207_),
    .B(_1208_),
    .X(_1209_));
 sky130_fd_sc_hd__o21ai_1 _4120_ (.A1(_2844_),
    .A2(_1148_),
    .B1(_1151_),
    .Y(_1210_));
 sky130_fd_sc_hd__xor2_1 _4121_ (.A(_1209_),
    .B(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__or2_1 _4122_ (.A(net136),
    .B(_1207_),
    .X(_1212_));
 sky130_fd_sc_hd__a22o_1 _4123_ (.A1(_0837_),
    .A2(_1209_),
    .B1(_1212_),
    .B2(_0825_),
    .X(_1213_));
 sky130_fd_sc_hd__a21o_1 _4124_ (.A1(_0836_),
    .A2(_1211_),
    .B1(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__o41a_2 _4125_ (.A1(_2838_),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A3(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A4(_0836_),
    .B1(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__xnor2_1 _4126_ (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B(_1162_),
    .Y(_1216_));
 sky130_fd_sc_hd__a21o_1 _4127_ (.A1(_1161_),
    .A2(_1163_),
    .B1(_1216_),
    .X(_1217_));
 sky130_fd_sc_hd__nand2_1 _4128_ (.A(_1163_),
    .B(_1216_),
    .Y(_1218_));
 sky130_fd_sc_hd__o211a_1 _4129_ (.A1(_1160_),
    .A2(_1218_),
    .B1(_1217_),
    .C1(_2849_),
    .X(_1219_));
 sky130_fd_sc_hd__xnor2_1 _4130_ (.A(_2845_),
    .B(_1165_),
    .Y(_1220_));
 sky130_fd_sc_hd__or2_1 _4131_ (.A(_1160_),
    .B(_1166_),
    .X(_1221_));
 sky130_fd_sc_hd__xnor2_1 _4132_ (.A(_1220_),
    .B(_1221_),
    .Y(_1222_));
 sky130_fd_sc_hd__a21oi_2 _4133_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1222_),
    .B1(_1219_),
    .Y(_1223_));
 sky130_fd_sc_hd__nor2_1 _4134_ (.A(_2881_),
    .B(_0843_),
    .Y(_1224_));
 sky130_fd_sc_hd__mux2_1 _4135_ (.A0(\z80.tv80s.i_tv80_core.BusA[5] ),
    .A1(net157),
    .S(net149),
    .X(_1225_));
 sky130_fd_sc_hd__a221o_1 _4136_ (.A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A2(_0856_),
    .B1(_1225_),
    .B2(_0846_),
    .C1(_0824_),
    .X(_1226_));
 sky130_fd_sc_hd__a211o_1 _4137_ (.A1(_2881_),
    .A2(_0850_),
    .B1(_1224_),
    .C1(_0842_),
    .X(_1227_));
 sky130_fd_sc_hd__a22o_1 _4138_ (.A1(_2881_),
    .A2(_0842_),
    .B1(_1227_),
    .B2(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(_1228_));
 sky130_fd_sc_hd__a211o_1 _4139_ (.A1(_0854_),
    .A2(_1223_),
    .B1(_1226_),
    .C1(_1228_),
    .X(_1229_));
 sky130_fd_sc_hd__o211a_1 _4140_ (.A1(_0823_),
    .A2(_1215_),
    .B1(_1229_),
    .C1(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(_1230_));
 sky130_fd_sc_hd__a21oi_1 _4141_ (.A1(_2835_),
    .A2(\z80.tv80s.di_reg[6] ),
    .B1(_1230_),
    .Y(_1231_));
 sky130_fd_sc_hd__mux2_4 _4142_ (.A0(_2848_),
    .A1(_1231_),
    .S(_0822_),
    .X(_1232_));
 sky130_fd_sc_hd__inv_2 _4143_ (.A(_1232_),
    .Y(_1233_));
 sky130_fd_sc_hd__o21a_1 _4144_ (.A1(net69),
    .A2(_1232_),
    .B1(net82),
    .X(_1234_));
 sky130_fd_sc_hd__a21bo_1 _4145_ (.A1(net69),
    .A2(_1205_),
    .B1_N(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__o21a_1 _4146_ (.A1(net246),
    .A2(net82),
    .B1(net84),
    .X(_1236_));
 sky130_fd_sc_hd__mux4_1 _4147_ (.A0(net357),
    .A1(net296),
    .A2(net300),
    .A3(net316),
    .S0(net72),
    .S1(net75),
    .X(_1237_));
 sky130_fd_sc_hd__a22o_2 _4148_ (.A1(_1235_),
    .A2(_1236_),
    .B1(_1237_),
    .B2(net85),
    .X(_1238_));
 sky130_fd_sc_hd__mux2_1 _4149_ (.A0(_1238_),
    .A1(net414),
    .S(_0813_),
    .X(_0047_));
 sky130_fd_sc_hd__a21o_1 _4150_ (.A1(_1202_),
    .A2(_1204_),
    .B1(_1200_),
    .X(_1239_));
 sky130_fd_sc_hd__a22o_1 _4151_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .A2(_0880_),
    .B1(_0882_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .X(_1240_));
 sky130_fd_sc_hd__a221o_1 _4152_ (.A1(net351),
    .A2(_0875_),
    .B1(_0877_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .C1(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__a22o_1 _4153_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .A2(_0885_),
    .B1(_0887_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .X(_1242_));
 sky130_fd_sc_hd__a221o_1 _4154_ (.A1(net418),
    .A2(_0811_),
    .B1(_0890_),
    .B2(net382),
    .C1(_1242_),
    .X(_1243_));
 sky130_fd_sc_hd__or2_1 _4155_ (.A(_1241_),
    .B(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__xnor2_1 _4156_ (.A(_0874_),
    .B(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__xnor2_1 _4157_ (.A(_1239_),
    .B(_1245_),
    .Y(_1246_));
 sky130_fd_sc_hd__and2_1 _4158_ (.A(net678),
    .B(_0821_),
    .X(_1247_));
 sky130_fd_sc_hd__a21o_1 _4159_ (.A1(_1209_),
    .A2(_1210_),
    .B1(_1207_),
    .X(_1248_));
 sky130_fd_sc_hd__xor2_1 _4160_ (.A(net157),
    .B(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__xor2_1 _4161_ (.A(net136),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(_1250_));
 sky130_fd_sc_hd__or2_1 _4162_ (.A(_1249_),
    .B(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__nand2_1 _4163_ (.A(_1249_),
    .B(_1250_),
    .Y(_1252_));
 sky130_fd_sc_hd__or2_1 _4164_ (.A(net157),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(_1253_));
 sky130_fd_sc_hd__nand2_1 _4165_ (.A(net157),
    .B(\z80.tv80s.i_tv80_core.BusB[7] ),
    .Y(_1254_));
 sky130_fd_sc_hd__nand2_1 _4166_ (.A(_2838_),
    .B(_1254_),
    .Y(_1255_));
 sky130_fd_sc_hd__a32o_1 _4167_ (.A1(_0837_),
    .A2(_1253_),
    .A3(_1254_),
    .B1(_1255_),
    .B2(_0825_),
    .X(_1256_));
 sky130_fd_sc_hd__a31o_1 _4168_ (.A1(_0836_),
    .A2(_1251_),
    .A3(_1252_),
    .B1(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__o41a_2 _4169_ (.A1(_2838_),
    .A2(net157),
    .A3(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A4(_0836_),
    .B1(_1257_),
    .X(_1258_));
 sky130_fd_sc_hd__xor2_1 _4170_ (.A(net157),
    .B(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(_1259_));
 sky130_fd_sc_hd__mux2_1 _4171_ (.A0(net157),
    .A1(_1259_),
    .S(_1162_),
    .X(_1260_));
 sky130_fd_sc_hd__and3b_1 _4172_ (.A_N(_1260_),
    .B(_1218_),
    .C(_1161_),
    .X(_1261_));
 sky130_fd_sc_hd__a21boi_1 _4173_ (.A1(_1161_),
    .A2(_1218_),
    .B1_N(_1260_),
    .Y(_1262_));
 sky130_fd_sc_hd__or3_1 _4174_ (.A(net157),
    .B(\z80.tv80s.i_tv80_core.BusA[6] ),
    .C(_1165_),
    .X(_1263_));
 sky130_fd_sc_hd__o21ai_1 _4175_ (.A1(\z80.tv80s.i_tv80_core.BusA[6] ),
    .A2(_1165_),
    .B1(net157),
    .Y(_1264_));
 sky130_fd_sc_hd__nand2_1 _4176_ (.A(_1263_),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__nor2_1 _4177_ (.A(_1166_),
    .B(_1220_),
    .Y(_1266_));
 sky130_fd_sc_hd__nor2_1 _4178_ (.A(_1265_),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__or2_1 _4179_ (.A(_1160_),
    .B(_1266_),
    .X(_1268_));
 sky130_fd_sc_hd__a221o_1 _4180_ (.A1(_1161_),
    .A2(_1267_),
    .B1(_1268_),
    .B2(_1265_),
    .C1(_2849_),
    .X(_1269_));
 sky130_fd_sc_hd__o31a_1 _4181_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1261_),
    .A3(_1262_),
    .B1(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__a22o_1 _4182_ (.A1(net157),
    .A2(_0856_),
    .B1(_1270_),
    .B2(_0854_),
    .X(_1271_));
 sky130_fd_sc_hd__nor2_1 _4183_ (.A(_2822_),
    .B(_2841_),
    .Y(_1272_));
 sky130_fd_sc_hd__a22o_1 _4184_ (.A1(_2822_),
    .A2(\z80.tv80s.i_tv80_core.BusA[6] ),
    .B1(_2870_),
    .B2(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__a211o_1 _4185_ (.A1(net157),
    .A2(_0459_),
    .B1(_1273_),
    .C1(_0456_),
    .X(_1274_));
 sky130_fd_sc_hd__nand2_1 _4186_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .B(_0467_),
    .Y(_1275_));
 sky130_fd_sc_hd__o211a_1 _4187_ (.A1(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A2(_0467_),
    .B1(_0841_),
    .C1(_1275_),
    .X(_1276_));
 sky130_fd_sc_hd__and3_1 _4188_ (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .B(_0467_),
    .C(_0850_),
    .X(_1277_));
 sky130_fd_sc_hd__a211o_1 _4189_ (.A1(_0846_),
    .A2(_1274_),
    .B1(_1276_),
    .C1(_1277_),
    .X(_1278_));
 sky130_fd_sc_hd__a211o_1 _4190_ (.A1(_0824_),
    .A2(_1258_),
    .B1(_1271_),
    .C1(_1278_),
    .X(_1279_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1279_),
    .S(net893),
    .X(_1280_));
 sky130_fd_sc_hd__a21oi_4 _4192_ (.A1(_0822_),
    .A2(_1280_),
    .B1(_1247_),
    .Y(_1281_));
 sky130_fd_sc_hd__inv_2 _4193_ (.A(_1281_),
    .Y(_1282_));
 sky130_fd_sc_hd__o21ai_1 _4194_ (.A1(net69),
    .A2(_1281_),
    .B1(net83),
    .Y(_1283_));
 sky130_fd_sc_hd__a21o_1 _4195_ (.A1(_0819_),
    .A2(_1246_),
    .B1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__o21a_1 _4196_ (.A1(net242),
    .A2(net82),
    .B1(net84),
    .X(_1285_));
 sky130_fd_sc_hd__nand2_8 _4197_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(_0781_),
    .Y(_1286_));
 sky130_fd_sc_hd__or3_1 _4198_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .B(net134),
    .C(net85),
    .X(_1287_));
 sky130_fd_sc_hd__o211a_1 _4199_ (.A1(net390),
    .A2(net76),
    .B1(net73),
    .C1(_1287_),
    .X(_1288_));
 sky130_fd_sc_hd__mux2_1 _4200_ (.A0(net366),
    .A1(net339),
    .S(net76),
    .X(_1289_));
 sky130_fd_sc_hd__o221a_1 _4201_ (.A1(net386),
    .A2(net134),
    .B1(net76),
    .B2(net382),
    .C1(net72),
    .X(_1290_));
 sky130_fd_sc_hd__o221a_1 _4202_ (.A1(net503),
    .A2(net134),
    .B1(net76),
    .B2(net418),
    .C1(net71),
    .X(_1291_));
 sky130_fd_sc_hd__a221o_1 _4203_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .A2(net84),
    .B1(net71),
    .B2(_1289_),
    .C1(_1288_),
    .X(_1292_));
 sky130_fd_sc_hd__o31a_1 _4204_ (.A1(_1286_),
    .A2(_1290_),
    .A3(_1291_),
    .B1(_1292_),
    .X(_1293_));
 sky130_fd_sc_hd__a22o_2 _4205_ (.A1(_1284_),
    .A2(_1285_),
    .B1(_1293_),
    .B2(net85),
    .X(_1294_));
 sky130_fd_sc_hd__mux2_1 _4206_ (.A0(_1294_),
    .A1(net418),
    .S(_0813_),
    .X(_0048_));
 sky130_fd_sc_hd__a32o_1 _4207_ (.A1(net125),
    .A2(_2882_),
    .A3(_2888_),
    .B1(_0417_),
    .B2(_0666_),
    .X(_1295_));
 sky130_fd_sc_hd__nor2_1 _4208_ (.A(_2882_),
    .B(_0483_),
    .Y(_1296_));
 sky130_fd_sc_hd__nor2_1 _4209_ (.A(_0426_),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__nand2_1 _4210_ (.A(_2825_),
    .B(net88),
    .Y(_1298_));
 sky130_fd_sc_hd__and3_1 _4211_ (.A(_2882_),
    .B(_2940_),
    .C(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__o31a_1 _4212_ (.A1(_1295_),
    .A2(_1297_),
    .A3(_1299_),
    .B1(net142),
    .X(_1300_));
 sky130_fd_sc_hd__a21oi_2 _4213_ (.A1(net88),
    .A2(_0484_),
    .B1(_2932_),
    .Y(_1301_));
 sky130_fd_sc_hd__and3_1 _4214_ (.A(net126),
    .B(_2868_),
    .C(net88),
    .X(_1302_));
 sky130_fd_sc_hd__a211oi_2 _4215_ (.A1(net140),
    .A2(_2992_),
    .B1(_2950_),
    .C1(_2887_),
    .Y(_1303_));
 sky130_fd_sc_hd__or2_1 _4216_ (.A(_1302_),
    .B(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__or2_1 _4217_ (.A(_1301_),
    .B(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__a311o_1 _4218_ (.A1(_2921_),
    .A2(_2964_),
    .A3(_0392_),
    .B1(_1300_),
    .C1(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__a22o_1 _4219_ (.A1(net154),
    .A2(\z80.tv80s.i_tv80_core.ISet[2] ),
    .B1(net160),
    .B2(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__or2_1 _4220_ (.A(_2942_),
    .B(_0762_),
    .X(_1308_));
 sky130_fd_sc_hd__or2_2 _4221_ (.A(_0383_),
    .B(_0545_),
    .X(_1309_));
 sky130_fd_sc_hd__and3b_2 _4222_ (.A_N(_2900_),
    .B(_2940_),
    .C(net113),
    .X(_1310_));
 sky130_fd_sc_hd__and3_1 _4223_ (.A(net125),
    .B(_2882_),
    .C(_1310_),
    .X(_1311_));
 sky130_fd_sc_hd__and3_1 _4224_ (.A(net147),
    .B(_0388_),
    .C(_0658_),
    .X(_1312_));
 sky130_fd_sc_hd__a21o_1 _4225_ (.A1(_2824_),
    .A2(_1312_),
    .B1(_1311_),
    .X(_1313_));
 sky130_fd_sc_hd__a211o_1 _4226_ (.A1(net142),
    .A2(_1313_),
    .B1(_1309_),
    .C1(_1308_),
    .X(_1314_));
 sky130_fd_sc_hd__o21ai_4 _4227_ (.A1(net99),
    .A2(_1307_),
    .B1(_1314_),
    .Y(_1315_));
 sky130_fd_sc_hd__nand2_1 _4228_ (.A(net142),
    .B(net125),
    .Y(_1316_));
 sky130_fd_sc_hd__a31o_1 _4229_ (.A1(_0417_),
    .A2(_0666_),
    .A3(_1316_),
    .B1(_1297_),
    .X(_1317_));
 sky130_fd_sc_hd__o21a_1 _4230_ (.A1(net124),
    .A2(_0540_),
    .B1(_0476_),
    .X(_1318_));
 sky130_fd_sc_hd__a31o_1 _4231_ (.A1(net147),
    .A2(_0501_),
    .A3(_0658_),
    .B1(_1318_),
    .X(_1319_));
 sky130_fd_sc_hd__a41o_1 _4232_ (.A1(net139),
    .A2(net125),
    .A3(_2880_),
    .A4(_2888_),
    .B1(_0692_),
    .X(_1320_));
 sky130_fd_sc_hd__a31o_1 _4233_ (.A1(_2911_),
    .A2(_2964_),
    .A3(_0392_),
    .B1(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__a211o_1 _4234_ (.A1(net139),
    .A2(_1317_),
    .B1(_1319_),
    .C1(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__a31o_1 _4235_ (.A1(\z80.tv80s.i_tv80_core.IR[5] ),
    .A2(_2880_),
    .A3(_1298_),
    .B1(net103),
    .X(_1323_));
 sky130_fd_sc_hd__o31a_1 _4236_ (.A1(_2940_),
    .A2(_1305_),
    .A3(_1322_),
    .B1(_1323_),
    .X(_1324_));
 sky130_fd_sc_hd__a21o_1 _4237_ (.A1(net151),
    .A2(\z80.tv80s.i_tv80_core.ISet[2] ),
    .B1(net100),
    .X(_1325_));
 sky130_fd_sc_hd__a21oi_1 _4238_ (.A1(net160),
    .A2(_1324_),
    .B1(_1325_),
    .Y(_1326_));
 sky130_fd_sc_hd__a41o_1 _4239_ (.A1(net139),
    .A2(net125),
    .A3(_2880_),
    .A4(_1310_),
    .B1(_1309_),
    .X(_1327_));
 sky130_fd_sc_hd__a21oi_1 _4240_ (.A1(_2911_),
    .A2(_1312_),
    .B1(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__a31o_2 _4241_ (.A1(_0683_),
    .A2(_0761_),
    .A3(_1328_),
    .B1(_1326_),
    .X(_1329_));
 sky130_fd_sc_hd__inv_2 _4242_ (.A(_1329_),
    .Y(_1330_));
 sky130_fd_sc_hd__nand2_1 _4243_ (.A(_0498_),
    .B(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__nand2b_1 _4244_ (.A_N(_1331_),
    .B(_1315_),
    .Y(_1332_));
 sky130_fd_sc_hd__mux2_1 _4245_ (.A0(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .A1(\z80.tv80s.i_tv80_core.Alternate ),
    .S(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(net218),
    .A1(_1333_),
    .S(net106),
    .X(_0049_));
 sky130_fd_sc_hd__or2_2 _4247_ (.A(net123),
    .B(net158),
    .X(_1334_));
 sky130_fd_sc_hd__nand2_1 _4248_ (.A(_2881_),
    .B(_2951_),
    .Y(_1335_));
 sky130_fd_sc_hd__a32o_1 _4249_ (.A1(_2881_),
    .A2(_2951_),
    .A3(_0513_),
    .B1(_0430_),
    .B2(_2888_),
    .X(_1336_));
 sky130_fd_sc_hd__a221o_1 _4250_ (.A1(net126),
    .A2(_2977_),
    .B1(_0662_),
    .B2(net130),
    .C1(_1336_),
    .X(_1337_));
 sky130_fd_sc_hd__a211o_1 _4251_ (.A1(net154),
    .A2(_1301_),
    .B1(_1302_),
    .C1(_2940_),
    .X(_1338_));
 sky130_fd_sc_hd__a31o_1 _4252_ (.A1(net142),
    .A2(_0395_),
    .A3(_0415_),
    .B1(_1338_),
    .X(_1339_));
 sky130_fd_sc_hd__a21o_1 _4253_ (.A1(net129),
    .A2(_2923_),
    .B1(_1297_),
    .X(_1340_));
 sky130_fd_sc_hd__a2111o_1 _4254_ (.A1(_2921_),
    .A2(_0692_),
    .B1(_1337_),
    .C1(_1339_),
    .D1(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__nand2_1 _4255_ (.A(net113),
    .B(_2881_),
    .Y(_1342_));
 sky130_fd_sc_hd__a31o_1 _4256_ (.A1(net154),
    .A2(_2885_),
    .A3(_1342_),
    .B1(net103),
    .X(_1343_));
 sky130_fd_sc_hd__nor3_2 _4257_ (.A(net113),
    .B(_2894_),
    .C(net102),
    .Y(_1344_));
 sky130_fd_sc_hd__a22o_1 _4258_ (.A1(_2944_),
    .A2(_0392_),
    .B1(_0442_),
    .B2(_0659_),
    .X(_1345_));
 sky130_fd_sc_hd__a21o_1 _4259_ (.A1(_2824_),
    .A2(_1345_),
    .B1(_1344_),
    .X(_1346_));
 sky130_fd_sc_hd__or2_1 _4260_ (.A(_0545_),
    .B(_1308_),
    .X(_1347_));
 sky130_fd_sc_hd__a221o_1 _4261_ (.A1(_3008_),
    .A2(_0395_),
    .B1(_1346_),
    .B2(net142),
    .C1(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__a32o_1 _4262_ (.A1(net160),
    .A2(_1341_),
    .A3(_1343_),
    .B1(_1348_),
    .B2(net100),
    .X(_1349_));
 sky130_fd_sc_hd__a22oi_4 _4263_ (.A1(net154),
    .A2(_1334_),
    .B1(_1349_),
    .B2(_2819_),
    .Y(_1350_));
 sky130_fd_sc_hd__inv_2 _4264_ (.A(_1350_),
    .Y(_1351_));
 sky130_fd_sc_hd__a31o_1 _4265_ (.A1(_2883_),
    .A2(_2940_),
    .A3(_1342_),
    .B1(_1301_),
    .X(_1352_));
 sky130_fd_sc_hd__a221o_1 _4266_ (.A1(_2911_),
    .A2(_0692_),
    .B1(_1352_),
    .B2(net151),
    .C1(_1318_),
    .X(_1353_));
 sky130_fd_sc_hd__a21oi_1 _4267_ (.A1(net114),
    .A2(_0501_),
    .B1(_2966_),
    .Y(_1354_));
 sky130_fd_sc_hd__nor2_1 _4268_ (.A(_0443_),
    .B(_1354_),
    .Y(_1355_));
 sky130_fd_sc_hd__a21o_1 _4269_ (.A1(_2823_),
    .A2(net125),
    .B1(net129),
    .X(_1356_));
 sky130_fd_sc_hd__nor2_1 _4270_ (.A(_2987_),
    .B(_0394_),
    .Y(_1357_));
 sky130_fd_sc_hd__a311o_1 _4271_ (.A1(net139),
    .A2(_0415_),
    .A3(_1356_),
    .B1(_1357_),
    .C1(_1302_),
    .X(_1358_));
 sky130_fd_sc_hd__a31o_1 _4272_ (.A1(_2974_),
    .A2(_0395_),
    .A3(_0473_),
    .B1(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__or4_1 _4273_ (.A(_1337_),
    .B(_1353_),
    .C(_1355_),
    .D(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__or2_1 _4274_ (.A(_0753_),
    .B(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__a22o_1 _4275_ (.A1(_3008_),
    .A2(_0483_),
    .B1(_1344_),
    .B2(net139),
    .X(_1362_));
 sky130_fd_sc_hd__a211o_1 _4276_ (.A1(_2911_),
    .A2(_1345_),
    .B1(_1347_),
    .C1(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__a22o_1 _4277_ (.A1(net160),
    .A2(_1361_),
    .B1(_1363_),
    .B2(net100),
    .X(_1364_));
 sky130_fd_sc_hd__a22o_4 _4278_ (.A1(net153),
    .A2(_1334_),
    .B1(_1364_),
    .B2(_2819_),
    .X(_1365_));
 sky130_fd_sc_hd__nand2_1 _4279_ (.A(_0498_),
    .B(_1365_),
    .Y(_1366_));
 sky130_fd_sc_hd__nor2_1 _4280_ (.A(_1351_),
    .B(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(\z80.tv80s.i_tv80_core.Alternate ),
    .A1(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .S(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__mux2_1 _4282_ (.A0(net538),
    .A1(_1368_),
    .S(net106),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _4283_ (.A(net101),
    .B(_0535_),
    .X(_1369_));
 sky130_fd_sc_hd__and3_4 _4284_ (.A(net150),
    .B(net101),
    .C(_0535_),
    .X(_1370_));
 sky130_fd_sc_hd__and3_2 _4285_ (.A(_2823_),
    .B(net116),
    .C(_1370_),
    .X(_1371_));
 sky130_fd_sc_hd__or3b_4 _4286_ (.A(net144),
    .B(_2831_),
    .C_N(_1370_),
    .X(_1372_));
 sky130_fd_sc_hd__xor2_1 _4287_ (.A(net723),
    .B(_0614_),
    .X(_1373_));
 sky130_fd_sc_hd__mux2_1 _4288_ (.A0(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A1(_1373_),
    .S(_1372_),
    .X(_1374_));
 sky130_fd_sc_hd__mux2_1 _4289_ (.A0(net723),
    .A1(_1374_),
    .S(net105),
    .X(_0051_));
 sky130_fd_sc_hd__a21oi_1 _4290_ (.A1(\z80.tv80s.i_tv80_core.R[0] ),
    .A2(_0614_),
    .B1(net578),
    .Y(_1375_));
 sky130_fd_sc_hd__a31o_1 _4291_ (.A1(\z80.tv80s.i_tv80_core.R[0] ),
    .A2(net578),
    .A3(_0614_),
    .B1(_1371_),
    .X(_1376_));
 sky130_fd_sc_hd__a2bb2o_1 _4292_ (.A1_N(_1375_),
    .A2_N(_1376_),
    .B1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .B2(_1371_),
    .X(_1377_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(net578),
    .A1(_1377_),
    .S(net105),
    .X(_0052_));
 sky130_fd_sc_hd__and2_1 _4294_ (.A(net105),
    .B(_1376_),
    .X(_1378_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A1(_2858_),
    .S(_1372_),
    .X(_1379_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(net624),
    .A1(_1379_),
    .S(_1378_),
    .X(_0053_));
 sky130_fd_sc_hd__a41o_1 _4297_ (.A1(\z80.tv80s.i_tv80_core.R[0] ),
    .A2(\z80.tv80s.i_tv80_core.R[1] ),
    .A3(\z80.tv80s.i_tv80_core.R[2] ),
    .A4(_0614_),
    .B1(net540),
    .X(_1380_));
 sky130_fd_sc_hd__and3_1 _4298_ (.A(\z80.tv80s.i_tv80_core.R[0] ),
    .B(net578),
    .C(\z80.tv80s.i_tv80_core.R[2] ),
    .X(_1381_));
 sky130_fd_sc_hd__and3_1 _4299_ (.A(net540),
    .B(_0598_),
    .C(_1381_),
    .X(_1382_));
 sky130_fd_sc_hd__nand2_1 _4300_ (.A(net95),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__a21o_1 _4301_ (.A1(_1372_),
    .A2(_1383_),
    .B1(net120),
    .X(_1384_));
 sky130_fd_sc_hd__a22o_1 _4302_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_1371_),
    .B1(_1380_),
    .B2(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__o21a_1 _4303_ (.A1(net105),
    .A2(net540),
    .B1(_1385_),
    .X(_0054_));
 sky130_fd_sc_hd__nor2_1 _4304_ (.A(net610),
    .B(_1383_),
    .Y(_1386_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A1(_1386_),
    .S(_1372_),
    .X(_1387_));
 sky130_fd_sc_hd__a22o_1 _4306_ (.A1(net610),
    .A2(_1384_),
    .B1(_1387_),
    .B2(net105),
    .X(_0055_));
 sky130_fd_sc_hd__and2_1 _4307_ (.A(\z80.tv80s.i_tv80_core.R[4] ),
    .B(_1382_),
    .X(_1388_));
 sky130_fd_sc_hd__a21oi_1 _4308_ (.A1(net131),
    .A2(_1388_),
    .B1(net586),
    .Y(_1389_));
 sky130_fd_sc_hd__and3_1 _4309_ (.A(net131),
    .B(net586),
    .C(_1388_),
    .X(_1390_));
 sky130_fd_sc_hd__or3_1 _4310_ (.A(_1371_),
    .B(_1389_),
    .C(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__o21ai_1 _4311_ (.A1(_2860_),
    .A2(_1372_),
    .B1(_1391_),
    .Y(_1392_));
 sky130_fd_sc_hd__mux2_1 _4312_ (.A0(net586),
    .A1(_1392_),
    .S(net108),
    .X(_0056_));
 sky130_fd_sc_hd__nand4_1 _4313_ (.A(net105),
    .B(net586),
    .C(net95),
    .D(_1388_),
    .Y(_1393_));
 sky130_fd_sc_hd__mux2_1 _4314_ (.A0(_1390_),
    .A1(_1393_),
    .S(net608),
    .X(_1394_));
 sky130_fd_sc_hd__or2_1 _4315_ (.A(_1371_),
    .B(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__nand2_1 _4316_ (.A(net105),
    .B(_1371_),
    .Y(_1396_));
 sky130_fd_sc_hd__o221a_1 _4317_ (.A1(net105),
    .A2(net608),
    .B1(_1396_),
    .B2(\z80.tv80s.i_tv80_core.ACC[6] ),
    .C1(_1395_),
    .X(_0057_));
 sky130_fd_sc_hd__nand2_2 _4318_ (.A(net161),
    .B(_2981_),
    .Y(_1397_));
 sky130_fd_sc_hd__and2_1 _4319_ (.A(net161),
    .B(_3019_),
    .X(_1398_));
 sky130_fd_sc_hd__nand2_1 _4320_ (.A(net161),
    .B(_3019_),
    .Y(_1399_));
 sky130_fd_sc_hd__nand2_1 _4321_ (.A(_1397_),
    .B(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__a21oi_1 _4322_ (.A1(net98),
    .A2(_1400_),
    .B1(net845),
    .Y(_1401_));
 sky130_fd_sc_hd__or2_1 _4323_ (.A(net845),
    .B(_1400_),
    .X(_1402_));
 sky130_fd_sc_hd__a22o_1 _4324_ (.A1(net553),
    .A2(_1401_),
    .B1(_1402_),
    .B2(net785),
    .X(_1403_));
 sky130_fd_sc_hd__mux2_1 _4325_ (.A0(net165),
    .A1(_1403_),
    .S(net106),
    .X(_0058_));
 sky130_fd_sc_hd__or2_1 _4326_ (.A(net106),
    .B(net164),
    .X(_1404_));
 sky130_fd_sc_hd__o31a_1 _4327_ (.A1(net119),
    .A2(_0492_),
    .A3(_1402_),
    .B1(_1404_),
    .X(_0059_));
 sky130_fd_sc_hd__nor2_4 _4328_ (.A(_0792_),
    .B(_0886_),
    .Y(_1405_));
 sky130_fd_sc_hd__mux2_1 _4329_ (.A0(net424),
    .A1(_0977_),
    .S(_1405_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4330_ (.A0(net416),
    .A1(_1018_),
    .S(_1405_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _4331_ (.A0(net433),
    .A1(_1059_),
    .S(_1405_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(net469),
    .A1(_1100_),
    .S(_1405_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _4333_ (.A0(net514),
    .A1(_1146_),
    .S(_1405_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(net362),
    .A1(_1193_),
    .S(_1405_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _4335_ (.A0(net364),
    .A1(_1238_),
    .S(_1405_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(net386),
    .A1(_1294_),
    .S(_1405_),
    .X(_0067_));
 sky130_fd_sc_hd__nor2_4 _4337_ (.A(_0792_),
    .B(_0878_),
    .Y(_1406_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(net314),
    .A1(_0977_),
    .S(_1406_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _4339_ (.A0(net268),
    .A1(_1018_),
    .S(_1406_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _4340_ (.A0(net280),
    .A1(_1059_),
    .S(_1406_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _4341_ (.A0(net324),
    .A1(_1100_),
    .S(_1406_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _4342_ (.A0(net294),
    .A1(_1146_),
    .S(_1406_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _4343_ (.A0(net360),
    .A1(_1193_),
    .S(_1406_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _4344_ (.A0(net296),
    .A1(_1238_),
    .S(_1406_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _4345_ (.A0(net390),
    .A1(_1294_),
    .S(_1406_),
    .X(_0075_));
 sky130_fd_sc_hd__nor2_2 _4346_ (.A(_3003_),
    .B(_0484_),
    .Y(_1407_));
 sky130_fd_sc_hd__or3_1 _4347_ (.A(net87),
    .B(_2975_),
    .C(_0511_),
    .X(_1408_));
 sky130_fd_sc_hd__nor2_1 _4348_ (.A(_0711_),
    .B(_1408_),
    .Y(_1409_));
 sky130_fd_sc_hd__or4b_1 _4349_ (.A(net111),
    .B(_0710_),
    .C(_1296_),
    .D_N(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__o2bb2ai_1 _4350_ (.A1_N(net101),
    .A2_N(_1407_),
    .B1(_1410_),
    .B2(_0707_),
    .Y(_1411_));
 sky130_fd_sc_hd__mux2_1 _4351_ (.A0(net521),
    .A1(_1411_),
    .S(net109),
    .X(_0076_));
 sky130_fd_sc_hd__nor2_4 _4352_ (.A(_0792_),
    .B(_0876_),
    .Y(_1412_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(net355),
    .A1(_0977_),
    .S(_1412_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(net343),
    .A1(_1018_),
    .S(_1412_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _4355_ (.A0(net326),
    .A1(_1059_),
    .S(_1412_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _4356_ (.A0(net380),
    .A1(_1100_),
    .S(_1412_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _4357_ (.A0(net337),
    .A1(_1146_),
    .S(_1412_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _4358_ (.A0(net463),
    .A1(_1193_),
    .S(_1412_),
    .X(_0082_));
 sky130_fd_sc_hd__mux2_1 _4359_ (.A0(net316),
    .A1(_1238_),
    .S(_1412_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _4360_ (.A0(net351),
    .A1(_1294_),
    .S(_1412_),
    .X(_0084_));
 sky130_fd_sc_hd__or3b_1 _4361_ (.A(_2854_),
    .B(_0790_),
    .C_N(_0788_),
    .X(_1413_));
 sky130_fd_sc_hd__a41o_4 _4362_ (.A1(_0778_),
    .A2(net84),
    .A3(net83),
    .A4(_1413_),
    .B1(net119),
    .X(_1414_));
 sky130_fd_sc_hd__nor2_4 _4363_ (.A(_0886_),
    .B(_1414_),
    .Y(_1415_));
 sky130_fd_sc_hd__mux4_1 _4364_ (.A0(net270),
    .A1(net312),
    .A2(net308),
    .A3(net322),
    .S0(net77),
    .S1(net73),
    .X(_1416_));
 sky130_fd_sc_hd__a21o_1 _4365_ (.A1(net69),
    .A2(_0960_),
    .B1(_0864_),
    .X(_1417_));
 sky130_fd_sc_hd__a21oi_1 _4366_ (.A1(_2864_),
    .A2(_0782_),
    .B1(net86),
    .Y(_1418_));
 sky130_fd_sc_hd__a22o_2 _4367_ (.A1(net86),
    .A2(_1416_),
    .B1(_1417_),
    .B2(_1418_),
    .X(_1419_));
 sky130_fd_sc_hd__mux2_1 _4368_ (.A0(net404),
    .A1(_1419_),
    .S(_1415_),
    .X(_0085_));
 sky130_fd_sc_hd__or3_1 _4369_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .B(net135),
    .C(net86),
    .X(_1420_));
 sky130_fd_sc_hd__o211a_1 _4370_ (.A1(net471),
    .A2(net77),
    .B1(net73),
    .C1(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__mux2_1 _4371_ (.A0(net284),
    .A1(net384),
    .S(net77),
    .X(_1422_));
 sky130_fd_sc_hd__o221a_1 _4372_ (.A1(net292),
    .A2(net135),
    .B1(net77),
    .B2(net274),
    .C1(net73),
    .X(_1423_));
 sky130_fd_sc_hd__o221a_1 _4373_ (.A1(net456),
    .A2(net135),
    .B1(net77),
    .B2(net332),
    .C1(net71),
    .X(_1424_));
 sky130_fd_sc_hd__a221o_1 _4374_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .A2(_0781_),
    .B1(net71),
    .B2(_1422_),
    .C1(_1421_),
    .X(_1425_));
 sky130_fd_sc_hd__o31a_1 _4375_ (.A1(_1286_),
    .A2(_1423_),
    .A3(_1424_),
    .B1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__nand2_1 _4376_ (.A(_0951_),
    .B(_0960_),
    .Y(_1427_));
 sky130_fd_sc_hd__o21a_1 _4377_ (.A1(_0951_),
    .A2(_0960_),
    .B1(_0819_),
    .X(_1428_));
 sky130_fd_sc_hd__a21o_1 _4378_ (.A1(_1427_),
    .A2(_1428_),
    .B1(_1005_),
    .X(_1429_));
 sky130_fd_sc_hd__a21oi_1 _4379_ (.A1(_2865_),
    .A2(_0782_),
    .B1(net86),
    .Y(_1430_));
 sky130_fd_sc_hd__a22o_2 _4380_ (.A1(net86),
    .A2(_1426_),
    .B1(_1429_),
    .B2(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__mux2_1 _4381_ (.A0(net292),
    .A1(_1431_),
    .S(_1415_),
    .X(_0086_));
 sky130_fd_sc_hd__or3_1 _4382_ (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .B(net135),
    .C(net86),
    .X(_1432_));
 sky130_fd_sc_hd__o211a_1 _4383_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .A2(net77),
    .B1(net73),
    .C1(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__mux2_1 _4384_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .S(net77),
    .X(_1434_));
 sky130_fd_sc_hd__o221a_1 _4385_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A2(net135),
    .B1(_0814_),
    .B2(net290),
    .C1(net73),
    .X(_1435_));
 sky130_fd_sc_hd__o221a_1 _4386_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A2(net135),
    .B1(net77),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .C1(net71),
    .X(_1436_));
 sky130_fd_sc_hd__a221o_1 _4387_ (.A1(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .A2(_0781_),
    .B1(net71),
    .B2(_1434_),
    .C1(_1433_),
    .X(_1437_));
 sky130_fd_sc_hd__o31a_1 _4388_ (.A1(_1286_),
    .A2(_1435_),
    .A3(_1436_),
    .B1(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__xor2_1 _4389_ (.A(_0961_),
    .B(_0962_),
    .X(_1439_));
 sky130_fd_sc_hd__a21o_1 _4390_ (.A1(_0819_),
    .A2(_1439_),
    .B1(_1055_),
    .X(_1440_));
 sky130_fd_sc_hd__o21a_1 _4391_ (.A1(net240),
    .A2(net83),
    .B1(net84),
    .X(_1441_));
 sky130_fd_sc_hd__a22o_2 _4392_ (.A1(net85),
    .A2(_1438_),
    .B1(_1440_),
    .B2(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__mux2_1 _4393_ (.A0(net262),
    .A1(_1442_),
    .S(_1415_),
    .X(_0087_));
 sky130_fd_sc_hd__xnor2_1 _4394_ (.A(_0873_),
    .B(_0927_),
    .Y(_1443_));
 sky130_fd_sc_hd__xnor2_1 _4395_ (.A(_0964_),
    .B(_1443_),
    .Y(_1444_));
 sky130_fd_sc_hd__nor2_1 _4396_ (.A(_0820_),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__o221a_1 _4397_ (.A1(net232),
    .A2(net82),
    .B1(_1088_),
    .B2(_1445_),
    .C1(net84),
    .X(_1446_));
 sky130_fd_sc_hd__mux4_2 _4398_ (.A0(net398),
    .A1(net276),
    .A2(net502),
    .A3(net258),
    .S0(net73),
    .S1(net77),
    .X(_1447_));
 sky130_fd_sc_hd__a21o_2 _4399_ (.A1(net85),
    .A2(_1447_),
    .B1(_1446_),
    .X(_1448_));
 sky130_fd_sc_hd__mux2_1 _4400_ (.A0(net478),
    .A1(_1448_),
    .S(_1415_),
    .X(_0088_));
 sky130_fd_sc_hd__xnor2_1 _4401_ (.A(_0922_),
    .B(_0966_),
    .Y(_1449_));
 sky130_fd_sc_hd__a21bo_1 _4402_ (.A1(net69),
    .A2(_1449_),
    .B1_N(_1142_),
    .X(_1450_));
 sky130_fd_sc_hd__o21a_1 _4403_ (.A1(net228),
    .A2(net82),
    .B1(net84),
    .X(_1451_));
 sky130_fd_sc_hd__mux4_2 _4404_ (.A0(net474),
    .A1(net278),
    .A2(net483),
    .A3(net310),
    .S0(net72),
    .S1(net75),
    .X(_1452_));
 sky130_fd_sc_hd__a22o_2 _4405_ (.A1(_1450_),
    .A2(_1451_),
    .B1(_1452_),
    .B2(net85),
    .X(_1453_));
 sky130_fd_sc_hd__mux2_1 _4406_ (.A0(net439),
    .A1(_1453_),
    .S(_1415_),
    .X(_0089_));
 sky130_fd_sc_hd__and2b_1 _4407_ (.A_N(_0921_),
    .B(_0967_),
    .X(_1454_));
 sky130_fd_sc_hd__xnor2_1 _4408_ (.A(_0915_),
    .B(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__nor2_1 _4409_ (.A(_0820_),
    .B(_1455_),
    .Y(_1456_));
 sky130_fd_sc_hd__o221a_1 _4410_ (.A1(net222),
    .A2(net82),
    .B1(_1179_),
    .B2(_1456_),
    .C1(net84),
    .X(_1457_));
 sky130_fd_sc_hd__mux4_2 _4411_ (.A0(net304),
    .A1(net266),
    .A2(net445),
    .A3(net358),
    .S0(net72),
    .S1(net75),
    .X(_1458_));
 sky130_fd_sc_hd__a21o_2 _4412_ (.A1(net85),
    .A2(_1458_),
    .B1(_1457_),
    .X(_1459_));
 sky130_fd_sc_hd__mux2_1 _4413_ (.A0(net468),
    .A1(_1459_),
    .S(_1415_),
    .X(_0090_));
 sky130_fd_sc_hd__a211o_1 _4414_ (.A1(net68),
    .A2(_0914_),
    .B1(_0921_),
    .C1(_0968_),
    .X(_1460_));
 sky130_fd_sc_hd__and2b_1 _4415_ (.A_N(_0908_),
    .B(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__xnor2_1 _4416_ (.A(_0908_),
    .B(_1460_),
    .Y(_1462_));
 sky130_fd_sc_hd__a21bo_1 _4417_ (.A1(net69),
    .A2(_1462_),
    .B1_N(_1234_),
    .X(_1463_));
 sky130_fd_sc_hd__o21a_1 _4418_ (.A1(net220),
    .A2(net82),
    .B1(net84),
    .X(_1464_));
 sky130_fd_sc_hd__mux4_1 _4419_ (.A0(net298),
    .A1(net353),
    .A2(net306),
    .A3(net376),
    .S0(net73),
    .S1(_0814_),
    .X(_1465_));
 sky130_fd_sc_hd__a22o_2 _4420_ (.A1(_1463_),
    .A2(_1464_),
    .B1(_1465_),
    .B2(net85),
    .X(_1466_));
 sky130_fd_sc_hd__mux2_1 _4421_ (.A0(net349),
    .A1(_1466_),
    .S(_1415_),
    .X(_0091_));
 sky130_fd_sc_hd__a21oi_1 _4422_ (.A1(_0874_),
    .A2(_0907_),
    .B1(_1461_),
    .Y(_1467_));
 sky130_fd_sc_hd__xnor2_1 _4423_ (.A(_0901_),
    .B(_1467_),
    .Y(_1468_));
 sky130_fd_sc_hd__nor2_1 _4424_ (.A(_0820_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__o22a_1 _4425_ (.A1(net224),
    .A2(net82),
    .B1(_1283_),
    .B2(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__mux4_1 _4426_ (.A0(net458),
    .A1(net282),
    .A2(net500),
    .A3(net288),
    .S0(net73),
    .S1(net77),
    .X(_1471_));
 sky130_fd_sc_hd__mux2_2 _4427_ (.A0(_1470_),
    .A1(_1471_),
    .S(net85),
    .X(_1472_));
 sky130_fd_sc_hd__mux2_1 _4428_ (.A0(net476),
    .A1(_1472_),
    .S(_1415_),
    .X(_0092_));
 sky130_fd_sc_hd__nor2_4 _4429_ (.A(_0792_),
    .B(_0891_),
    .Y(_1473_));
 sky130_fd_sc_hd__mux2_1 _4430_ (.A0(net495),
    .A1(_0977_),
    .S(_1473_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4431_ (.A0(net402),
    .A1(_1018_),
    .S(_1473_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4432_ (.A0(net437),
    .A1(_1059_),
    .S(_1473_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4433_ (.A0(net446),
    .A1(_1100_),
    .S(_1473_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4434_ (.A0(net443),
    .A1(_1146_),
    .S(_1473_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _4435_ (.A0(net499),
    .A1(_1193_),
    .S(_1473_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _4436_ (.A0(net415),
    .A1(_1238_),
    .S(_1473_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _4437_ (.A0(net382),
    .A1(_1294_),
    .S(_1473_),
    .X(_0100_));
 sky130_fd_sc_hd__nor2_4 _4438_ (.A(_0878_),
    .B(_1414_),
    .Y(_1474_));
 sky130_fd_sc_hd__mux2_1 _4439_ (.A0(net308),
    .A1(_1419_),
    .S(_1474_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _4440_ (.A0(net471),
    .A1(_1431_),
    .S(_1474_),
    .X(_0102_));
 sky130_fd_sc_hd__mux2_1 _4441_ (.A0(net272),
    .A1(_1442_),
    .S(_1474_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _4442_ (.A0(net276),
    .A1(_1448_),
    .S(_1474_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _4443_ (.A0(net278),
    .A1(_1453_),
    .S(_1474_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _4444_ (.A0(net266),
    .A1(_1459_),
    .S(_1474_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4445_ (.A0(net353),
    .A1(_1466_),
    .S(_1474_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _4446_ (.A0(net282),
    .A1(_1472_),
    .S(_1474_),
    .X(_0108_));
 sky130_fd_sc_hd__or2_4 _4447_ (.A(_0792_),
    .B(_0883_),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_1 _4448_ (.A0(_0977_),
    .A1(net450),
    .S(_1475_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4449_ (.A0(_1018_),
    .A1(net420),
    .S(_1475_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4450_ (.A0(_1059_),
    .A1(net400),
    .S(_1475_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4451_ (.A0(_1100_),
    .A1(net488),
    .S(_1475_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4452_ (.A0(_1146_),
    .A1(net452),
    .S(_1475_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4453_ (.A0(_1193_),
    .A1(net302),
    .S(_1475_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_1 _4454_ (.A0(_1238_),
    .A1(net357),
    .S(_1475_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _4455_ (.A0(_1294_),
    .A1(net366),
    .S(_1475_),
    .X(_0116_));
 sky130_fd_sc_hd__or2_4 _4456_ (.A(_0881_),
    .B(_1414_),
    .X(_1476_));
 sky130_fd_sc_hd__mux2_1 _4457_ (.A0(_1419_),
    .A1(net312),
    .S(_1476_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _4458_ (.A0(_1431_),
    .A1(net384),
    .S(_1476_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _4459_ (.A0(_1442_),
    .A1(net328),
    .S(_1476_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _4460_ (.A0(_1448_),
    .A1(net502),
    .S(_1476_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _4461_ (.A0(_1453_),
    .A1(net483),
    .S(_1476_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4462_ (.A0(_1459_),
    .A1(net445),
    .S(_1476_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4463_ (.A0(_1466_),
    .A1(net306),
    .S(_1476_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4464_ (.A0(_1472_),
    .A1(net500),
    .S(_1476_),
    .X(_0124_));
 sky130_fd_sc_hd__or2_4 _4465_ (.A(_0883_),
    .B(_1414_),
    .X(_1477_));
 sky130_fd_sc_hd__mux2_1 _4466_ (.A0(_1419_),
    .A1(net270),
    .S(_1477_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4467_ (.A0(_1431_),
    .A1(net284),
    .S(_1477_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4468_ (.A0(_1442_),
    .A1(net260),
    .S(_1477_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _4469_ (.A0(_1448_),
    .A1(net398),
    .S(_1477_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4470_ (.A0(_1453_),
    .A1(net474),
    .S(_1477_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _4471_ (.A0(_1459_),
    .A1(net304),
    .S(_1477_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4472_ (.A0(_1466_),
    .A1(net298),
    .S(_1477_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4473_ (.A0(_1472_),
    .A1(net458),
    .S(_1477_),
    .X(_0132_));
 sky130_fd_sc_hd__or2_4 _4474_ (.A(_0812_),
    .B(_1414_),
    .X(_1478_));
 sky130_fd_sc_hd__mux2_1 _4475_ (.A0(_1419_),
    .A1(net431),
    .S(_1478_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4476_ (.A0(_1431_),
    .A1(net332),
    .S(_1478_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4477_ (.A0(_1442_),
    .A1(net372),
    .S(_1478_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4478_ (.A0(_1448_),
    .A1(net489),
    .S(_1478_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4479_ (.A0(_1453_),
    .A1(net435),
    .S(_1478_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4480_ (.A0(_1459_),
    .A1(net427),
    .S(_1478_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4481_ (.A0(_1466_),
    .A1(net410),
    .S(_1478_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4482_ (.A0(_1472_),
    .A1(net493),
    .S(_1478_),
    .X(_0140_));
 sky130_fd_sc_hd__nor2_4 _4483_ (.A(_0876_),
    .B(_1414_),
    .Y(_1479_));
 sky130_fd_sc_hd__mux2_1 _4484_ (.A0(net322),
    .A1(_1419_),
    .S(_1479_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4485_ (.A0(net491),
    .A1(_1431_),
    .S(_1479_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_1 _4486_ (.A0(net256),
    .A1(_1442_),
    .S(_1479_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4487_ (.A0(net258),
    .A1(_1448_),
    .S(_1479_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4488_ (.A0(net310),
    .A1(_1453_),
    .S(_1479_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4489_ (.A0(net358),
    .A1(_1459_),
    .S(_1479_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4490_ (.A0(net376),
    .A1(_1466_),
    .S(_1479_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _4491_ (.A0(net288),
    .A1(_1472_),
    .S(_1479_),
    .X(_0148_));
 sky130_fd_sc_hd__or2_4 _4492_ (.A(_0792_),
    .B(_0888_),
    .X(_1480_));
 sky130_fd_sc_hd__mux2_1 _4493_ (.A0(_0977_),
    .A1(net509),
    .S(_1480_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4494_ (.A0(_1018_),
    .A1(net455),
    .S(_1480_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4495_ (.A0(_1059_),
    .A1(net461),
    .S(_1480_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4496_ (.A0(_1100_),
    .A1(net498),
    .S(_1480_),
    .X(_0152_));
 sky130_fd_sc_hd__mux2_1 _4497_ (.A0(_1146_),
    .A1(net501),
    .S(_1480_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4498_ (.A0(_1193_),
    .A1(net480),
    .S(_1480_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4499_ (.A0(_1238_),
    .A1(net460),
    .S(_1480_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4500_ (.A0(_1294_),
    .A1(net503),
    .S(_1480_),
    .X(_0156_));
 sky130_fd_sc_hd__nor2_4 _4501_ (.A(_0891_),
    .B(_1414_),
    .Y(_1481_));
 sky130_fd_sc_hd__mux2_1 _4502_ (.A0(net341),
    .A1(_1419_),
    .S(_1481_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _4503_ (.A0(net274),
    .A1(_1431_),
    .S(_1481_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4504_ (.A0(net290),
    .A1(_1442_),
    .S(_1481_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4505_ (.A0(net378),
    .A1(_1448_),
    .S(_1481_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4506_ (.A0(net394),
    .A1(_1453_),
    .S(_1481_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _4507_ (.A0(net406),
    .A1(_1459_),
    .S(_1481_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _4508_ (.A0(net370),
    .A1(_1466_),
    .S(_1481_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4509_ (.A0(net368),
    .A1(_1472_),
    .S(_1481_),
    .X(_0164_));
 sky130_fd_sc_hd__or2_4 _4510_ (.A(_0792_),
    .B(_0881_),
    .X(_1482_));
 sky130_fd_sc_hd__mux2_1 _4511_ (.A0(_0977_),
    .A1(net396),
    .S(_1482_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_1 _4512_ (.A0(_1018_),
    .A1(net426),
    .S(_1482_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_1 _4513_ (.A0(_1059_),
    .A1(net505),
    .S(_1482_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_1 _4514_ (.A0(_1100_),
    .A1(net448),
    .S(_1482_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_1 _4515_ (.A0(_1146_),
    .A1(net429),
    .S(_1482_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _4516_ (.A0(_1193_),
    .A1(net320),
    .S(_1482_),
    .X(_0170_));
 sky130_fd_sc_hd__mux2_1 _4517_ (.A0(_1238_),
    .A1(net300),
    .S(_1482_),
    .X(_0171_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(_1294_),
    .A1(net339),
    .S(_1482_),
    .X(_0172_));
 sky130_fd_sc_hd__and2_4 _4519_ (.A(net161),
    .B(_2960_),
    .X(_1483_));
 sky130_fd_sc_hd__nand2_2 _4520_ (.A(net162),
    .B(_2960_),
    .Y(_1484_));
 sky130_fd_sc_hd__and3_4 _4521_ (.A(net108),
    .B(net92),
    .C(_1483_),
    .X(_1485_));
 sky130_fd_sc_hd__or4_2 _4522_ (.A(net111),
    .B(_2871_),
    .C(_2887_),
    .D(_2901_),
    .X(_1486_));
 sky130_fd_sc_hd__or2_2 _4523_ (.A(net97),
    .B(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__mux2_1 _4524_ (.A0(net703),
    .A1(\z80.tv80s.i_tv80_core.ACC[0] ),
    .S(_1485_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_1 _4525_ (.A0(net670),
    .A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .S(_1485_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_1 _4526_ (.A0(net668),
    .A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .S(_1485_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_1 _4527_ (.A0(net705),
    .A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .S(_1485_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_1 _4528_ (.A0(net693),
    .A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .S(_1485_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_1 _4529_ (.A0(net683),
    .A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .S(_1485_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_1 _4530_ (.A0(net660),
    .A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .S(_1485_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_1 _4531_ (.A0(net662),
    .A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .S(_1485_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_1 _4532_ (.A0(net707),
    .A1(net138),
    .S(_1485_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_1 _4533_ (.A0(net745),
    .A1(\z80.tv80s.i_tv80_core.F[1] ),
    .S(_1485_),
    .X(_0182_));
 sky130_fd_sc_hd__mux2_1 _4534_ (.A0(net681),
    .A1(\z80.tv80s.i_tv80_core.F[2] ),
    .S(_1485_),
    .X(_0183_));
 sky130_fd_sc_hd__mux2_1 _4535_ (.A0(net697),
    .A1(\z80.tv80s.i_tv80_core.F[3] ),
    .S(_1485_),
    .X(_0184_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(net699),
    .A1(\z80.tv80s.i_tv80_core.F[4] ),
    .S(_1485_),
    .X(_0185_));
 sky130_fd_sc_hd__mux2_1 _4537_ (.A0(net695),
    .A1(\z80.tv80s.i_tv80_core.F[5] ),
    .S(_1485_),
    .X(_0186_));
 sky130_fd_sc_hd__mux2_1 _4538_ (.A0(net676),
    .A1(\z80.tv80s.i_tv80_core.F[6] ),
    .S(_1485_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _4539_ (.A0(net685),
    .A1(\z80.tv80s.i_tv80_core.F[7] ),
    .S(_1485_),
    .X(_0188_));
 sky130_fd_sc_hd__a21o_1 _4540_ (.A1(_2948_),
    .A2(_1312_),
    .B1(_2942_),
    .X(_1488_));
 sky130_fd_sc_hd__and4_1 _4541_ (.A(net125),
    .B(net113),
    .C(_2948_),
    .D(_0417_),
    .X(_1489_));
 sky130_fd_sc_hd__a31o_1 _4542_ (.A1(_2948_),
    .A2(_2964_),
    .A3(_0392_),
    .B1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__a22oi_4 _4543_ (.A1(net99),
    .A2(_1488_),
    .B1(_1490_),
    .B2(net160),
    .Y(_1491_));
 sky130_fd_sc_hd__inv_2 _4544_ (.A(_1491_),
    .Y(_1492_));
 sky130_fd_sc_hd__nand2_2 _4545_ (.A(_1315_),
    .B(_1329_),
    .Y(_1493_));
 sky130_fd_sc_hd__a21oi_4 _4546_ (.A1(_1492_),
    .A2(_1493_),
    .B1(net119),
    .Y(_1494_));
 sky130_fd_sc_hd__a21oi_1 _4547_ (.A1(_2920_),
    .A2(_0651_),
    .B1(_2887_),
    .Y(_1495_));
 sky130_fd_sc_hd__o21a_1 _4548_ (.A1(_0476_),
    .A2(_1495_),
    .B1(net125),
    .X(_1496_));
 sky130_fd_sc_hd__o21a_1 _4549_ (.A1(_2829_),
    .A2(_2949_),
    .B1(_2825_),
    .X(_1497_));
 sky130_fd_sc_hd__nor3_1 _4550_ (.A(net129),
    .B(_0418_),
    .C(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__a21oi_2 _4551_ (.A1(net125),
    .A2(_2948_),
    .B1(_1497_),
    .Y(_1499_));
 sky130_fd_sc_hd__a221o_1 _4552_ (.A1(net146),
    .A2(_0425_),
    .B1(_1499_),
    .B2(_2964_),
    .C1(_2940_),
    .X(_1500_));
 sky130_fd_sc_hd__a311o_1 _4553_ (.A1(net146),
    .A2(_0501_),
    .A3(_0541_),
    .B1(_1498_),
    .C1(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__a21o_1 _4554_ (.A1(net146),
    .A2(_1298_),
    .B1(net103),
    .X(_1502_));
 sky130_fd_sc_hd__o31a_1 _4555_ (.A1(_1305_),
    .A2(_1496_),
    .A3(_1501_),
    .B1(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__a211o_1 _4556_ (.A1(net147),
    .A2(_1310_),
    .B1(_0440_),
    .C1(_2944_),
    .X(_1504_));
 sky130_fd_sc_hd__or2_1 _4557_ (.A(_2830_),
    .B(_2949_),
    .X(_1505_));
 sky130_fd_sc_hd__nand2_1 _4558_ (.A(_2830_),
    .B(_2949_),
    .Y(_1506_));
 sky130_fd_sc_hd__a32o_1 _4559_ (.A1(_1312_),
    .A2(_1505_),
    .A3(_1506_),
    .B1(_1504_),
    .B2(net124),
    .X(_1507_));
 sky130_fd_sc_hd__o21a_1 _4560_ (.A1(_0545_),
    .A2(_1507_),
    .B1(net99),
    .X(_1508_));
 sky130_fd_sc_hd__a221o_4 _4561_ (.A1(net156),
    .A2(net158),
    .B1(net159),
    .B2(_1503_),
    .C1(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__nor2_2 _4562_ (.A(_1315_),
    .B(_1329_),
    .Y(_1510_));
 sky130_fd_sc_hd__nor2_4 _4563_ (.A(_1492_),
    .B(_1510_),
    .Y(_1511_));
 sky130_fd_sc_hd__inv_2 _4564_ (.A(_1511_),
    .Y(_1512_));
 sky130_fd_sc_hd__mux2_1 _4565_ (.A0(_0893_),
    .A1(_0960_),
    .S(_1509_),
    .X(_1513_));
 sky130_fd_sc_hd__nor2_1 _4566_ (.A(_1512_),
    .B(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__nor3_4 _4567_ (.A(_1491_),
    .B(_1493_),
    .C(_1509_),
    .Y(_1515_));
 sky130_fd_sc_hd__and4_2 _4568_ (.A(_1315_),
    .B(_1329_),
    .C(_1492_),
    .D(_1509_),
    .X(_1516_));
 sky130_fd_sc_hd__and2b_2 _4569_ (.A_N(_1509_),
    .B(_1510_),
    .X(_1517_));
 sky130_fd_sc_hd__and2_2 _4570_ (.A(_1509_),
    .B(_1510_),
    .X(_1518_));
 sky130_fd_sc_hd__a221o_1 _4571_ (.A1(\z80.tv80s.di_reg[0] ),
    .A2(_1517_),
    .B1(_1518_),
    .B2(\z80.tv80s.i_tv80_core.ACC[0] ),
    .C1(_1514_),
    .X(_1519_));
 sky130_fd_sc_hd__a221o_1 _4572_ (.A1(\z80.tv80s.i_tv80_core.SP[0] ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\z80.tv80s.i_tv80_core.SP[8] ),
    .C1(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__a22o_1 _4573_ (.A1(net120),
    .A2(net646),
    .B1(_1494_),
    .B2(_1520_),
    .X(_0189_));
 sky130_fd_sc_hd__nand2_1 _4574_ (.A(_0947_),
    .B(_1509_),
    .Y(_1521_));
 sky130_fd_sc_hd__o211a_1 _4575_ (.A1(_1011_),
    .A2(_1509_),
    .B1(_1511_),
    .C1(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__a221o_1 _4576_ (.A1(\z80.tv80s.di_reg[1] ),
    .A2(_1517_),
    .B1(_1518_),
    .B2(\z80.tv80s.i_tv80_core.ACC[1] ),
    .C1(_1522_),
    .X(_1523_));
 sky130_fd_sc_hd__a221o_1 _4577_ (.A1(net654),
    .A2(_1515_),
    .B1(_1516_),
    .B2(net604),
    .C1(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__a22o_1 _4578_ (.A1(net120),
    .A2(net766),
    .B1(_1494_),
    .B2(_1524_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4579_ (.A0(_1023_),
    .A1(_0937_),
    .S(_1509_),
    .X(_1525_));
 sky130_fd_sc_hd__a22o_1 _4580_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_1517_),
    .B1(_1518_),
    .B2(\z80.tv80s.i_tv80_core.ACC[2] ),
    .X(_1526_));
 sky130_fd_sc_hd__a221o_1 _4581_ (.A1(net652),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\z80.tv80s.i_tv80_core.SP[10] ),
    .C1(_1526_),
    .X(_1527_));
 sky130_fd_sc_hd__a21o_1 _4582_ (.A1(_1511_),
    .A2(_1525_),
    .B1(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__a22o_1 _4583_ (.A1(net120),
    .A2(net658),
    .B1(_1494_),
    .B2(_1528_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _4584_ (.A0(_1093_),
    .A1(_0927_),
    .S(_1509_),
    .X(_1529_));
 sky130_fd_sc_hd__a22o_1 _4585_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_1517_),
    .B1(_1518_),
    .B2(\z80.tv80s.i_tv80_core.ACC[3] ),
    .X(_1530_));
 sky130_fd_sc_hd__a221o_1 _4586_ (.A1(net672),
    .A2(_1515_),
    .B1(_1516_),
    .B2(net628),
    .C1(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__a21o_1 _4587_ (.A1(_1511_),
    .A2(_1529_),
    .B1(_1531_),
    .X(_1532_));
 sky130_fd_sc_hd__a22o_1 _4588_ (.A1(net120),
    .A2(net687),
    .B1(_1494_),
    .B2(_1532_),
    .X(_0192_));
 sky130_fd_sc_hd__mux2_1 _4589_ (.A0(_1110_),
    .A1(_0920_),
    .S(_1509_),
    .X(_1533_));
 sky130_fd_sc_hd__a22o_1 _4590_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_1517_),
    .B1(_1518_),
    .B2(\z80.tv80s.i_tv80_core.ACC[4] ),
    .X(_1534_));
 sky130_fd_sc_hd__a221o_1 _4591_ (.A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(net616),
    .C1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__a21o_1 _4592_ (.A1(_1511_),
    .A2(_1533_),
    .B1(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__a22o_1 _4593_ (.A1(net120),
    .A2(net637),
    .B1(_1494_),
    .B2(_1536_),
    .X(_0193_));
 sky130_fd_sc_hd__nand2_1 _4594_ (.A(_0913_),
    .B(_1509_),
    .Y(_1537_));
 sky130_fd_sc_hd__o211a_1 _4595_ (.A1(_1185_),
    .A2(_1509_),
    .B1(_1511_),
    .C1(_1537_),
    .X(_1538_));
 sky130_fd_sc_hd__a221o_1 _4596_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_1517_),
    .B1(_1518_),
    .B2(\z80.tv80s.i_tv80_core.ACC[5] ),
    .C1(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__a221o_1 _4597_ (.A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\z80.tv80s.i_tv80_core.SP[13] ),
    .C1(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__a22o_1 _4598_ (.A1(net120),
    .A2(net717),
    .B1(_1494_),
    .B2(_1540_),
    .X(_0194_));
 sky130_fd_sc_hd__nand2_1 _4599_ (.A(_0906_),
    .B(_1509_),
    .Y(_1541_));
 sky130_fd_sc_hd__o211a_1 _4600_ (.A1(_1199_),
    .A2(_1509_),
    .B1(_1511_),
    .C1(_1541_),
    .X(_1542_));
 sky130_fd_sc_hd__a221o_1 _4601_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_1517_),
    .B1(_1518_),
    .B2(\z80.tv80s.i_tv80_core.ACC[6] ),
    .C1(_1542_),
    .X(_1543_));
 sky130_fd_sc_hd__a221o_1 _4602_ (.A1(net631),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\z80.tv80s.i_tv80_core.SP[14] ),
    .C1(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__a22o_1 _4603_ (.A1(net120),
    .A2(net749),
    .B1(_1494_),
    .B2(_1544_),
    .X(_0195_));
 sky130_fd_sc_hd__mux2_1 _4604_ (.A0(_1244_),
    .A1(_0900_),
    .S(_1509_),
    .X(_1545_));
 sky130_fd_sc_hd__a22o_1 _4605_ (.A1(\z80.tv80s.di_reg[7] ),
    .A2(_1517_),
    .B1(_1518_),
    .B2(\z80.tv80s.i_tv80_core.ACC[7] ),
    .X(_1546_));
 sky130_fd_sc_hd__a221o_1 _4606_ (.A1(\z80.tv80s.i_tv80_core.SP[7] ),
    .A2(_1515_),
    .B1(_1516_),
    .B2(\z80.tv80s.i_tv80_core.SP[15] ),
    .C1(_1546_),
    .X(_1547_));
 sky130_fd_sc_hd__a21o_1 _4607_ (.A1(_1511_),
    .A2(_1545_),
    .B1(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__a22o_1 _4608_ (.A1(\z80.tv80s.i_tv80_core.BusAck ),
    .A2(net533),
    .B1(_1494_),
    .B2(_1548_),
    .X(_0196_));
 sky130_fd_sc_hd__and2b_1 _4609_ (.A_N(net10),
    .B(net584),
    .X(_1549_));
 sky130_fd_sc_hd__o21ba_1 _4610_ (.A1(net484),
    .A2(_1549_),
    .B1_N(\z80.tv80s.i_tv80_core.NMICycle ),
    .X(_0197_));
 sky130_fd_sc_hd__a211o_1 _4611_ (.A1(net648),
    .A2(net576),
    .B1(net773),
    .C1(net890),
    .X(_1550_));
 sky130_fd_sc_hd__nand2_2 _4612_ (.A(net97),
    .B(_1550_),
    .Y(_1551_));
 sky130_fd_sc_hd__and2_1 _4613_ (.A(net9),
    .B(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__a21o_1 _4614_ (.A1(net804),
    .A2(net158),
    .B1(net97),
    .X(_1553_));
 sky130_fd_sc_hd__and2_4 _4615_ (.A(_0600_),
    .B(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__nand2_1 _4616_ (.A(net648),
    .B(net412),
    .Y(_1555_));
 sky130_fd_sc_hd__o21ai_4 _4617_ (.A1(net92),
    .A2(_1555_),
    .B1(_1554_),
    .Y(_1556_));
 sky130_fd_sc_hd__o22a_1 _4618_ (.A1(net464),
    .A2(_1554_),
    .B1(_1556_),
    .B2(_1552_),
    .X(_0198_));
 sky130_fd_sc_hd__and2_1 _4619_ (.A(net8),
    .B(_1551_),
    .X(_1557_));
 sky130_fd_sc_hd__o22a_1 _4620_ (.A1(net155),
    .A2(_1554_),
    .B1(_1556_),
    .B2(_1557_),
    .X(_0199_));
 sky130_fd_sc_hd__and2_1 _4621_ (.A(net6),
    .B(_1551_),
    .X(_1558_));
 sky130_fd_sc_hd__o22a_1 _4622_ (.A1(net152),
    .A2(_1554_),
    .B1(_1556_),
    .B2(_1558_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_1 _4623_ (.A(net3),
    .B(_1551_),
    .X(_1559_));
 sky130_fd_sc_hd__o22a_1 _4624_ (.A1(net148),
    .A2(_1554_),
    .B1(_1556_),
    .B2(_1559_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_1 _4625_ (.A(net2),
    .B(_1551_),
    .X(_1560_));
 sky130_fd_sc_hd__o22a_1 _4626_ (.A1(net143),
    .A2(_1554_),
    .B1(_1556_),
    .B2(_1560_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _4627_ (.A(net4),
    .B(_1551_),
    .X(_1561_));
 sky130_fd_sc_hd__o22a_1 _4628_ (.A1(net141),
    .A2(_1554_),
    .B1(_1556_),
    .B2(_1561_),
    .X(_0203_));
 sky130_fd_sc_hd__and2_1 _4629_ (.A(net5),
    .B(_1551_),
    .X(_1562_));
 sky130_fd_sc_hd__o22a_1 _4630_ (.A1(net814),
    .A2(_1554_),
    .B1(_1556_),
    .B2(_1562_),
    .X(_0204_));
 sky130_fd_sc_hd__and2_1 _4631_ (.A(net7),
    .B(_1551_),
    .X(_1563_));
 sky130_fd_sc_hd__o22a_1 _4632_ (.A1(net841),
    .A2(_1554_),
    .B1(_1556_),
    .B2(_1563_),
    .X(_0205_));
 sky130_fd_sc_hd__and4_1 _4633_ (.A(_2855_),
    .B(net535),
    .C(_0788_),
    .D(_0789_),
    .X(_1564_));
 sky130_fd_sc_hd__nand2_2 _4634_ (.A(_2854_),
    .B(_1564_),
    .Y(_1565_));
 sky130_fd_sc_hd__a21oi_4 _4635_ (.A1(_0786_),
    .A2(net70),
    .B1(net121),
    .Y(_1566_));
 sky130_fd_sc_hd__nor2_1 _4636_ (.A(_0863_),
    .B(_1565_),
    .Y(_1567_));
 sky130_fd_sc_hd__or3b_4 _4637_ (.A(_0383_),
    .B(_0542_),
    .C_N(_0684_),
    .X(_1568_));
 sky130_fd_sc_hd__mux2_1 _4638_ (.A0(\z80.tv80s.i_tv80_core.BusA[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[0] ),
    .S(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__and4_4 _4639_ (.A(_2822_),
    .B(net101),
    .C(_0384_),
    .D(_0541_),
    .X(_1570_));
 sky130_fd_sc_hd__mux2_1 _4640_ (.A0(_1569_),
    .A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .S(_1570_),
    .X(_1571_));
 sky130_fd_sc_hd__o21a_1 _4641_ (.A1(_0786_),
    .A2(_1571_),
    .B1(net70),
    .X(_1572_));
 sky130_fd_sc_hd__o32a_1 _4642_ (.A1(net121),
    .A2(_1567_),
    .A3(_1572_),
    .B1(net527),
    .B2(_1566_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_1 _4643_ (.A0(\z80.tv80s.i_tv80_core.BusA[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[1] ),
    .S(_1568_),
    .X(_1573_));
 sky130_fd_sc_hd__mux2_1 _4644_ (.A0(_1573_),
    .A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .S(_1570_),
    .X(_1574_));
 sky130_fd_sc_hd__nor2_1 _4645_ (.A(_1003_),
    .B(net70),
    .Y(_1575_));
 sky130_fd_sc_hd__o21a_1 _4646_ (.A1(_0786_),
    .A2(_1574_),
    .B1(net70),
    .X(_1576_));
 sky130_fd_sc_hd__o32a_1 _4647_ (.A1(net121),
    .A2(_1575_),
    .A3(_1576_),
    .B1(net529),
    .B2(_1566_),
    .X(_0207_));
 sky130_fd_sc_hd__mux2_1 _4648_ (.A0(\z80.tv80s.i_tv80_core.BusA[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[2] ),
    .S(_1568_),
    .X(_1577_));
 sky130_fd_sc_hd__mux2_1 _4649_ (.A0(_1577_),
    .A1(\z80.tv80s.i_tv80_core.BusB[6] ),
    .S(_1570_),
    .X(_1578_));
 sky130_fd_sc_hd__nor2_1 _4650_ (.A(_1053_),
    .B(net70),
    .Y(_1579_));
 sky130_fd_sc_hd__o21a_1 _4651_ (.A1(_0786_),
    .A2(_1578_),
    .B1(net70),
    .X(_1580_));
 sky130_fd_sc_hd__o32a_1 _4652_ (.A1(net121),
    .A2(_1579_),
    .A3(_1580_),
    .B1(net545),
    .B2(_1566_),
    .X(_0208_));
 sky130_fd_sc_hd__nor2_1 _4653_ (.A(_1086_),
    .B(net70),
    .Y(_1581_));
 sky130_fd_sc_hd__mux2_1 _4654_ (.A0(\z80.tv80s.i_tv80_core.BusA[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .S(_1568_),
    .X(_1582_));
 sky130_fd_sc_hd__mux2_1 _4655_ (.A0(_1582_),
    .A1(\z80.tv80s.i_tv80_core.BusB[7] ),
    .S(_1570_),
    .X(_1583_));
 sky130_fd_sc_hd__o21a_1 _4656_ (.A1(_0786_),
    .A2(_1583_),
    .B1(net70),
    .X(_1584_));
 sky130_fd_sc_hd__o32a_1 _4657_ (.A1(net121),
    .A2(_1581_),
    .A3(_1584_),
    .B1(net565),
    .B2(_1566_),
    .X(_0209_));
 sky130_fd_sc_hd__nor2_1 _4658_ (.A(_1140_),
    .B(net70),
    .Y(_1585_));
 sky130_fd_sc_hd__mux2_1 _4659_ (.A0(\z80.tv80s.i_tv80_core.BusB[0] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .S(_1568_),
    .X(_1586_));
 sky130_fd_sc_hd__mux2_1 _4660_ (.A0(_1586_),
    .A1(\z80.tv80s.i_tv80_core.BusA[0] ),
    .S(_1570_),
    .X(_1587_));
 sky130_fd_sc_hd__o21a_1 _4661_ (.A1(_0786_),
    .A2(_1587_),
    .B1(net70),
    .X(_1588_));
 sky130_fd_sc_hd__o32a_1 _4662_ (.A1(net121),
    .A2(_1585_),
    .A3(_1588_),
    .B1(net561),
    .B2(_1566_),
    .X(_0210_));
 sky130_fd_sc_hd__nor2_1 _4663_ (.A(_1177_),
    .B(net70),
    .Y(_1589_));
 sky130_fd_sc_hd__mux2_1 _4664_ (.A0(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .S(_1568_),
    .X(_1590_));
 sky130_fd_sc_hd__mux2_1 _4665_ (.A0(_1590_),
    .A1(\z80.tv80s.i_tv80_core.BusA[1] ),
    .S(_1570_),
    .X(_1591_));
 sky130_fd_sc_hd__o21a_1 _4666_ (.A1(_0786_),
    .A2(_1591_),
    .B1(net70),
    .X(_1592_));
 sky130_fd_sc_hd__o32a_1 _4667_ (.A1(net121),
    .A2(_1589_),
    .A3(_1592_),
    .B1(net572),
    .B2(_1566_),
    .X(_0211_));
 sky130_fd_sc_hd__nor2_1 _4668_ (.A(_1232_),
    .B(net70),
    .Y(_1593_));
 sky130_fd_sc_hd__mux2_1 _4669_ (.A0(\z80.tv80s.i_tv80_core.BusB[2] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[6] ),
    .S(_1568_),
    .X(_1594_));
 sky130_fd_sc_hd__mux2_1 _4670_ (.A0(_1594_),
    .A1(\z80.tv80s.i_tv80_core.BusA[2] ),
    .S(_1570_),
    .X(_1595_));
 sky130_fd_sc_hd__o21a_1 _4671_ (.A1(_0786_),
    .A2(_1595_),
    .B1(net70),
    .X(_1596_));
 sky130_fd_sc_hd__o32a_1 _4672_ (.A1(net121),
    .A2(_1593_),
    .A3(_1596_),
    .B1(net551),
    .B2(_1566_),
    .X(_0212_));
 sky130_fd_sc_hd__nor2_1 _4673_ (.A(_1281_),
    .B(net70),
    .Y(_1597_));
 sky130_fd_sc_hd__mux2_1 _4674_ (.A0(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A1(\z80.tv80s.i_tv80_core.BusB[7] ),
    .S(_1568_),
    .X(_1598_));
 sky130_fd_sc_hd__mux2_1 _4675_ (.A0(_1598_),
    .A1(\z80.tv80s.i_tv80_core.BusA[3] ),
    .S(_1570_),
    .X(_1599_));
 sky130_fd_sc_hd__o21a_1 _4676_ (.A1(_0786_),
    .A2(_1599_),
    .B1(net70),
    .X(_1600_));
 sky130_fd_sc_hd__o32a_1 _4677_ (.A1(net121),
    .A2(_1597_),
    .A3(_1600_),
    .B1(net549),
    .B2(_1566_),
    .X(_0213_));
 sky130_fd_sc_hd__nand2_4 _4678_ (.A(net630),
    .B(_1564_),
    .Y(_1601_));
 sky130_fd_sc_hd__or4_4 _4679_ (.A(_2822_),
    .B(net111),
    .C(_2906_),
    .D(_2950_),
    .X(_1602_));
 sky130_fd_sc_hd__or2_2 _4680_ (.A(net56),
    .B(_1602_),
    .X(_1603_));
 sky130_fd_sc_hd__a21o_2 _4681_ (.A1(_1484_),
    .A2(_1603_),
    .B1(net97),
    .X(_1604_));
 sky130_fd_sc_hd__o22a_1 _4682_ (.A1(\z80.tv80s.i_tv80_core.Ap[0] ),
    .A2(_1484_),
    .B1(_1603_),
    .B2(_2857_),
    .X(_1605_));
 sky130_fd_sc_hd__a2bb2o_1 _4683_ (.A1_N(net97),
    .A2_N(_1605_),
    .B1(_1604_),
    .B2(_2857_),
    .X(_1606_));
 sky130_fd_sc_hd__and3_2 _4684_ (.A(net144),
    .B(net116),
    .C(_1369_),
    .X(_1607_));
 sky130_fd_sc_hd__or3b_4 _4685_ (.A(_2823_),
    .B(_2831_),
    .C_N(_1369_),
    .X(_1608_));
 sky130_fd_sc_hd__mux2_1 _4686_ (.A0(net614),
    .A1(net723),
    .S(_1370_),
    .X(_1609_));
 sky130_fd_sc_hd__o21ai_1 _4687_ (.A1(_1608_),
    .A2(_1609_),
    .B1(_1601_),
    .Y(_1610_));
 sky130_fd_sc_hd__a21o_1 _4688_ (.A1(_1606_),
    .A2(_1608_),
    .B1(_1610_),
    .X(_1611_));
 sky130_fd_sc_hd__o21ai_1 _4689_ (.A1(_0863_),
    .A2(_1601_),
    .B1(_1611_),
    .Y(_1612_));
 sky130_fd_sc_hd__mux2_1 _4690_ (.A0(net866),
    .A1(_1612_),
    .S(net110),
    .X(_0214_));
 sky130_fd_sc_hd__a2bb2o_1 _4691_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2_N(_1603_),
    .B1(_1483_),
    .B2(net670),
    .X(_1613_));
 sky130_fd_sc_hd__a22o_1 _4692_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_1604_),
    .B1(_1613_),
    .B2(net93),
    .X(_1614_));
 sky130_fd_sc_hd__mux2_1 _4693_ (.A0(net594),
    .A1(net578),
    .S(_1370_),
    .X(_1615_));
 sky130_fd_sc_hd__mux2_1 _4694_ (.A0(_1614_),
    .A1(_1615_),
    .S(_1607_),
    .X(_1616_));
 sky130_fd_sc_hd__mux2_1 _4695_ (.A0(_1004_),
    .A1(_1616_),
    .S(_1601_),
    .X(_1617_));
 sky130_fd_sc_hd__mux2_1 _4696_ (.A0(net870),
    .A1(_1617_),
    .S(net108),
    .X(_0215_));
 sky130_fd_sc_hd__mux2_1 _4697_ (.A0(net633),
    .A1(net624),
    .S(_1370_),
    .X(_1618_));
 sky130_fd_sc_hd__a2bb2o_1 _4698_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2_N(_1603_),
    .B1(_1483_),
    .B2(net668),
    .X(_1619_));
 sky130_fd_sc_hd__a22o_1 _4699_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_1604_),
    .B1(_1619_),
    .B2(net92),
    .X(_1620_));
 sky130_fd_sc_hd__mux2_1 _4700_ (.A0(_1618_),
    .A1(_1620_),
    .S(_1608_),
    .X(_1621_));
 sky130_fd_sc_hd__mux2_1 _4701_ (.A0(_1054_),
    .A1(_1621_),
    .S(_1601_),
    .X(_1622_));
 sky130_fd_sc_hd__mux2_1 _4702_ (.A0(net865),
    .A1(_1622_),
    .S(net110),
    .X(_0216_));
 sky130_fd_sc_hd__a2bb2o_1 _4703_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2_N(_1603_),
    .B1(_1483_),
    .B2(net705),
    .X(_1623_));
 sky130_fd_sc_hd__a22o_1 _4704_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_1604_),
    .B1(_1623_),
    .B2(net92),
    .X(_1624_));
 sky130_fd_sc_hd__mux2_1 _4705_ (.A0(net701),
    .A1(net540),
    .S(_1370_),
    .X(_1625_));
 sky130_fd_sc_hd__mux2_1 _4706_ (.A0(_1624_),
    .A1(_1625_),
    .S(_1607_),
    .X(_1626_));
 sky130_fd_sc_hd__mux2_1 _4707_ (.A0(_1087_),
    .A1(_1626_),
    .S(_1601_),
    .X(_1627_));
 sky130_fd_sc_hd__mux2_1 _4708_ (.A0(net879),
    .A1(_1627_),
    .S(net108),
    .X(_0217_));
 sky130_fd_sc_hd__a2bb2o_1 _4709_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2_N(_1603_),
    .B1(_1483_),
    .B2(net693),
    .X(_1628_));
 sky130_fd_sc_hd__a22o_1 _4710_ (.A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(_1604_),
    .B1(_1628_),
    .B2(net93),
    .X(_1629_));
 sky130_fd_sc_hd__mux2_1 _4711_ (.A0(net719),
    .A1(net610),
    .S(_1370_),
    .X(_1630_));
 sky130_fd_sc_hd__mux2_1 _4712_ (.A0(_1629_),
    .A1(_1630_),
    .S(_1607_),
    .X(_1631_));
 sky130_fd_sc_hd__mux2_1 _4713_ (.A0(_1141_),
    .A1(_1631_),
    .S(_1601_),
    .X(_1632_));
 sky130_fd_sc_hd__mux2_1 _4714_ (.A0(net863),
    .A1(_1632_),
    .S(net110),
    .X(_0218_));
 sky130_fd_sc_hd__a2bb2o_1 _4715_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2_N(_1603_),
    .B1(_1483_),
    .B2(net683),
    .X(_1633_));
 sky130_fd_sc_hd__a22o_1 _4716_ (.A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2(_1604_),
    .B1(_1633_),
    .B2(net92),
    .X(_1634_));
 sky130_fd_sc_hd__mux2_1 _4717_ (.A0(net751),
    .A1(net586),
    .S(_1370_),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _4718_ (.A0(_1634_),
    .A1(_1635_),
    .S(_1607_),
    .X(_1636_));
 sky130_fd_sc_hd__mux2_1 _4719_ (.A0(_1178_),
    .A1(_1636_),
    .S(_1601_),
    .X(_1637_));
 sky130_fd_sc_hd__mux2_1 _4720_ (.A0(net875),
    .A1(_1637_),
    .S(net108),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_1 _4721_ (.A0(net622),
    .A1(net608),
    .S(_1370_),
    .X(_1638_));
 sky130_fd_sc_hd__a2bb2o_1 _4722_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2_N(_1603_),
    .B1(_1483_),
    .B2(net660),
    .X(_1639_));
 sky130_fd_sc_hd__a22o_1 _4723_ (.A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_1604_),
    .B1(_1639_),
    .B2(net92),
    .X(_1640_));
 sky130_fd_sc_hd__mux2_1 _4724_ (.A0(_1638_),
    .A1(_1640_),
    .S(_1608_),
    .X(_1641_));
 sky130_fd_sc_hd__mux2_1 _4725_ (.A0(_1233_),
    .A1(_1641_),
    .S(_1601_),
    .X(_1642_));
 sky130_fd_sc_hd__mux2_1 _4726_ (.A0(net864),
    .A1(_1642_),
    .S(net108),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_1 _4727_ (.A0(net777),
    .A1(net374),
    .S(_1370_),
    .X(_1643_));
 sky130_fd_sc_hd__a2bb2o_1 _4728_ (.A1_N(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2_N(_1603_),
    .B1(_1483_),
    .B2(net662),
    .X(_1644_));
 sky130_fd_sc_hd__a22o_1 _4729_ (.A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(_1604_),
    .B1(_1644_),
    .B2(net92),
    .X(_1645_));
 sky130_fd_sc_hd__mux2_1 _4730_ (.A0(_1643_),
    .A1(_1645_),
    .S(_1608_),
    .X(_1646_));
 sky130_fd_sc_hd__mux2_1 _4731_ (.A0(_1282_),
    .A1(_1646_),
    .S(_1601_),
    .X(_1647_));
 sky130_fd_sc_hd__mux2_1 _4732_ (.A0(net836),
    .A1(_1647_),
    .S(net110),
    .X(_0221_));
 sky130_fd_sc_hd__a21oi_2 _4733_ (.A1(net56),
    .A2(net93),
    .B1(_0603_),
    .Y(_1648_));
 sky130_fd_sc_hd__and3b_1 _4734_ (.A_N(_0469_),
    .B(_0513_),
    .C(_0408_),
    .X(_1649_));
 sky130_fd_sc_hd__a2bb2o_1 _4735_ (.A1_N(_0419_),
    .A2_N(_0656_),
    .B1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .B2(_2988_),
    .X(_1650_));
 sky130_fd_sc_hd__a211o_1 _4736_ (.A1(_0632_),
    .A2(_0868_),
    .B1(_1649_),
    .C1(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__a21o_4 _4737_ (.A1(net161),
    .A2(_1651_),
    .B1(_0738_),
    .X(_1652_));
 sky130_fd_sc_hd__inv_2 _4738_ (.A(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__mux4_1 _4739_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .S0(net164),
    .S1(net133),
    .X(_1654_));
 sky130_fd_sc_hd__mux4_1 _4740_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .S0(net164),
    .S1(net133),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_4 _4741_ (.A0(_1655_),
    .A1(_1654_),
    .S(net165),
    .X(_1656_));
 sky130_fd_sc_hd__o21a_1 _4742_ (.A1(net79),
    .A2(_1656_),
    .B1(net67),
    .X(_1657_));
 sky130_fd_sc_hd__or4_1 _4743_ (.A(_0425_),
    .B(_0506_),
    .C(_0708_),
    .D(_1408_),
    .X(_1658_));
 sky130_fd_sc_hd__and3_1 _4744_ (.A(net155),
    .B(net152),
    .C(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(_1659_));
 sky130_fd_sc_hd__or4b_2 _4745_ (.A(net111),
    .B(_0656_),
    .C(_1658_),
    .D_N(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__inv_2 _4746_ (.A(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__and4bb_1 _4747_ (.A_N(_2924_),
    .B_N(_2939_),
    .C(_2987_),
    .D(_0426_),
    .X(_1662_));
 sky130_fd_sc_hd__and4bb_1 _4748_ (.A_N(_0409_),
    .B_N(_0410_),
    .C(_1409_),
    .D(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__a41o_2 _4749_ (.A1(net162),
    .A2(_0706_),
    .A3(_0867_),
    .A4(_1663_),
    .B1(_1661_),
    .X(_1664_));
 sky130_fd_sc_hd__and2_2 _4750_ (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .B(_0725_),
    .X(_1665_));
 sky130_fd_sc_hd__nor2_1 _4751_ (.A(net63),
    .B(_1665_),
    .Y(_1666_));
 sky130_fd_sc_hd__and3_2 _4752_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .B(\z80.tv80s.i_tv80_core.IntCycle ),
    .C(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .X(_1667_));
 sky130_fd_sc_hd__nand3_2 _4753_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .B(\z80.tv80s.i_tv80_core.IntCycle ),
    .C(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .Y(_1668_));
 sky130_fd_sc_hd__and2_4 _4754_ (.A(_0453_),
    .B(_0492_),
    .X(_1669_));
 sky130_fd_sc_hd__nand2_2 _4755_ (.A(_0453_),
    .B(_0492_),
    .Y(_1670_));
 sky130_fd_sc_hd__nor3_4 _4756_ (.A(_0437_),
    .B(_0452_),
    .C(_0492_),
    .Y(_1671_));
 sky130_fd_sc_hd__nor2_8 _4757_ (.A(_0438_),
    .B(_0492_),
    .Y(_1672_));
 sky130_fd_sc_hd__and3b_4 _4758_ (.A_N(_0492_),
    .B(_0438_),
    .C(_0452_),
    .X(_1673_));
 sky130_fd_sc_hd__a22o_1 _4759_ (.A1(_1656_),
    .A2(_1672_),
    .B1(_1673_),
    .B2(\z80.tv80s.di_reg[0] ),
    .X(_1674_));
 sky130_fd_sc_hd__a21o_1 _4760_ (.A1(\z80.tv80s.i_tv80_core.SP[0] ),
    .A2(_1671_),
    .B1(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__mux2_1 _4761_ (.A0(\z80.tv80s.i_tv80_core.PC[0] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1676_));
 sky130_fd_sc_hd__mux2_1 _4762_ (.A0(_1656_),
    .A1(_1676_),
    .S(_0497_),
    .X(_1677_));
 sky130_fd_sc_hd__and2b_4 _4763_ (.A_N(_0439_),
    .B(_0493_),
    .X(_1678_));
 sky130_fd_sc_hd__a2111o_1 _4764_ (.A1(_2870_),
    .A2(_2939_),
    .B1(_0709_),
    .C1(_1658_),
    .D1(_2924_),
    .X(_1679_));
 sky130_fd_sc_hd__or2_1 _4765_ (.A(_2938_),
    .B(_0703_),
    .X(_1680_));
 sky130_fd_sc_hd__inv_2 _4766_ (.A(_1680_),
    .Y(_1681_));
 sky130_fd_sc_hd__and3_1 _4767_ (.A(net161),
    .B(_0541_),
    .C(_0704_),
    .X(_1682_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_0702_),
    .B(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__or4_2 _4769_ (.A(_0699_),
    .B(_1679_),
    .C(_1680_),
    .D(_1683_),
    .X(_1684_));
 sky130_fd_sc_hd__o21ai_4 _4770_ (.A1(_0542_),
    .A2(_0634_),
    .B1(_1684_),
    .Y(_1685_));
 sky130_fd_sc_hd__a31o_1 _4771_ (.A1(_2825_),
    .A2(_0388_),
    .A3(_0540_),
    .B1(_0383_),
    .X(_1686_));
 sky130_fd_sc_hd__nor2_1 _4772_ (.A(_0699_),
    .B(_1679_),
    .Y(_1687_));
 sky130_fd_sc_hd__a41o_1 _4773_ (.A1(_0702_),
    .A2(_1681_),
    .A3(_1682_),
    .A4(_1687_),
    .B1(net101),
    .X(_1688_));
 sky130_fd_sc_hd__nand2_1 _4774_ (.A(_1686_),
    .B(_1688_),
    .Y(_1689_));
 sky130_fd_sc_hd__xor2_1 _4775_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(_1685_),
    .X(_1690_));
 sky130_fd_sc_hd__a22o_1 _4776_ (.A1(net57),
    .A2(_1677_),
    .B1(_1678_),
    .B2(_1690_),
    .X(_1691_));
 sky130_fd_sc_hd__a211o_1 _4777_ (.A1(\z80.tv80s.i_tv80_core.PC[0] ),
    .A2(_1669_),
    .B1(_1675_),
    .C1(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A1(_1692_),
    .S(net90),
    .X(_1693_));
 sky130_fd_sc_hd__a221o_1 _4779_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(net63),
    .B1(net61),
    .B2(_1693_),
    .C1(net80),
    .X(_1694_));
 sky130_fd_sc_hd__a221o_1 _4780_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(_1652_),
    .B1(_1657_),
    .B2(_1694_),
    .C1(net97),
    .X(_1695_));
 sky130_fd_sc_hd__o21a_1 _4781_ (.A1(\z80.tv80s.i_tv80_core.R[0] ),
    .A2(net91),
    .B1(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__mux2_1 _4782_ (.A0(net547),
    .A1(_1696_),
    .S(net55),
    .X(_0222_));
 sky130_fd_sc_hd__a21o_1 _4783_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .A2(_1667_),
    .B1(_1665_),
    .X(_1697_));
 sky130_fd_sc_hd__mux4_1 _4784_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .S0(net164),
    .S1(net133),
    .X(_1698_));
 sky130_fd_sc_hd__mux4_1 _4785_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .S0(net164),
    .S1(net133),
    .X(_1699_));
 sky130_fd_sc_hd__mux2_2 _4786_ (.A0(_1699_),
    .A1(_1698_),
    .S(net165),
    .X(_1700_));
 sky130_fd_sc_hd__mux2_1 _4787_ (.A0(\z80.tv80s.i_tv80_core.PC[1] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(_0499_),
    .X(_1701_));
 sky130_fd_sc_hd__or2_1 _4788_ (.A(net98),
    .B(_1700_),
    .X(_1702_));
 sky130_fd_sc_hd__o211a_1 _4789_ (.A1(_0496_),
    .A2(_1701_),
    .B1(_1702_),
    .C1(net57),
    .X(_1703_));
 sky130_fd_sc_hd__a21o_1 _4790_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(_1685_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .X(_1704_));
 sky130_fd_sc_hd__and2_1 _4791_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .X(_1705_));
 sky130_fd_sc_hd__and2_1 _4792_ (.A(_1685_),
    .B(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__and3b_1 _4793_ (.A_N(_1706_),
    .B(_1678_),
    .C(_1704_),
    .X(_1707_));
 sky130_fd_sc_hd__a221o_1 _4794_ (.A1(\z80.tv80s.i_tv80_core.SP[1] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(_1700_),
    .C1(_1669_),
    .X(_1708_));
 sky130_fd_sc_hd__a2111o_1 _4795_ (.A1(\z80.tv80s.di_reg[1] ),
    .A2(_1673_),
    .B1(_1703_),
    .C1(_1707_),
    .D1(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__or2_1 _4796_ (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .B(_1670_),
    .X(_1710_));
 sky130_fd_sc_hd__a31o_1 _4797_ (.A1(net90),
    .A2(_1709_),
    .A3(_1710_),
    .B1(_1697_),
    .X(_1711_));
 sky130_fd_sc_hd__mux2_1 _4798_ (.A0(_1711_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net63),
    .X(_1712_));
 sky130_fd_sc_hd__nand2_1 _4799_ (.A(net79),
    .B(_1712_),
    .Y(_1713_));
 sky130_fd_sc_hd__a21oi_1 _4800_ (.A1(net80),
    .A2(_1700_),
    .B1(_1652_),
    .Y(_1714_));
 sky130_fd_sc_hd__a221o_1 _4801_ (.A1(_2861_),
    .A2(_1652_),
    .B1(_1713_),
    .B2(_1714_),
    .C1(net97),
    .X(_1715_));
 sky130_fd_sc_hd__a21bo_1 _4802_ (.A1(net578),
    .A2(net95),
    .B1_N(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__mux2_1 _4803_ (.A0(net590),
    .A1(_1716_),
    .S(net55),
    .X(_0223_));
 sky130_fd_sc_hd__a21o_1 _4804_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .A2(_1667_),
    .B1(_1665_),
    .X(_1717_));
 sky130_fd_sc_hd__mux4_1 _4805_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .S0(net133),
    .S1(net164),
    .X(_1718_));
 sky130_fd_sc_hd__mux4_1 _4806_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .S0(net133),
    .S1(net164),
    .X(_1719_));
 sky130_fd_sc_hd__mux2_4 _4807_ (.A0(_1719_),
    .A1(_1718_),
    .S(net165),
    .X(_1720_));
 sky130_fd_sc_hd__or2_1 _4808_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B(_1706_),
    .X(_1721_));
 sky130_fd_sc_hd__or3b_1 _4809_ (.A(_2862_),
    .B(_1689_),
    .C_N(_1705_),
    .X(_1722_));
 sky130_fd_sc_hd__mux2_1 _4810_ (.A0(\z80.tv80s.i_tv80_core.PC[2] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1723_));
 sky130_fd_sc_hd__mux2_1 _4811_ (.A0(_1720_),
    .A1(_1723_),
    .S(net98),
    .X(_1724_));
 sky130_fd_sc_hd__a221o_1 _4812_ (.A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .A2(net58),
    .B1(_1672_),
    .B2(_1720_),
    .C1(_1669_),
    .X(_1725_));
 sky130_fd_sc_hd__a22o_1 _4813_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_1673_),
    .B1(_1724_),
    .B2(net57),
    .X(_1726_));
 sky130_fd_sc_hd__a31o_1 _4814_ (.A1(_1678_),
    .A2(_1721_),
    .A3(_1722_),
    .B1(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__o22a_1 _4815_ (.A1(\z80.tv80s.i_tv80_core.PC[2] ),
    .A2(_1670_),
    .B1(_1725_),
    .B2(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__a21o_1 _4816_ (.A1(net90),
    .A2(_1728_),
    .B1(_1717_),
    .X(_1729_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(_1729_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(net63),
    .X(_1730_));
 sky130_fd_sc_hd__nand2_1 _4818_ (.A(net79),
    .B(_1730_),
    .Y(_1731_));
 sky130_fd_sc_hd__a21oi_1 _4819_ (.A1(net80),
    .A2(_1720_),
    .B1(_1652_),
    .Y(_1732_));
 sky130_fd_sc_hd__a221o_1 _4820_ (.A1(_2862_),
    .A2(_1652_),
    .B1(_1731_),
    .B2(_1732_),
    .C1(net95),
    .X(_1733_));
 sky130_fd_sc_hd__o21ai_1 _4821_ (.A1(_2858_),
    .A2(net91),
    .B1(_1733_),
    .Y(_1734_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(net555),
    .A1(_1734_),
    .S(net55),
    .X(_0224_));
 sky130_fd_sc_hd__mux4_1 _4823_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .S0(net133),
    .S1(net164),
    .X(_1735_));
 sky130_fd_sc_hd__mux4_1 _4824_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .S0(net133),
    .S1(net164),
    .X(_1736_));
 sky130_fd_sc_hd__mux2_4 _4825_ (.A0(_1736_),
    .A1(_1735_),
    .S(net165),
    .X(_1737_));
 sky130_fd_sc_hd__a21o_1 _4826_ (.A1(net80),
    .A2(_1737_),
    .B1(_1652_),
    .X(_1738_));
 sky130_fd_sc_hd__and3_1 _4827_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .C(_1706_),
    .X(_1739_));
 sky130_fd_sc_hd__xnor2_1 _4828_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .B(_1722_),
    .Y(_1740_));
 sky130_fd_sc_hd__mux2_1 _4829_ (.A0(\z80.tv80s.i_tv80_core.PC[3] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .S(_0499_),
    .X(_1741_));
 sky130_fd_sc_hd__or2_1 _4830_ (.A(net98),
    .B(_1737_),
    .X(_1742_));
 sky130_fd_sc_hd__o211a_1 _4831_ (.A1(_0496_),
    .A2(_1741_),
    .B1(_1742_),
    .C1(net57),
    .X(_1743_));
 sky130_fd_sc_hd__a221o_1 _4832_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(_1737_),
    .C1(_1669_),
    .X(_1744_));
 sky130_fd_sc_hd__a221o_1 _4833_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_1673_),
    .B1(_1678_),
    .B2(_1740_),
    .C1(_1743_),
    .X(_1745_));
 sky130_fd_sc_hd__o22a_1 _4834_ (.A1(\z80.tv80s.i_tv80_core.PC[3] ),
    .A2(_1670_),
    .B1(_1744_),
    .B2(_1745_),
    .X(_1746_));
 sky130_fd_sc_hd__mux2_1 _4835_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A1(_1746_),
    .S(net90),
    .X(_1747_));
 sky130_fd_sc_hd__a22o_1 _4836_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net63),
    .B1(net61),
    .B2(_1747_),
    .X(_1748_));
 sky130_fd_sc_hd__a21o_1 _4837_ (.A1(net79),
    .A2(_1748_),
    .B1(_1738_),
    .X(_1749_));
 sky130_fd_sc_hd__o211a_1 _4838_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net67),
    .B1(_1749_),
    .C1(net91),
    .X(_1750_));
 sky130_fd_sc_hd__a21bo_1 _4839_ (.A1(net540),
    .A2(net95),
    .B1_N(net55),
    .X(_1751_));
 sky130_fd_sc_hd__o22a_1 _4840_ (.A1(net602),
    .A2(net55),
    .B1(_1750_),
    .B2(_1751_),
    .X(_0225_));
 sky130_fd_sc_hd__mux4_1 _4841_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .S0(net132),
    .S1(net163),
    .X(_1752_));
 sky130_fd_sc_hd__mux4_1 _4842_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .S0(net132),
    .S1(net163),
    .X(_1753_));
 sky130_fd_sc_hd__mux2_4 _4843_ (.A0(_1753_),
    .A1(_1752_),
    .S(net165),
    .X(_1754_));
 sky130_fd_sc_hd__a21o_1 _4844_ (.A1(net80),
    .A2(_1754_),
    .B1(_1652_),
    .X(_1755_));
 sky130_fd_sc_hd__or2_1 _4845_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .B(_1739_),
    .X(_1756_));
 sky130_fd_sc_hd__and2_1 _4846_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .B(_1739_),
    .X(_1757_));
 sky130_fd_sc_hd__and3b_1 _4847_ (.A_N(_1757_),
    .B(_1678_),
    .C(_1756_),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _4848_ (.A0(\z80.tv80s.i_tv80_core.PC[4] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1759_));
 sky130_fd_sc_hd__mux2_1 _4849_ (.A0(_1754_),
    .A1(_1759_),
    .S(net98),
    .X(_1760_));
 sky130_fd_sc_hd__a221o_1 _4850_ (.A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(_1754_),
    .C1(_1669_),
    .X(_1761_));
 sky130_fd_sc_hd__a22o_1 _4851_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_1673_),
    .B1(_1760_),
    .B2(net57),
    .X(_1762_));
 sky130_fd_sc_hd__or3_1 _4852_ (.A(_1758_),
    .B(_1761_),
    .C(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__o21a_1 _4853_ (.A1(\z80.tv80s.i_tv80_core.PC[4] ),
    .A2(_1670_),
    .B1(net89),
    .X(_1764_));
 sky130_fd_sc_hd__a22o_1 _4854_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(_1667_),
    .B1(_1763_),
    .B2(_1764_),
    .X(_1765_));
 sky130_fd_sc_hd__a22o_1 _4855_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net62),
    .B1(net61),
    .B2(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__a21o_1 _4856_ (.A1(net79),
    .A2(_1766_),
    .B1(_1755_),
    .X(_1767_));
 sky130_fd_sc_hd__o211a_1 _4857_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net67),
    .B1(_1767_),
    .C1(net91),
    .X(_1768_));
 sky130_fd_sc_hd__a21bo_1 _4858_ (.A1(\z80.tv80s.i_tv80_core.R[4] ),
    .A2(net95),
    .B1_N(net55),
    .X(_1769_));
 sky130_fd_sc_hd__o22a_1 _4859_ (.A1(net536),
    .A2(net55),
    .B1(_1768_),
    .B2(_1769_),
    .X(_0226_));
 sky130_fd_sc_hd__mux4_1 _4860_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .S0(net132),
    .S1(net163),
    .X(_1770_));
 sky130_fd_sc_hd__mux4_1 _4861_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .S0(net132),
    .S1(net163),
    .X(_1771_));
 sky130_fd_sc_hd__mux2_2 _4862_ (.A0(_1771_),
    .A1(_1770_),
    .S(net165),
    .X(_1772_));
 sky130_fd_sc_hd__nand2_1 _4863_ (.A(net80),
    .B(_1772_),
    .Y(_1773_));
 sky130_fd_sc_hd__a21o_1 _4864_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A2(_1667_),
    .B1(_1665_),
    .X(_1774_));
 sky130_fd_sc_hd__or2_1 _4865_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .B(_1757_),
    .X(_1775_));
 sky130_fd_sc_hd__and2_1 _4866_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .B(_1757_),
    .X(_1776_));
 sky130_fd_sc_hd__and3b_1 _4867_ (.A_N(_1776_),
    .B(_1678_),
    .C(_1775_),
    .X(_1777_));
 sky130_fd_sc_hd__mux2_1 _4868_ (.A0(\z80.tv80s.i_tv80_core.PC[5] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1778_));
 sky130_fd_sc_hd__mux2_1 _4869_ (.A0(_1772_),
    .A1(_1778_),
    .S(net98),
    .X(_1779_));
 sky130_fd_sc_hd__a221o_1 _4870_ (.A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(_1772_),
    .C1(_1669_),
    .X(_1780_));
 sky130_fd_sc_hd__a22o_1 _4871_ (.A1(\z80.tv80s.di_reg[5] ),
    .A2(_1673_),
    .B1(_1779_),
    .B2(net57),
    .X(_1781_));
 sky130_fd_sc_hd__o32a_1 _4872_ (.A1(_1777_),
    .A2(_1780_),
    .A3(_1781_),
    .B1(_1670_),
    .B2(\z80.tv80s.i_tv80_core.PC[5] ),
    .X(_1782_));
 sky130_fd_sc_hd__a21o_1 _4873_ (.A1(net90),
    .A2(_1782_),
    .B1(_1774_),
    .X(_1783_));
 sky130_fd_sc_hd__mux2_1 _4874_ (.A0(_1783_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net63),
    .X(_1784_));
 sky130_fd_sc_hd__a21bo_1 _4875_ (.A1(net79),
    .A2(_1784_),
    .B1_N(_1773_),
    .X(_1785_));
 sky130_fd_sc_hd__mux2_1 _4876_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A1(_1785_),
    .S(net67),
    .X(_1786_));
 sky130_fd_sc_hd__mux2_1 _4877_ (.A0(net586),
    .A1(_1786_),
    .S(net93),
    .X(_1787_));
 sky130_fd_sc_hd__mux2_1 _4878_ (.A0(net598),
    .A1(_1787_),
    .S(net55),
    .X(_0227_));
 sky130_fd_sc_hd__mux4_1 _4879_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .S0(net133),
    .S1(net164),
    .X(_1788_));
 sky130_fd_sc_hd__mux4_1 _4880_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .S0(net133),
    .S1(net164),
    .X(_1789_));
 sky130_fd_sc_hd__mux2_2 _4881_ (.A0(_1789_),
    .A1(_1788_),
    .S(net165),
    .X(_1790_));
 sky130_fd_sc_hd__nand2_1 _4882_ (.A(net80),
    .B(_1790_),
    .Y(_1791_));
 sky130_fd_sc_hd__a21o_1 _4883_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A2(_1667_),
    .B1(_1665_),
    .X(_1792_));
 sky130_fd_sc_hd__mux2_1 _4884_ (.A0(\z80.tv80s.i_tv80_core.PC[6] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(_0499_),
    .X(_1793_));
 sky130_fd_sc_hd__mux2_1 _4885_ (.A0(_1790_),
    .A1(_1793_),
    .S(net98),
    .X(_1794_));
 sky130_fd_sc_hd__a21boi_1 _4886_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A2(_1776_),
    .B1_N(_1678_),
    .Y(_1795_));
 sky130_fd_sc_hd__o21a_1 _4887_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A2(_1776_),
    .B1(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__a221o_1 _4888_ (.A1(\z80.tv80s.i_tv80_core.SP[6] ),
    .A2(net58),
    .B1(_1672_),
    .B2(_1790_),
    .C1(_1669_),
    .X(_1797_));
 sky130_fd_sc_hd__a22o_1 _4889_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_1673_),
    .B1(_1794_),
    .B2(net57),
    .X(_1798_));
 sky130_fd_sc_hd__o32a_1 _4890_ (.A1(_1796_),
    .A2(_1797_),
    .A3(_1798_),
    .B1(_1670_),
    .B2(\z80.tv80s.i_tv80_core.PC[6] ),
    .X(_1799_));
 sky130_fd_sc_hd__a21o_1 _4891_ (.A1(net90),
    .A2(_1799_),
    .B1(_1792_),
    .X(_1800_));
 sky130_fd_sc_hd__mux2_1 _4892_ (.A0(_1800_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net63),
    .X(_1801_));
 sky130_fd_sc_hd__a21bo_1 _4893_ (.A1(net79),
    .A2(_1801_),
    .B1_N(_1791_),
    .X(_1802_));
 sky130_fd_sc_hd__mux2_1 _4894_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A1(_1802_),
    .S(net67),
    .X(_1803_));
 sky130_fd_sc_hd__mux2_1 _4895_ (.A0(\z80.tv80s.i_tv80_core.R[6] ),
    .A1(_1803_),
    .S(net93),
    .X(_1804_));
 sky130_fd_sc_hd__mux2_1 _4896_ (.A0(net588),
    .A1(_1804_),
    .S(_1648_),
    .X(_0228_));
 sky130_fd_sc_hd__mux4_1 _4897_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .S0(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .S1(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(_1805_));
 sky130_fd_sc_hd__mux4_1 _4898_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .S0(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .S1(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(_1806_));
 sky130_fd_sc_hd__mux2_2 _4899_ (.A0(_1806_),
    .A1(_1805_),
    .S(\z80.tv80s.i_tv80_core.RegAddrC[2] ),
    .X(_1807_));
 sky130_fd_sc_hd__nand2_1 _4900_ (.A(net80),
    .B(_1807_),
    .Y(_1808_));
 sky130_fd_sc_hd__mux2_1 _4901_ (.A0(\z80.tv80s.i_tv80_core.PC[7] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .S(_0499_),
    .X(_1809_));
 sky130_fd_sc_hd__mux2_1 _4902_ (.A0(_1807_),
    .A1(_1809_),
    .S(net98),
    .X(_1810_));
 sky130_fd_sc_hd__a31o_1 _4903_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A2(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A3(_1757_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(_1811_));
 sky130_fd_sc_hd__and4_1 _4904_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .C(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .D(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(_1812_));
 sky130_fd_sc_hd__and4_2 _4905_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .C(_1705_),
    .D(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__inv_2 _4906_ (.A(_1813_),
    .Y(_1814_));
 sky130_fd_sc_hd__o211a_1 _4907_ (.A1(_1689_),
    .A2(_1814_),
    .B1(_1811_),
    .C1(_1678_),
    .X(_1815_));
 sky130_fd_sc_hd__a221o_1 _4908_ (.A1(\z80.tv80s.i_tv80_core.SP[7] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(_1807_),
    .C1(_1669_),
    .X(_1816_));
 sky130_fd_sc_hd__a221o_1 _4909_ (.A1(\z80.tv80s.di_reg[7] ),
    .A2(_1673_),
    .B1(_1810_),
    .B2(_0494_),
    .C1(_1815_),
    .X(_1817_));
 sky130_fd_sc_hd__o22a_1 _4910_ (.A1(\z80.tv80s.i_tv80_core.PC[7] ),
    .A2(_1670_),
    .B1(_1816_),
    .B2(_1817_),
    .X(_1818_));
 sky130_fd_sc_hd__mux2_1 _4911_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(_1818_),
    .S(net90),
    .X(_1819_));
 sky130_fd_sc_hd__a22o_1 _4912_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A2(net63),
    .B1(net61),
    .B2(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__a21bo_1 _4913_ (.A1(net79),
    .A2(_1820_),
    .B1_N(_1808_),
    .X(_1821_));
 sky130_fd_sc_hd__mux2_1 _4914_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(_1821_),
    .S(net67),
    .X(_1822_));
 sky130_fd_sc_hd__mux2_1 _4915_ (.A0(net374),
    .A1(_1822_),
    .S(net93),
    .X(_1823_));
 sky130_fd_sc_hd__mux2_1 _4916_ (.A0(net563),
    .A1(_1823_),
    .S(_1648_),
    .X(_0229_));
 sky130_fd_sc_hd__mux4_1 _4917_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .S0(net163),
    .S1(net132),
    .X(_1824_));
 sky130_fd_sc_hd__mux4_1 _4918_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .S0(net163),
    .S1(net133),
    .X(_1825_));
 sky130_fd_sc_hd__mux2_2 _4919_ (.A0(_1825_),
    .A1(_1824_),
    .S(net165),
    .X(_1826_));
 sky130_fd_sc_hd__nand2_1 _4920_ (.A(net80),
    .B(_1826_),
    .Y(_1827_));
 sky130_fd_sc_hd__a22o_1 _4921_ (.A1(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A2(_1673_),
    .B1(_1826_),
    .B2(_1672_),
    .X(_1828_));
 sky130_fd_sc_hd__a21o_1 _4922_ (.A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .A2(net58),
    .B1(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__mux2_1 _4923_ (.A0(\z80.tv80s.i_tv80_core.PC[8] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1830_));
 sky130_fd_sc_hd__mux2_1 _4924_ (.A0(_1826_),
    .A1(_1830_),
    .S(net98),
    .X(_1831_));
 sky130_fd_sc_hd__xor2_1 _4925_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .B(_1813_),
    .X(_1832_));
 sky130_fd_sc_hd__mux2_1 _4926_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_1832_),
    .S(_1685_),
    .X(_1833_));
 sky130_fd_sc_hd__a22o_1 _4927_ (.A1(net57),
    .A2(_1831_),
    .B1(_1833_),
    .B2(_1678_),
    .X(_1834_));
 sky130_fd_sc_hd__a211o_1 _4928_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(_1669_),
    .B1(_1829_),
    .C1(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_1 _4929_ (.A0(\z80.tv80s.i_tv80_core.I[0] ),
    .A1(_1835_),
    .S(net89),
    .X(_1836_));
 sky130_fd_sc_hd__a22o_1 _4930_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .A2(net63),
    .B1(net60),
    .B2(_1836_),
    .X(_1837_));
 sky130_fd_sc_hd__a21bo_1 _4931_ (.A1(net79),
    .A2(_1837_),
    .B1_N(_1827_),
    .X(_1838_));
 sky130_fd_sc_hd__mux2_1 _4932_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_1838_),
    .S(net66),
    .X(_1839_));
 sky130_fd_sc_hd__mux2_1 _4933_ (.A0(net614),
    .A1(_1839_),
    .S(net91),
    .X(_1840_));
 sky130_fd_sc_hd__mux2_1 _4934_ (.A0(net644),
    .A1(_1840_),
    .S(net55),
    .X(_0230_));
 sky130_fd_sc_hd__mux4_1 _4935_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .S0(net132),
    .S1(net163),
    .X(_1841_));
 sky130_fd_sc_hd__mux4_1 _4936_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .S0(net132),
    .S1(net163),
    .X(_1842_));
 sky130_fd_sc_hd__mux2_2 _4937_ (.A0(_1842_),
    .A1(_1841_),
    .S(net165),
    .X(_1843_));
 sky130_fd_sc_hd__nand2_1 _4938_ (.A(net80),
    .B(_1843_),
    .Y(_1844_));
 sky130_fd_sc_hd__a22o_1 _4939_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_1673_),
    .B1(_1843_),
    .B2(_1672_),
    .X(_1845_));
 sky130_fd_sc_hd__a21o_1 _4940_ (.A1(\z80.tv80s.i_tv80_core.SP[9] ),
    .A2(net58),
    .B1(_1845_),
    .X(_1846_));
 sky130_fd_sc_hd__mux2_1 _4941_ (.A0(\z80.tv80s.i_tv80_core.PC[9] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1847_));
 sky130_fd_sc_hd__mux2_1 _4942_ (.A0(_1843_),
    .A1(_1847_),
    .S(net98),
    .X(_1848_));
 sky130_fd_sc_hd__and3_1 _4943_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .C(_1813_),
    .X(_1849_));
 sky130_fd_sc_hd__a21oi_1 _4944_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .A2(_1813_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .Y(_1850_));
 sky130_fd_sc_hd__nor2_1 _4945_ (.A(_1849_),
    .B(_1850_),
    .Y(_1851_));
 sky130_fd_sc_hd__mux2_1 _4946_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_1851_),
    .S(_1685_),
    .X(_1852_));
 sky130_fd_sc_hd__a22o_1 _4947_ (.A1(net57),
    .A2(_1848_),
    .B1(_1852_),
    .B2(_1678_),
    .X(_1853_));
 sky130_fd_sc_hd__a211o_1 _4948_ (.A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .A2(_1669_),
    .B1(_1846_),
    .C1(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__mux2_1 _4949_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(_1854_),
    .S(net89),
    .X(_1855_));
 sky130_fd_sc_hd__a22o_1 _4950_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .A2(net62),
    .B1(net60),
    .B2(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__a21bo_1 _4951_ (.A1(net78),
    .A2(_1856_),
    .B1_N(_1844_),
    .X(_1857_));
 sky130_fd_sc_hd__mux2_1 _4952_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_1857_),
    .S(net66),
    .X(_1858_));
 sky130_fd_sc_hd__mux2_1 _4953_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(_1858_),
    .S(net91),
    .X(_1859_));
 sky130_fd_sc_hd__mux2_1 _4954_ (.A0(net557),
    .A1(_1859_),
    .S(net55),
    .X(_0231_));
 sky130_fd_sc_hd__mux4_1 _4955_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .S0(net132),
    .S1(net163),
    .X(_1860_));
 sky130_fd_sc_hd__mux4_1 _4956_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .S0(net132),
    .S1(net163),
    .X(_1861_));
 sky130_fd_sc_hd__mux2_2 _4957_ (.A0(_1861_),
    .A1(_1860_),
    .S(net165),
    .X(_1862_));
 sky130_fd_sc_hd__nand2_1 _4958_ (.A(net80),
    .B(_1862_),
    .Y(_1863_));
 sky130_fd_sc_hd__a22o_1 _4959_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_1673_),
    .B1(_1862_),
    .B2(_1672_),
    .X(_1864_));
 sky130_fd_sc_hd__a21o_1 _4960_ (.A1(\z80.tv80s.i_tv80_core.SP[10] ),
    .A2(net58),
    .B1(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__mux2_1 _4961_ (.A0(\z80.tv80s.i_tv80_core.PC[10] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1866_));
 sky130_fd_sc_hd__mux2_1 _4962_ (.A0(_1862_),
    .A1(_1866_),
    .S(net98),
    .X(_1867_));
 sky130_fd_sc_hd__xor2_1 _4963_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .B(_1849_),
    .X(_1868_));
 sky130_fd_sc_hd__mux2_1 _4964_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_1868_),
    .S(_1685_),
    .X(_1869_));
 sky130_fd_sc_hd__a22o_1 _4965_ (.A1(net57),
    .A2(_1867_),
    .B1(_1869_),
    .B2(_1678_),
    .X(_1870_));
 sky130_fd_sc_hd__a211o_1 _4966_ (.A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .A2(_1669_),
    .B1(_1865_),
    .C1(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__mux2_1 _4967_ (.A0(\z80.tv80s.i_tv80_core.I[2] ),
    .A1(_1871_),
    .S(net89),
    .X(_1872_));
 sky130_fd_sc_hd__a22o_1 _4968_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(net62),
    .B1(net60),
    .B2(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__a21bo_1 _4969_ (.A1(net78),
    .A2(_1873_),
    .B1_N(_1863_),
    .X(_1874_));
 sky130_fd_sc_hd__mux2_1 _4970_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_1874_),
    .S(net66),
    .X(_1875_));
 sky130_fd_sc_hd__mux2_1 _4971_ (.A0(\z80.tv80s.i_tv80_core.I[2] ),
    .A1(_1875_),
    .S(net91),
    .X(_1876_));
 sky130_fd_sc_hd__mux2_1 _4972_ (.A0(net580),
    .A1(_1876_),
    .S(net55),
    .X(_0232_));
 sky130_fd_sc_hd__mux4_1 _4973_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .S0(net132),
    .S1(net163),
    .X(_1877_));
 sky130_fd_sc_hd__mux4_1 _4974_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .S0(net132),
    .S1(net163),
    .X(_1878_));
 sky130_fd_sc_hd__mux2_2 _4975_ (.A0(_1878_),
    .A1(_1877_),
    .S(net165),
    .X(_1879_));
 sky130_fd_sc_hd__nand2_1 _4976_ (.A(net80),
    .B(_1879_),
    .Y(_1880_));
 sky130_fd_sc_hd__a22o_1 _4977_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_1673_),
    .B1(_1879_),
    .B2(_1672_),
    .X(_1881_));
 sky130_fd_sc_hd__a21o_1 _4978_ (.A1(\z80.tv80s.i_tv80_core.SP[11] ),
    .A2(net58),
    .B1(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__mux2_1 _4979_ (.A0(\z80.tv80s.i_tv80_core.PC[11] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1883_));
 sky130_fd_sc_hd__mux2_1 _4980_ (.A0(_1879_),
    .A1(_1883_),
    .S(net98),
    .X(_1884_));
 sky130_fd_sc_hd__and3_1 _4981_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .C(_1849_),
    .X(_1885_));
 sky130_fd_sc_hd__a21oi_1 _4982_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .A2(_1849_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .Y(_1886_));
 sky130_fd_sc_hd__nor2_1 _4983_ (.A(_1885_),
    .B(_1886_),
    .Y(_1887_));
 sky130_fd_sc_hd__mux2_1 _4984_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_1887_),
    .S(_1685_),
    .X(_1888_));
 sky130_fd_sc_hd__a22o_1 _4985_ (.A1(net57),
    .A2(_1884_),
    .B1(_1888_),
    .B2(_1678_),
    .X(_1889_));
 sky130_fd_sc_hd__a211o_1 _4986_ (.A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .A2(_1669_),
    .B1(_1882_),
    .C1(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__mux2_1 _4987_ (.A0(\z80.tv80s.i_tv80_core.I[3] ),
    .A1(_1890_),
    .S(net89),
    .X(_1891_));
 sky130_fd_sc_hd__a22o_1 _4988_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2(net62),
    .B1(net60),
    .B2(_1891_),
    .X(_1892_));
 sky130_fd_sc_hd__a21bo_1 _4989_ (.A1(net78),
    .A2(_1892_),
    .B1_N(_1880_),
    .X(_1893_));
 sky130_fd_sc_hd__mux2_1 _4990_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_1893_),
    .S(net66),
    .X(_1894_));
 sky130_fd_sc_hd__mux2_1 _4991_ (.A0(\z80.tv80s.i_tv80_core.I[3] ),
    .A1(_1894_),
    .S(net91),
    .X(_1895_));
 sky130_fd_sc_hd__mux2_1 _4992_ (.A0(net606),
    .A1(_1895_),
    .S(net55),
    .X(_0233_));
 sky130_fd_sc_hd__mux4_1 _4993_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .S0(net132),
    .S1(net164),
    .X(_1896_));
 sky130_fd_sc_hd__mux4_1 _4994_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .S0(net132),
    .S1(net164),
    .X(_1897_));
 sky130_fd_sc_hd__mux2_2 _4995_ (.A0(_1897_),
    .A1(_1896_),
    .S(net165),
    .X(_1898_));
 sky130_fd_sc_hd__nand2_1 _4996_ (.A(net80),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__a22o_1 _4997_ (.A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(_1673_),
    .B1(_1898_),
    .B2(_1672_),
    .X(_1900_));
 sky130_fd_sc_hd__a21o_1 _4998_ (.A1(\z80.tv80s.i_tv80_core.SP[12] ),
    .A2(net58),
    .B1(_1900_),
    .X(_1901_));
 sky130_fd_sc_hd__mux2_1 _4999_ (.A0(\z80.tv80s.i_tv80_core.PC[12] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1902_));
 sky130_fd_sc_hd__mux2_1 _5000_ (.A0(_1898_),
    .A1(_1902_),
    .S(net98),
    .X(_1903_));
 sky130_fd_sc_hd__and2_1 _5001_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .B(_1885_),
    .X(_1904_));
 sky130_fd_sc_hd__nor2_1 _5002_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .B(_1885_),
    .Y(_1905_));
 sky130_fd_sc_hd__o21ai_1 _5003_ (.A1(_1904_),
    .A2(_1905_),
    .B1(_1685_),
    .Y(_1906_));
 sky130_fd_sc_hd__o21a_1 _5004_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_1685_),
    .B1(_1906_),
    .X(_1907_));
 sky130_fd_sc_hd__a22o_1 _5005_ (.A1(net57),
    .A2(_1903_),
    .B1(_1907_),
    .B2(_1678_),
    .X(_1908_));
 sky130_fd_sc_hd__a211o_1 _5006_ (.A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .A2(_1669_),
    .B1(_1901_),
    .C1(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__mux2_1 _5007_ (.A0(\z80.tv80s.i_tv80_core.I[4] ),
    .A1(_1909_),
    .S(net89),
    .X(_1910_));
 sky130_fd_sc_hd__a22o_1 _5008_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(net62),
    .B1(net60),
    .B2(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__a21bo_1 _5009_ (.A1(net78),
    .A2(_1911_),
    .B1_N(_1899_),
    .X(_1912_));
 sky130_fd_sc_hd__mux2_1 _5010_ (.A0(\z80.tv80s.di_reg[4] ),
    .A1(_1912_),
    .S(net66),
    .X(_1913_));
 sky130_fd_sc_hd__mux2_1 _5011_ (.A0(\z80.tv80s.i_tv80_core.I[4] ),
    .A1(_1913_),
    .S(net91),
    .X(_1914_));
 sky130_fd_sc_hd__mux2_1 _5012_ (.A0(net618),
    .A1(_1914_),
    .S(net55),
    .X(_0234_));
 sky130_fd_sc_hd__mux4_1 _5013_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .S0(net133),
    .S1(net164),
    .X(_1915_));
 sky130_fd_sc_hd__mux4_1 _5014_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .S0(net133),
    .S1(net164),
    .X(_1916_));
 sky130_fd_sc_hd__mux2_2 _5015_ (.A0(_1916_),
    .A1(_1915_),
    .S(net165),
    .X(_1917_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(net80),
    .B(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__a22o_1 _5017_ (.A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2(_1673_),
    .B1(_1917_),
    .B2(_1672_),
    .X(_1919_));
 sky130_fd_sc_hd__a21o_1 _5018_ (.A1(\z80.tv80s.i_tv80_core.SP[13] ),
    .A2(net58),
    .B1(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__mux2_1 _5019_ (.A0(\z80.tv80s.i_tv80_core.PC[13] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1921_));
 sky130_fd_sc_hd__mux2_1 _5020_ (.A0(_1917_),
    .A1(_1921_),
    .S(net98),
    .X(_1922_));
 sky130_fd_sc_hd__xor2_1 _5021_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .B(_1904_),
    .X(_1923_));
 sky130_fd_sc_hd__mux2_1 _5022_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1923_),
    .S(_1685_),
    .X(_1924_));
 sky130_fd_sc_hd__a22o_1 _5023_ (.A1(net57),
    .A2(_1922_),
    .B1(_1924_),
    .B2(_1678_),
    .X(_1925_));
 sky130_fd_sc_hd__a211o_1 _5024_ (.A1(\z80.tv80s.i_tv80_core.PC[13] ),
    .A2(_1669_),
    .B1(_1920_),
    .C1(_1925_),
    .X(_1926_));
 sky130_fd_sc_hd__mux2_1 _5025_ (.A0(\z80.tv80s.i_tv80_core.I[5] ),
    .A1(_1926_),
    .S(net89),
    .X(_1927_));
 sky130_fd_sc_hd__a22o_1 _5026_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(net62),
    .B1(net60),
    .B2(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__a21bo_1 _5027_ (.A1(net78),
    .A2(_1928_),
    .B1_N(_1918_),
    .X(_1929_));
 sky130_fd_sc_hd__mux2_1 _5028_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_1929_),
    .S(net66),
    .X(_1930_));
 sky130_fd_sc_hd__mux2_1 _5029_ (.A0(\z80.tv80s.i_tv80_core.I[5] ),
    .A1(_1930_),
    .S(net93),
    .X(_1931_));
 sky130_fd_sc_hd__mux2_1 _5030_ (.A0(net620),
    .A1(_1931_),
    .S(net55),
    .X(_0235_));
 sky130_fd_sc_hd__mux4_1 _5031_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .S0(net132),
    .S1(net163),
    .X(_1932_));
 sky130_fd_sc_hd__mux4_1 _5032_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .S0(net132),
    .S1(net163),
    .X(_1933_));
 sky130_fd_sc_hd__mux2_2 _5033_ (.A0(_1933_),
    .A1(_1932_),
    .S(net165),
    .X(_1934_));
 sky130_fd_sc_hd__nand2_1 _5034_ (.A(net80),
    .B(_1934_),
    .Y(_1935_));
 sky130_fd_sc_hd__a22o_1 _5035_ (.A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_1673_),
    .B1(_1934_),
    .B2(_1672_),
    .X(_1936_));
 sky130_fd_sc_hd__a21o_1 _5036_ (.A1(\z80.tv80s.i_tv80_core.SP[14] ),
    .A2(net58),
    .B1(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__mux2_1 _5037_ (.A0(\z80.tv80s.i_tv80_core.PC[14] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1938_));
 sky130_fd_sc_hd__mux2_1 _5038_ (.A0(_1934_),
    .A1(_1938_),
    .S(net98),
    .X(_1939_));
 sky130_fd_sc_hd__and3_1 _5039_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .B(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .C(_1904_),
    .X(_1940_));
 sky130_fd_sc_hd__a21oi_1 _5040_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(_1904_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .Y(_1941_));
 sky130_fd_sc_hd__nor2_1 _5041_ (.A(_1940_),
    .B(_1941_),
    .Y(_1942_));
 sky130_fd_sc_hd__mux2_1 _5042_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_1942_),
    .S(_1685_),
    .X(_1943_));
 sky130_fd_sc_hd__a22o_1 _5043_ (.A1(net57),
    .A2(_1939_),
    .B1(_1943_),
    .B2(_1678_),
    .X(_1944_));
 sky130_fd_sc_hd__a211o_1 _5044_ (.A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .A2(_1669_),
    .B1(_1937_),
    .C1(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__mux2_1 _5045_ (.A0(\z80.tv80s.i_tv80_core.I[6] ),
    .A1(_1945_),
    .S(net89),
    .X(_1946_));
 sky130_fd_sc_hd__a22o_1 _5046_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2(net62),
    .B1(net60),
    .B2(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__a21bo_1 _5047_ (.A1(net78),
    .A2(_1947_),
    .B1_N(_1935_),
    .X(_1948_));
 sky130_fd_sc_hd__mux2_1 _5048_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_1948_),
    .S(net66),
    .X(_1949_));
 sky130_fd_sc_hd__mux2_1 _5049_ (.A0(net622),
    .A1(_1949_),
    .S(net91),
    .X(_1950_));
 sky130_fd_sc_hd__mux2_1 _5050_ (.A0(net626),
    .A1(_1950_),
    .S(net55),
    .X(_0236_));
 sky130_fd_sc_hd__mux4_1 _5051_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .S0(net132),
    .S1(net163),
    .X(_1951_));
 sky130_fd_sc_hd__mux4_1 _5052_ (.A0(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .A2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .A3(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .S0(net133),
    .S1(net163),
    .X(_1952_));
 sky130_fd_sc_hd__mux2_2 _5053_ (.A0(_1952_),
    .A1(_1951_),
    .S(net165),
    .X(_1953_));
 sky130_fd_sc_hd__nand2_1 _5054_ (.A(net80),
    .B(_1953_),
    .Y(_1954_));
 sky130_fd_sc_hd__a22o_1 _5055_ (.A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(_1673_),
    .B1(_1953_),
    .B2(_1672_),
    .X(_1955_));
 sky130_fd_sc_hd__a21o_1 _5056_ (.A1(\z80.tv80s.i_tv80_core.SP[15] ),
    .A2(net58),
    .B1(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__mux2_1 _5057_ (.A0(\z80.tv80s.i_tv80_core.PC[15] ),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .S(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(_1957_));
 sky130_fd_sc_hd__mux2_1 _5058_ (.A0(_1953_),
    .A1(_1957_),
    .S(net98),
    .X(_1958_));
 sky130_fd_sc_hd__xor2_1 _5059_ (.A(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .B(_1940_),
    .X(_1959_));
 sky130_fd_sc_hd__mux2_1 _5060_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1959_),
    .S(_1685_),
    .X(_1960_));
 sky130_fd_sc_hd__a22o_1 _5061_ (.A1(net57),
    .A2(_1958_),
    .B1(_1960_),
    .B2(_1678_),
    .X(_1961_));
 sky130_fd_sc_hd__a211o_1 _5062_ (.A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .A2(_1669_),
    .B1(_1956_),
    .C1(_1961_),
    .X(_1962_));
 sky130_fd_sc_hd__mux2_1 _5063_ (.A0(\z80.tv80s.i_tv80_core.I[7] ),
    .A1(_1962_),
    .S(net89),
    .X(_1963_));
 sky130_fd_sc_hd__a22o_1 _5064_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .A2(net62),
    .B1(net60),
    .B2(_1963_),
    .X(_1964_));
 sky130_fd_sc_hd__a21bo_1 _5065_ (.A1(net78),
    .A2(_1964_),
    .B1_N(_1954_),
    .X(_1965_));
 sky130_fd_sc_hd__mux2_1 _5066_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_1965_),
    .S(net66),
    .X(_1966_));
 sky130_fd_sc_hd__mux2_1 _5067_ (.A0(\z80.tv80s.i_tv80_core.I[7] ),
    .A1(_1966_),
    .S(net91),
    .X(_1967_));
 sky130_fd_sc_hd__mux2_1 _5068_ (.A0(net664),
    .A1(_1967_),
    .S(net55),
    .X(_0237_));
 sky130_fd_sc_hd__or3b_1 _5069_ (.A(_2854_),
    .B(_2856_),
    .C_N(_0788_),
    .X(_1968_));
 sky130_fd_sc_hd__or4b_4 _5070_ (.A(net525),
    .B(_2855_),
    .C(_1968_),
    .D_N(net511),
    .X(_1969_));
 sky130_fd_sc_hd__inv_2 _5071_ (.A(_1969_),
    .Y(_1970_));
 sky130_fd_sc_hd__nor2_1 _5072_ (.A(_0863_),
    .B(_1969_),
    .Y(_1971_));
 sky130_fd_sc_hd__a21oi_4 _5073_ (.A1(net840),
    .A2(_0721_),
    .B1(_0850_),
    .Y(_1972_));
 sky130_fd_sc_hd__a21o_2 _5074_ (.A1(net896),
    .A2(_0721_),
    .B1(_0850_),
    .X(_1973_));
 sky130_fd_sc_hd__or2_1 _5075_ (.A(net56),
    .B(_1483_),
    .X(_1974_));
 sky130_fd_sc_hd__inv_2 _5076_ (.A(_1974_),
    .Y(_1975_));
 sky130_fd_sc_hd__nand2_4 _5077_ (.A(net162),
    .B(_0700_),
    .Y(_1976_));
 sky130_fd_sc_hd__a21oi_1 _5078_ (.A1(net150),
    .A2(net138),
    .B1(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__a211o_1 _5079_ (.A1(net138),
    .A2(_1976_),
    .B1(_1977_),
    .C1(_1974_),
    .X(_1978_));
 sky130_fd_sc_hd__o21ai_1 _5080_ (.A1(net707),
    .A2(_1484_),
    .B1(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__or2_2 _5081_ (.A(_0574_),
    .B(net97),
    .X(_1980_));
 sky130_fd_sc_hd__and2_1 _5082_ (.A(_1487_),
    .B(_1980_),
    .X(_1981_));
 sky130_fd_sc_hd__nand2_1 _5083_ (.A(_1487_),
    .B(_1980_),
    .Y(_1982_));
 sky130_fd_sc_hd__a2bb2o_1 _5084_ (.A1_N(net138),
    .A2_N(_1982_),
    .B1(_1979_),
    .B2(net92),
    .X(_1983_));
 sky130_fd_sc_hd__o21ai_1 _5085_ (.A1(net521),
    .A2(_1972_),
    .B1(_1983_),
    .Y(_1984_));
 sky130_fd_sc_hd__a21bo_1 _5086_ (.A1(net157),
    .A2(_1248_),
    .B1_N(_1252_),
    .X(_1985_));
 sky130_fd_sc_hd__nor2_1 _5087_ (.A(_2838_),
    .B(_0825_),
    .Y(_1986_));
 sky130_fd_sc_hd__nor2_1 _5088_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .B(net136),
    .Y(_1987_));
 sky130_fd_sc_hd__mux2_1 _5089_ (.A0(_1986_),
    .A1(_1987_),
    .S(_1985_),
    .X(_1988_));
 sky130_fd_sc_hd__o211a_1 _5090_ (.A1(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .A2(net136),
    .B1(\z80.tv80s.i_tv80_core.F[0] ),
    .C1(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_1989_));
 sky130_fd_sc_hd__a21o_1 _5091_ (.A1(net114),
    .A2(net157),
    .B1(_1272_),
    .X(_1990_));
 sky130_fd_sc_hd__a2111o_1 _5092_ (.A1(_0846_),
    .A2(_1990_),
    .B1(_1972_),
    .C1(net521),
    .D1(_1989_),
    .X(_1991_));
 sky130_fd_sc_hd__a221o_1 _5093_ (.A1(_0854_),
    .A2(_1161_),
    .B1(_1988_),
    .B2(_2836_),
    .C1(_1991_),
    .X(_1992_));
 sky130_fd_sc_hd__a31o_1 _5094_ (.A1(_1969_),
    .A2(_1984_),
    .A3(_1992_),
    .B1(_1971_),
    .X(_1993_));
 sky130_fd_sc_hd__mux2_1 _5095_ (.A0(net138),
    .A1(_1993_),
    .S(net108),
    .X(_0238_));
 sky130_fd_sc_hd__and4_2 _5096_ (.A(net124),
    .B(net99),
    .C(_0575_),
    .D(_1310_),
    .X(_1994_));
 sky130_fd_sc_hd__nor3_2 _5097_ (.A(_2832_),
    .B(_3002_),
    .C(_0677_),
    .Y(_1995_));
 sky130_fd_sc_hd__nor3_1 _5098_ (.A(_1970_),
    .B(_1994_),
    .C(_1995_),
    .Y(_1996_));
 sky130_fd_sc_hd__o221a_1 _5099_ (.A1(_2836_),
    .A2(\z80.tv80s.i_tv80_core.F[1] ),
    .B1(_0854_),
    .B2(_1986_),
    .C1(_1973_),
    .X(_1997_));
 sky130_fd_sc_hd__a21boi_1 _5100_ (.A1(_2849_),
    .A2(_1602_),
    .B1_N(_1976_),
    .Y(_1998_));
 sky130_fd_sc_hd__o22a_1 _5101_ (.A1(\z80.tv80s.i_tv80_core.Fp[1] ),
    .A2(_1484_),
    .B1(_1974_),
    .B2(_1998_),
    .X(_1999_));
 sky130_fd_sc_hd__nor2_1 _5102_ (.A(_1607_),
    .B(_1973_),
    .Y(_2000_));
 sky130_fd_sc_hd__o22a_1 _5103_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1982_),
    .B1(_1999_),
    .B2(net97),
    .X(_2001_));
 sky130_fd_sc_hd__a21o_1 _5104_ (.A1(_2000_),
    .A2(_2001_),
    .B1(_1997_),
    .X(_2002_));
 sky130_fd_sc_hd__a22o_1 _5105_ (.A1(_1004_),
    .A2(_1970_),
    .B1(_1996_),
    .B2(_2002_),
    .X(_2003_));
 sky130_fd_sc_hd__mux2_1 _5106_ (.A0(net886),
    .A1(_2003_),
    .S(net108),
    .X(_0239_));
 sky130_fd_sc_hd__or3b_1 _5107_ (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .B(_1250_),
    .C_N(_1248_),
    .X(_2004_));
 sky130_fd_sc_hd__o21ai_1 _5108_ (.A1(_1248_),
    .A2(_1252_),
    .B1(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__xnor2_1 _5109_ (.A(_1215_),
    .B(_1258_),
    .Y(_2006_));
 sky130_fd_sc_hd__xor2_1 _5110_ (.A(_1131_),
    .B(_1156_),
    .X(_2007_));
 sky130_fd_sc_hd__xor2_1 _5111_ (.A(_0840_),
    .B(_0987_),
    .X(_2008_));
 sky130_fd_sc_hd__xnor2_1 _5112_ (.A(_1039_),
    .B(_1069_),
    .Y(_2009_));
 sky130_fd_sc_hd__xnor2_1 _5113_ (.A(_2008_),
    .B(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__xnor2_1 _5114_ (.A(_2007_),
    .B(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__nor2_1 _5115_ (.A(_2006_),
    .B(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__a21o_1 _5116_ (.A1(_2006_),
    .A2(_2011_),
    .B1(_0836_),
    .X(_2013_));
 sky130_fd_sc_hd__o22a_1 _5117_ (.A1(_0835_),
    .A2(_2005_),
    .B1(_2012_),
    .B2(_2013_),
    .X(_2014_));
 sky130_fd_sc_hd__mux2_1 _5118_ (.A0(\z80.tv80s.i_tv80_core.F[2] ),
    .A1(_2014_),
    .S(_2851_),
    .X(_2015_));
 sky130_fd_sc_hd__xnor2_1 _5119_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_0998_),
    .Y(_2016_));
 sky130_fd_sc_hd__xor2_1 _5120_ (.A(_1223_),
    .B(_1270_),
    .X(_2017_));
 sky130_fd_sc_hd__xnor2_1 _5121_ (.A(_2016_),
    .B(_2017_),
    .Y(_2018_));
 sky130_fd_sc_hd__xnor2_1 _5122_ (.A(_1117_),
    .B(_1168_),
    .Y(_2019_));
 sky130_fd_sc_hd__xnor2_1 _5123_ (.A(_1042_),
    .B(_1075_),
    .Y(_2020_));
 sky130_fd_sc_hd__xnor2_1 _5124_ (.A(_2019_),
    .B(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__xnor2_1 _5125_ (.A(_2018_),
    .B(_2021_),
    .Y(_2022_));
 sky130_fd_sc_hd__nor2_1 _5126_ (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .B(_1159_),
    .Y(_2023_));
 sky130_fd_sc_hd__a211o_1 _5127_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_1267_),
    .B1(_2023_),
    .C1(_1160_),
    .X(_2024_));
 sky130_fd_sc_hd__xnor2_1 _5128_ (.A(_2022_),
    .B(_2024_),
    .Y(_2025_));
 sky130_fd_sc_hd__xor2_1 _5129_ (.A(_1225_),
    .B(_1274_),
    .X(_2026_));
 sky130_fd_sc_hd__xor2_1 _5130_ (.A(_0849_),
    .B(_0989_),
    .X(_2027_));
 sky130_fd_sc_hd__xor2_1 _5131_ (.A(_1044_),
    .B(_1077_),
    .X(_2028_));
 sky130_fd_sc_hd__xor2_1 _5132_ (.A(_1119_),
    .B(_1171_),
    .X(_2029_));
 sky130_fd_sc_hd__xnor2_1 _5133_ (.A(_2028_),
    .B(_2029_),
    .Y(_2030_));
 sky130_fd_sc_hd__xnor2_1 _5134_ (.A(_2027_),
    .B(_2030_),
    .Y(_2031_));
 sky130_fd_sc_hd__nor2_1 _5135_ (.A(_2026_),
    .B(_2031_),
    .Y(_2032_));
 sky130_fd_sc_hd__a21o_1 _5136_ (.A1(_2026_),
    .A2(_2031_),
    .B1(net162),
    .X(_2033_));
 sky130_fd_sc_hd__o22a_1 _5137_ (.A1(net111),
    .A2(\z80.tv80s.i_tv80_core.F[2] ),
    .B1(_2032_),
    .B2(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__xor2_1 _5138_ (.A(_1043_),
    .B(_1076_),
    .X(_2035_));
 sky130_fd_sc_hd__xor2_1 _5139_ (.A(_0858_),
    .B(_0988_),
    .X(_2036_));
 sky130_fd_sc_hd__xnor2_1 _5140_ (.A(_2035_),
    .B(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__xor2_1 _5141_ (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .B(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(_2038_));
 sky130_fd_sc_hd__xnor2_1 _5142_ (.A(_1259_),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__xnor2_1 _5143_ (.A(_2037_),
    .B(_2039_),
    .Y(_2040_));
 sky130_fd_sc_hd__a22o_1 _5144_ (.A1(\z80.tv80s.i_tv80_core.BusB[1] ),
    .A2(_0464_),
    .B1(_1046_),
    .B2(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(_2041_));
 sky130_fd_sc_hd__a22o_1 _5145_ (.A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A2(_0459_),
    .B1(_0465_),
    .B2(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(_2042_));
 sky130_fd_sc_hd__a221o_1 _5146_ (.A1(\z80.tv80s.i_tv80_core.BusB[6] ),
    .A2(_2881_),
    .B1(_0455_),
    .B2(\z80.tv80s.i_tv80_core.BusB[3] ),
    .C1(_2042_),
    .X(_2043_));
 sky130_fd_sc_hd__a211o_1 _5147_ (.A1(\z80.tv80s.i_tv80_core.BusB[7] ),
    .A2(_0467_),
    .B1(_0851_),
    .C1(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__a211o_1 _5148_ (.A1(\z80.tv80s.i_tv80_core.BusB[4] ),
    .A2(_0460_),
    .B1(_2041_),
    .C1(_2044_),
    .X(_2045_));
 sky130_fd_sc_hd__and2_1 _5149_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_1986_),
    .X(_2046_));
 sky130_fd_sc_hd__nand2_1 _5150_ (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .B(_1986_),
    .Y(_2047_));
 sky130_fd_sc_hd__a22o_1 _5151_ (.A1(_0846_),
    .A2(_2034_),
    .B1(_2040_),
    .B2(_0856_),
    .X(_2048_));
 sky130_fd_sc_hd__a221o_1 _5152_ (.A1(_0854_),
    .A2(_2025_),
    .B1(_2046_),
    .B2(\z80.tv80s.i_tv80_core.F[2] ),
    .C1(_1972_),
    .X(_2049_));
 sky130_fd_sc_hd__a21o_1 _5153_ (.A1(_2836_),
    .A2(_2015_),
    .B1(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__or3b_1 _5154_ (.A(_2048_),
    .B(_2050_),
    .C_N(_2045_),
    .X(_2051_));
 sky130_fd_sc_hd__mux2_1 _5155_ (.A0(\z80.tv80s.i_tv80_core.Fp[2] ),
    .A1(\z80.tv80s.i_tv80_core.F[2] ),
    .S(_1487_),
    .X(_2052_));
 sky130_fd_sc_hd__mux2_1 _5156_ (.A0(net805),
    .A1(_2052_),
    .S(_1608_),
    .X(_2053_));
 sky130_fd_sc_hd__o21ba_1 _5157_ (.A1(_1973_),
    .A2(_2053_),
    .B1_N(_1994_),
    .X(_2054_));
 sky130_fd_sc_hd__nor2_1 _5158_ (.A(_3004_),
    .B(_0677_),
    .Y(_2055_));
 sky130_fd_sc_hd__xor2_1 _5159_ (.A(\z80.tv80s.di_reg[5] ),
    .B(\z80.tv80s.di_reg[4] ),
    .X(_2056_));
 sky130_fd_sc_hd__xor2_1 _5160_ (.A(\z80.tv80s.di_reg[1] ),
    .B(\z80.tv80s.di_reg[0] ),
    .X(_2057_));
 sky130_fd_sc_hd__xor2_1 _5161_ (.A(\z80.tv80s.di_reg[7] ),
    .B(\z80.tv80s.di_reg[6] ),
    .X(_2058_));
 sky130_fd_sc_hd__xor2_1 _5162_ (.A(\z80.tv80s.di_reg[3] ),
    .B(\z80.tv80s.di_reg[2] ),
    .X(_2059_));
 sky130_fd_sc_hd__xnor2_1 _5163_ (.A(_2058_),
    .B(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__xnor2_1 _5164_ (.A(_2057_),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__xnor2_1 _5165_ (.A(_2056_),
    .B(_2061_),
    .Y(_2062_));
 sky130_fd_sc_hd__a221o_1 _5166_ (.A1(_2051_),
    .A2(_2054_),
    .B1(_2062_),
    .B2(_1994_),
    .C1(_2055_),
    .X(_2063_));
 sky130_fd_sc_hd__o311a_1 _5167_ (.A1(net574),
    .A2(_3004_),
    .A3(_0677_),
    .B1(_1969_),
    .C1(_2063_),
    .X(_2064_));
 sky130_fd_sc_hd__o21ai_1 _5168_ (.A1(_1053_),
    .A2(_1969_),
    .B1(net108),
    .Y(_2065_));
 sky130_fd_sc_hd__o22a_1 _5169_ (.A1(net827),
    .A2(net108),
    .B1(_2064_),
    .B2(_2065_),
    .X(_0240_));
 sky130_fd_sc_hd__mux2_1 _5170_ (.A0(_2859_),
    .A1(\z80.tv80s.i_tv80_core.F[3] ),
    .S(_1602_),
    .X(_2066_));
 sky130_fd_sc_hd__mux2_1 _5171_ (.A0(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A1(_2066_),
    .S(_1976_),
    .X(_2067_));
 sky130_fd_sc_hd__a22o_1 _5172_ (.A1(\z80.tv80s.i_tv80_core.Fp[3] ),
    .A2(_1483_),
    .B1(_1975_),
    .B2(_2067_),
    .X(_2068_));
 sky130_fd_sc_hd__a221o_1 _5173_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_1981_),
    .B1(_2068_),
    .B2(net92),
    .C1(_1973_),
    .X(_2069_));
 sky130_fd_sc_hd__mux2_1 _5174_ (.A0(net656),
    .A1(_1069_),
    .S(_0785_),
    .X(_2070_));
 sky130_fd_sc_hd__a31o_1 _5175_ (.A1(\z80.tv80s.i_tv80_core.BusB[3] ),
    .A2(_2885_),
    .A3(_0850_),
    .B1(_1078_),
    .X(_2071_));
 sky130_fd_sc_hd__a2111o_1 _5176_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_2046_),
    .B1(_2071_),
    .C1(_1079_),
    .D1(_1972_),
    .X(_2072_));
 sky130_fd_sc_hd__a21oi_1 _5177_ (.A1(_2836_),
    .A2(_2070_),
    .B1(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__nor2_1 _5178_ (.A(_1995_),
    .B(_2073_),
    .Y(_2074_));
 sky130_fd_sc_hd__a22o_1 _5179_ (.A1(_1083_),
    .A2(_1995_),
    .B1(_2069_),
    .B2(_2074_),
    .X(_2075_));
 sky130_fd_sc_hd__mux2_1 _5180_ (.A0(_1087_),
    .A1(_2075_),
    .S(_1969_),
    .X(_2076_));
 sky130_fd_sc_hd__mux2_1 _5181_ (.A0(net816),
    .A1(_2076_),
    .S(net108),
    .X(_0241_));
 sky130_fd_sc_hd__nand2_1 _5182_ (.A(_1125_),
    .B(_1987_),
    .Y(_2077_));
 sky130_fd_sc_hd__o311a_1 _5183_ (.A1(_2838_),
    .A2(_0825_),
    .A3(_1125_),
    .B1(_2077_),
    .C1(_0853_),
    .X(_2078_));
 sky130_fd_sc_hd__o22a_1 _5184_ (.A1(_0855_),
    .A2(_1116_),
    .B1(_2078_),
    .B2(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_2079_));
 sky130_fd_sc_hd__o211ai_1 _5185_ (.A1(_2850_),
    .A2(_2047_),
    .B1(_2079_),
    .C1(_0851_),
    .Y(_2080_));
 sky130_fd_sc_hd__o311a_1 _5186_ (.A1(net114),
    .A2(_1976_),
    .A3(_1980_),
    .B1(_2850_),
    .C1(_1604_),
    .X(_2081_));
 sky130_fd_sc_hd__a2bb2o_1 _5187_ (.A1_N(\z80.tv80s.i_tv80_core.Fp[4] ),
    .A2_N(_1484_),
    .B1(_1975_),
    .B2(_1977_),
    .X(_2082_));
 sky130_fd_sc_hd__a21bo_1 _5188_ (.A1(net92),
    .A2(_2082_),
    .B1_N(_2000_),
    .X(_2083_));
 sky130_fd_sc_hd__a2bb2o_1 _5189_ (.A1_N(_2081_),
    .A2_N(_2083_),
    .B1(_1973_),
    .B2(_2080_),
    .X(_2084_));
 sky130_fd_sc_hd__a22o_1 _5190_ (.A1(_1141_),
    .A2(_1970_),
    .B1(_1996_),
    .B2(_2084_),
    .X(_2085_));
 sky130_fd_sc_hd__mux2_1 _5191_ (.A0(net830),
    .A1(_2085_),
    .S(net109),
    .X(_0242_));
 sky130_fd_sc_hd__mux2_1 _5192_ (.A0(_2860_),
    .A1(\z80.tv80s.i_tv80_core.F[5] ),
    .S(_1602_),
    .X(_2086_));
 sky130_fd_sc_hd__mux2_1 _5193_ (.A0(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A1(_2086_),
    .S(_1976_),
    .X(_2087_));
 sky130_fd_sc_hd__a22o_1 _5194_ (.A1(\z80.tv80s.i_tv80_core.Fp[5] ),
    .A2(_1483_),
    .B1(_1975_),
    .B2(_2087_),
    .X(_2088_));
 sky130_fd_sc_hd__a221o_1 _5195_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_1981_),
    .B1(_2088_),
    .B2(net92),
    .C1(_1973_),
    .X(_2089_));
 sky130_fd_sc_hd__mux2_1 _5196_ (.A0(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A1(_1156_),
    .S(_0785_),
    .X(_2090_));
 sky130_fd_sc_hd__a31o_1 _5197_ (.A1(\z80.tv80s.i_tv80_core.BusB[5] ),
    .A2(_2885_),
    .A3(_0850_),
    .B1(_1170_),
    .X(_2091_));
 sky130_fd_sc_hd__a221o_1 _5198_ (.A1(_0846_),
    .A2(_1171_),
    .B1(_2046_),
    .B2(\z80.tv80s.i_tv80_core.F[5] ),
    .C1(_2091_),
    .X(_2092_));
 sky130_fd_sc_hd__a21oi_1 _5199_ (.A1(_2836_),
    .A2(_2090_),
    .B1(_2092_),
    .Y(_2093_));
 sky130_fd_sc_hd__a21oi_1 _5200_ (.A1(_1973_),
    .A2(_2093_),
    .B1(_1995_),
    .Y(_2094_));
 sky130_fd_sc_hd__a22o_1 _5201_ (.A1(_1000_),
    .A2(_1995_),
    .B1(_2089_),
    .B2(_2094_),
    .X(_2095_));
 sky130_fd_sc_hd__mux2_1 _5202_ (.A0(_1178_),
    .A1(_2095_),
    .S(_1969_),
    .X(_2096_));
 sky130_fd_sc_hd__mux2_1 _5203_ (.A0(net817),
    .A1(_2096_),
    .S(net109),
    .X(_0243_));
 sky130_fd_sc_hd__a211o_1 _5204_ (.A1(_2828_),
    .A2(\z80.tv80s.i_tv80_core.Z16_r ),
    .B1(_0840_),
    .C1(_0987_),
    .X(_2097_));
 sky130_fd_sc_hd__or3b_1 _5205_ (.A(_2097_),
    .B(_1069_),
    .C_N(_1039_),
    .X(_2098_));
 sky130_fd_sc_hd__or3b_1 _5206_ (.A(_2098_),
    .B(_1156_),
    .C_N(_1131_),
    .X(_2099_));
 sky130_fd_sc_hd__o31a_1 _5207_ (.A1(_1215_),
    .A2(_1258_),
    .A3(_2099_),
    .B1(_2851_),
    .X(_2100_));
 sky130_fd_sc_hd__a211o_1 _5208_ (.A1(_2828_),
    .A2(\z80.tv80s.i_tv80_core.Arith16_r ),
    .B1(_2100_),
    .C1(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(_2101_));
 sky130_fd_sc_hd__or3b_1 _5209_ (.A(_0855_),
    .B(_1042_),
    .C_N(_1075_),
    .X(_2102_));
 sky130_fd_sc_hd__or3_1 _5210_ (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .B(_0999_),
    .C(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__or4_1 _5211_ (.A(_1044_),
    .B(_1077_),
    .C(_1119_),
    .D(_1171_),
    .X(_2104_));
 sky130_fd_sc_hd__or3_1 _5212_ (.A(_1225_),
    .B(_1274_),
    .C(_2104_),
    .X(_2105_));
 sky130_fd_sc_hd__o31a_1 _5213_ (.A1(_0849_),
    .A2(_0989_),
    .A3(_2105_),
    .B1(net111),
    .X(_2106_));
 sky130_fd_sc_hd__o21ai_1 _5214_ (.A1(net111),
    .A2(\z80.tv80s.i_tv80_core.F[6] ),
    .B1(_0846_),
    .Y(_2107_));
 sky130_fd_sc_hd__or2_1 _5215_ (.A(_2106_),
    .B(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__or4_1 _5216_ (.A(_0858_),
    .B(_0988_),
    .C(_1043_),
    .D(_1076_),
    .X(_2109_));
 sky130_fd_sc_hd__or4_1 _5217_ (.A(net157),
    .B(\z80.tv80s.i_tv80_core.BusA[4] ),
    .C(\z80.tv80s.i_tv80_core.BusA[5] ),
    .D(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(_2110_));
 sky130_fd_sc_hd__o311a_1 _5218_ (.A1(_0857_),
    .A2(_2109_),
    .A3(_2110_),
    .B1(_2045_),
    .C1(_2047_),
    .X(_2111_));
 sky130_fd_sc_hd__or4_1 _5219_ (.A(_1118_),
    .B(_1168_),
    .C(_1270_),
    .D(_2103_),
    .X(_2112_));
 sky130_fd_sc_hd__o211a_1 _5220_ (.A1(_1223_),
    .A2(_2112_),
    .B1(_2111_),
    .C1(_2108_),
    .X(_2113_));
 sky130_fd_sc_hd__o2bb2a_2 _5221_ (.A1_N(_2113_),
    .A2_N(_2101_),
    .B1(_2047_),
    .B2(\z80.tv80s.i_tv80_core.F[6] ),
    .X(_2114_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(\z80.tv80s.i_tv80_core.Fp[6] ),
    .A1(\z80.tv80s.i_tv80_core.F[6] ),
    .S(_1487_),
    .X(_2115_));
 sky130_fd_sc_hd__or4_1 _5223_ (.A(\z80.tv80s.i_tv80_core.I[5] ),
    .B(\z80.tv80s.i_tv80_core.I[4] ),
    .C(\z80.tv80s.i_tv80_core.I[7] ),
    .D(\z80.tv80s.i_tv80_core.I[6] ),
    .X(_2116_));
 sky130_fd_sc_hd__or4_1 _5224_ (.A(\z80.tv80s.i_tv80_core.I[1] ),
    .B(\z80.tv80s.i_tv80_core.I[0] ),
    .C(\z80.tv80s.i_tv80_core.I[3] ),
    .D(\z80.tv80s.i_tv80_core.I[2] ),
    .X(_2117_));
 sky130_fd_sc_hd__nor2_1 _5225_ (.A(_2116_),
    .B(_2117_),
    .Y(_2118_));
 sky130_fd_sc_hd__and4_1 _5226_ (.A(net144),
    .B(\z80.tv80s.i_tv80_core.ts[3] ),
    .C(_1369_),
    .D(_2118_),
    .X(_2119_));
 sky130_fd_sc_hd__a21o_1 _5227_ (.A1(_1608_),
    .A2(_2115_),
    .B1(_2119_),
    .X(_2120_));
 sky130_fd_sc_hd__mux2_1 _5228_ (.A0(_2114_),
    .A1(_2120_),
    .S(_1972_),
    .X(_2121_));
 sky130_fd_sc_hd__or4_1 _5229_ (.A(\z80.tv80s.di_reg[1] ),
    .B(\z80.tv80s.di_reg[0] ),
    .C(\z80.tv80s.di_reg[5] ),
    .D(\z80.tv80s.di_reg[4] ),
    .X(_2122_));
 sky130_fd_sc_hd__or4_1 _5230_ (.A(\z80.tv80s.di_reg[3] ),
    .B(\z80.tv80s.di_reg[2] ),
    .C(\z80.tv80s.di_reg[7] ),
    .D(\z80.tv80s.di_reg[6] ),
    .X(_2123_));
 sky130_fd_sc_hd__o21ai_1 _5231_ (.A1(_2122_),
    .A2(_2123_),
    .B1(_1994_),
    .Y(_2124_));
 sky130_fd_sc_hd__o21a_1 _5232_ (.A1(_1994_),
    .A2(_2121_),
    .B1(_2124_),
    .X(_2125_));
 sky130_fd_sc_hd__mux2_1 _5233_ (.A0(_1233_),
    .A1(_2125_),
    .S(_1969_),
    .X(_2126_));
 sky130_fd_sc_hd__mux2_1 _5234_ (.A0(net869),
    .A1(_2126_),
    .S(net108),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5235_ (.A0(\z80.tv80s.i_tv80_core.F[7] ),
    .A1(_1258_),
    .S(_2851_),
    .X(_2127_));
 sky130_fd_sc_hd__mux2_1 _5236_ (.A0(\z80.tv80s.i_tv80_core.F[7] ),
    .A1(_1274_),
    .S(net112),
    .X(_2128_));
 sky130_fd_sc_hd__a22o_1 _5237_ (.A1(_2836_),
    .A2(_2127_),
    .B1(_2128_),
    .B2(_0846_),
    .X(_2129_));
 sky130_fd_sc_hd__a2111o_1 _5238_ (.A1(\z80.tv80s.i_tv80_core.F[7] ),
    .A2(_2046_),
    .B1(_2129_),
    .C1(_1271_),
    .D1(_1277_),
    .X(_2130_));
 sky130_fd_sc_hd__mux2_1 _5239_ (.A0(\z80.tv80s.i_tv80_core.Fp[7] ),
    .A1(\z80.tv80s.i_tv80_core.F[7] ),
    .S(_1487_),
    .X(_2131_));
 sky130_fd_sc_hd__mux2_1 _5240_ (.A0(net777),
    .A1(_2131_),
    .S(_1608_),
    .X(_2132_));
 sky130_fd_sc_hd__mux2_1 _5241_ (.A0(_2130_),
    .A1(_2132_),
    .S(_1972_),
    .X(_2133_));
 sky130_fd_sc_hd__mux2_1 _5242_ (.A0(_2133_),
    .A1(\z80.tv80s.di_reg[7] ),
    .S(_1994_),
    .X(_2134_));
 sky130_fd_sc_hd__mux2_1 _5243_ (.A0(_1282_),
    .A1(_2134_),
    .S(_1969_),
    .X(_2135_));
 sky130_fd_sc_hd__mux2_1 _5244_ (.A0(net834),
    .A1(_2135_),
    .S(net109),
    .X(_0245_));
 sky130_fd_sc_hd__o2111ai_4 _5245_ (.A1(net117),
    .A2(_0793_),
    .B1(_0776_),
    .C1(_0769_),
    .D1(_0766_),
    .Y(_2136_));
 sky130_fd_sc_hd__inv_2 _5246_ (.A(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__or2_1 _5247_ (.A(_2835_),
    .B(_0721_),
    .X(_2138_));
 sky130_fd_sc_hd__a21oi_1 _5248_ (.A1(_2136_),
    .A2(_2138_),
    .B1(net122),
    .Y(_2139_));
 sky130_fd_sc_hd__or4_1 _5249_ (.A(_0951_),
    .B(_0960_),
    .C(_0962_),
    .D(_2136_),
    .X(_2140_));
 sky130_fd_sc_hd__or4b_1 _5250_ (.A(_0974_),
    .B(_1449_),
    .C(_2140_),
    .D_N(_1444_),
    .X(_2141_));
 sky130_fd_sc_hd__or4b_1 _5251_ (.A(_1014_),
    .B(_1462_),
    .C(_2141_),
    .D_N(_1455_),
    .X(_2142_));
 sky130_fd_sc_hd__or3b_1 _5252_ (.A(_2142_),
    .B(_1029_),
    .C_N(_1468_),
    .X(_2143_));
 sky130_fd_sc_hd__or4b_1 _5253_ (.A(_1096_),
    .B(_1189_),
    .C(_2143_),
    .D_N(_1114_),
    .X(_2144_));
 sky130_fd_sc_hd__o32a_1 _5254_ (.A1(_1205_),
    .A2(_1246_),
    .A3(_2144_),
    .B1(_2137_),
    .B2(_2114_),
    .X(_2145_));
 sky130_fd_sc_hd__mux2_1 _5255_ (.A0(net574),
    .A1(_2145_),
    .S(_2139_),
    .X(_0246_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(net102),
    .B(_0530_),
    .Y(_2146_));
 sky130_fd_sc_hd__o221a_1 _5257_ (.A1(net146),
    .A2(_0530_),
    .B1(_2146_),
    .B2(_2931_),
    .C1(net88),
    .X(_2147_));
 sky130_fd_sc_hd__nor2_1 _5258_ (.A(net129),
    .B(net88),
    .Y(_2148_));
 sky130_fd_sc_hd__a21oi_1 _5259_ (.A1(_2897_),
    .A2(_2930_),
    .B1(_2934_),
    .Y(_2149_));
 sky130_fd_sc_hd__nor3_1 _5260_ (.A(_3010_),
    .B(_3018_),
    .C(_2149_),
    .Y(_2150_));
 sky130_fd_sc_hd__o21ai_1 _5261_ (.A1(net88),
    .A2(net102),
    .B1(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__o22a_1 _5262_ (.A1(net146),
    .A2(net129),
    .B1(_2148_),
    .B2(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__o21a_1 _5263_ (.A1(_2147_),
    .A2(_2152_),
    .B1(\z80.tv80s.i_tv80_core.ISet[2] ),
    .X(_2153_));
 sky130_fd_sc_hd__nor2_1 _5264_ (.A(_2942_),
    .B(_0536_),
    .Y(_2154_));
 sky130_fd_sc_hd__nor2_1 _5265_ (.A(net127),
    .B(_3007_),
    .Y(_2155_));
 sky130_fd_sc_hd__or4_1 _5266_ (.A(_2945_),
    .B(_0485_),
    .C(_2154_),
    .D(_2155_),
    .X(_2156_));
 sky130_fd_sc_hd__a211o_1 _5267_ (.A1(_2944_),
    .A2(_0392_),
    .B1(_1407_),
    .C1(net147),
    .X(_2157_));
 sky130_fd_sc_hd__a221o_1 _5268_ (.A1(net147),
    .A2(_2944_),
    .B1(_2156_),
    .B2(_2157_),
    .C1(_0684_),
    .X(_2158_));
 sky130_fd_sc_hd__a211o_1 _5269_ (.A1(_2980_),
    .A2(_2992_),
    .B1(_0408_),
    .C1(_0501_),
    .X(_2159_));
 sky130_fd_sc_hd__or3_1 _5270_ (.A(net87),
    .B(_2975_),
    .C(_2988_),
    .X(_2160_));
 sky130_fd_sc_hd__or4b_1 _5271_ (.A(_2982_),
    .B(_2983_),
    .C(_0411_),
    .D_N(_0419_),
    .X(_2161_));
 sky130_fd_sc_hd__or4_1 _5272_ (.A(_0508_),
    .B(_0709_),
    .C(_1680_),
    .D(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__or4_2 _5273_ (.A(_3022_),
    .B(_2159_),
    .C(_2160_),
    .D(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__a22o_1 _5274_ (.A1(_2825_),
    .A2(_0511_),
    .B1(_2163_),
    .B2(net146),
    .X(_2164_));
 sky130_fd_sc_hd__a221o_1 _5275_ (.A1(net99),
    .A2(_2158_),
    .B1(_2164_),
    .B2(net160),
    .C1(_2153_),
    .X(_2165_));
 sky130_fd_sc_hd__a221o_1 _5276_ (.A1(_2879_),
    .A2(_0484_),
    .B1(_0511_),
    .B2(_0391_),
    .C1(_2163_),
    .X(_2166_));
 sky130_fd_sc_hd__a21oi_1 _5277_ (.A1(net130),
    .A2(_2885_),
    .B1(_0531_),
    .Y(_2167_));
 sky130_fd_sc_hd__a211o_1 _5278_ (.A1(_2944_),
    .A2(_0391_),
    .B1(_2154_),
    .C1(_2155_),
    .X(_2168_));
 sky130_fd_sc_hd__a32o_1 _5279_ (.A1(net114),
    .A2(_2823_),
    .A3(_2980_),
    .B1(_2166_),
    .B2(net140),
    .X(_2169_));
 sky130_fd_sc_hd__a21o_1 _5280_ (.A1(net139),
    .A2(_2168_),
    .B1(_0486_),
    .X(_2170_));
 sky130_fd_sc_hd__a32o_1 _5281_ (.A1(net139),
    .A2(\z80.tv80s.i_tv80_core.ISet[2] ),
    .A3(_2167_),
    .B1(_2170_),
    .B2(net100),
    .X(_2171_));
 sky130_fd_sc_hd__a21oi_1 _5282_ (.A1(net162),
    .A2(_2169_),
    .B1(_2171_),
    .Y(_2172_));
 sky130_fd_sc_hd__inv_2 _5283_ (.A(_2172_),
    .Y(_2173_));
 sky130_fd_sc_hd__and3_1 _5284_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .B(\z80.tv80s.i_tv80_core.ISet[1] ),
    .C(net109),
    .X(_2174_));
 sky130_fd_sc_hd__a32o_1 _5285_ (.A1(_2165_),
    .A2(_2172_),
    .A3(_2174_),
    .B1(net330),
    .B2(net122),
    .X(_0247_));
 sky130_fd_sc_hd__nor2_2 _5286_ (.A(net121),
    .B(_1980_),
    .Y(_2175_));
 sky130_fd_sc_hd__a22o_1 _5287_ (.A1(net121),
    .A2(net852),
    .B1(_2165_),
    .B2(_2175_),
    .X(_0248_));
 sky130_fd_sc_hd__o21ai_1 _5288_ (.A1(\z80.tv80s.i_tv80_core.IR[5] ),
    .A2(_2926_),
    .B1(_2898_),
    .Y(_2176_));
 sky130_fd_sc_hd__o21bai_1 _5289_ (.A1(_2914_),
    .A2(_2917_),
    .B1_N(_3027_),
    .Y(_2177_));
 sky130_fd_sc_hd__a311o_1 _5290_ (.A1(_2868_),
    .A2(_2949_),
    .A3(_2176_),
    .B1(_2177_),
    .C1(_2973_),
    .X(_2178_));
 sky130_fd_sc_hd__or3b_1 _5291_ (.A(_2977_),
    .B(_0403_),
    .C_N(_0419_),
    .X(_2179_));
 sky130_fd_sc_hd__or4_1 _5292_ (.A(_2984_),
    .B(_3022_),
    .C(_0560_),
    .D(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__or3_1 _5293_ (.A(_2989_),
    .B(_2178_),
    .C(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__or4_1 _5294_ (.A(_3010_),
    .B(_3018_),
    .C(_2149_),
    .D(_2181_),
    .X(_2182_));
 sky130_fd_sc_hd__a22o_1 _5295_ (.A1(net841),
    .A2(_0531_),
    .B1(_2167_),
    .B2(net142),
    .X(_2183_));
 sky130_fd_sc_hd__a21o_1 _5296_ (.A1(_0446_),
    .A2(_2182_),
    .B1(_2183_),
    .X(_2184_));
 sky130_fd_sc_hd__a31o_1 _5297_ (.A1(net147),
    .A2(_2944_),
    .A3(_0391_),
    .B1(_0485_),
    .X(_2185_));
 sky130_fd_sc_hd__o22a_1 _5298_ (.A1(net145),
    .A2(_1407_),
    .B1(_2185_),
    .B2(_0537_),
    .X(_2186_));
 sky130_fd_sc_hd__o21a_1 _5299_ (.A1(net142),
    .A2(_0392_),
    .B1(_2945_),
    .X(_2187_));
 sky130_fd_sc_hd__a221o_1 _5300_ (.A1(_3008_),
    .A2(_0446_),
    .B1(_0545_),
    .B2(net114),
    .C1(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__o31a_1 _5301_ (.A1(_2942_),
    .A2(_2186_),
    .A3(_2188_),
    .B1(net100),
    .X(_2189_));
 sky130_fd_sc_hd__a211o_1 _5302_ (.A1(_0391_),
    .A2(_0511_),
    .B1(_1296_),
    .C1(_2163_),
    .X(_2190_));
 sky130_fd_sc_hd__nor2_1 _5303_ (.A(_2887_),
    .B(_2918_),
    .Y(_2191_));
 sky130_fd_sc_hd__a211o_1 _5304_ (.A1(net145),
    .A2(_2190_),
    .B1(_2191_),
    .C1(_2923_),
    .X(_2192_));
 sky130_fd_sc_hd__a221o_1 _5305_ (.A1(net158),
    .A2(_2184_),
    .B1(_2192_),
    .B2(net160),
    .C1(_2189_),
    .X(_2193_));
 sky130_fd_sc_hd__a22o_1 _5306_ (.A1(net121),
    .A2(net137),
    .B1(_2175_),
    .B2(_2193_),
    .X(_0249_));
 sky130_fd_sc_hd__a22o_1 _5307_ (.A1(net121),
    .A2(net843),
    .B1(_2173_),
    .B2(_2175_),
    .X(_0250_));
 sky130_fd_sc_hd__and2b_1 _5308_ (.A_N(_2167_),
    .B(net158),
    .X(_2194_));
 sky130_fd_sc_hd__a211o_1 _5309_ (.A1(net162),
    .A2(_1303_),
    .B1(_2194_),
    .C1(net101),
    .X(_2195_));
 sky130_fd_sc_hd__a32o_1 _5310_ (.A1(_1309_),
    .A2(_2175_),
    .A3(_2195_),
    .B1(net833),
    .B2(net122),
    .X(_0251_));
 sky130_fd_sc_hd__o21ai_1 _5311_ (.A1(net88),
    .A2(_2940_),
    .B1(_2150_),
    .Y(_2196_));
 sky130_fd_sc_hd__a2bb2o_1 _5312_ (.A1_N(_2885_),
    .A2_N(_2146_),
    .B1(_2196_),
    .B2(net129),
    .X(_2197_));
 sky130_fd_sc_hd__and2_1 _5313_ (.A(net158),
    .B(_2197_),
    .X(_2198_));
 sky130_fd_sc_hd__or2_1 _5314_ (.A(_1304_),
    .B(_1340_),
    .X(_2199_));
 sky130_fd_sc_hd__or3_1 _5315_ (.A(_0692_),
    .B(_1301_),
    .C(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__o221a_1 _5316_ (.A1(net113),
    .A2(_3007_),
    .B1(_0385_),
    .B2(_0514_),
    .C1(_0683_),
    .X(_2201_));
 sky130_fd_sc_hd__or3b_1 _5317_ (.A(_2942_),
    .B(_1407_),
    .C_N(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__a221o_1 _5318_ (.A1(net160),
    .A2(_2200_),
    .B1(_2202_),
    .B2(net100),
    .C1(_2198_),
    .X(_2203_));
 sky130_fd_sc_hd__a22o_1 _5319_ (.A1(net121),
    .A2(net840),
    .B1(_2175_),
    .B2(_2203_),
    .X(_0252_));
 sky130_fd_sc_hd__nor2_1 _5320_ (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .B(_0678_),
    .Y(_2204_));
 sky130_fd_sc_hd__mux2_1 _5321_ (.A0(net345),
    .A1(_2204_),
    .S(_2175_),
    .X(_0253_));
 sky130_fd_sc_hd__or4_1 _5322_ (.A(_2980_),
    .B(_2983_),
    .C(_3024_),
    .D(_0411_),
    .X(_2205_));
 sky130_fd_sc_hd__or3_1 _5323_ (.A(_2964_),
    .B(_2982_),
    .C(_0415_),
    .X(_2206_));
 sky130_fd_sc_hd__or4_1 _5324_ (.A(_0425_),
    .B(_0506_),
    .C(_0662_),
    .D(_2206_),
    .X(_2207_));
 sky130_fd_sc_hd__nand2_1 _5325_ (.A(_2936_),
    .B(_0433_),
    .Y(_2208_));
 sky130_fd_sc_hd__or4_1 _5326_ (.A(_0477_),
    .B(_0505_),
    .C(_1408_),
    .D(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__or4_1 _5327_ (.A(_0710_),
    .B(_2205_),
    .C(_2207_),
    .D(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__and3_1 _5328_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .B(_2951_),
    .C(_0467_),
    .X(_2211_));
 sky130_fd_sc_hd__a31o_1 _5329_ (.A1(net147),
    .A2(_2975_),
    .A3(_0513_),
    .B1(_2211_),
    .X(_2212_));
 sky130_fd_sc_hd__mux2_1 _5330_ (.A0(net126),
    .A1(_2212_),
    .S(_2210_),
    .X(_2213_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(_2942_),
    .A2(net99),
    .B1(_2213_),
    .B2(net159),
    .X(_2214_));
 sky130_fd_sc_hd__inv_2 _5332_ (.A(_2214_),
    .Y(_2215_));
 sky130_fd_sc_hd__o21a_1 _5333_ (.A1(_1509_),
    .A2(_2214_),
    .B1(_0575_),
    .X(_2216_));
 sky130_fd_sc_hd__mux2_1 _5334_ (.A0(net630),
    .A1(_2216_),
    .S(net106),
    .X(_0254_));
 sky130_fd_sc_hd__a21oi_1 _5335_ (.A1(_1315_),
    .A2(_2215_),
    .B1(_0574_),
    .Y(_2217_));
 sky130_fd_sc_hd__mux2_1 _5336_ (.A0(net511),
    .A1(_2217_),
    .S(net106),
    .X(_0255_));
 sky130_fd_sc_hd__a21oi_1 _5337_ (.A1(_1329_),
    .A2(_2215_),
    .B1(_0574_),
    .Y(_2218_));
 sky130_fd_sc_hd__mux2_1 _5338_ (.A0(net525),
    .A1(_2218_),
    .S(net106),
    .X(_0256_));
 sky130_fd_sc_hd__or4_1 _5339_ (.A(net119),
    .B(_0574_),
    .C(_1491_),
    .D(_2214_),
    .X(_2219_));
 sky130_fd_sc_hd__o21ai_1 _5340_ (.A1(net106),
    .A2(_2855_),
    .B1(_2219_),
    .Y(_0257_));
 sky130_fd_sc_hd__or3b_1 _5341_ (.A(_1311_),
    .B(_1312_),
    .C_N(_2201_),
    .X(_2220_));
 sky130_fd_sc_hd__a211o_1 _5342_ (.A1(_0392_),
    .A2(_0405_),
    .B1(_1295_),
    .C1(_1301_),
    .X(_2221_));
 sky130_fd_sc_hd__or4_1 _5343_ (.A(_1299_),
    .B(_1319_),
    .C(_2199_),
    .D(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__a221o_1 _5344_ (.A1(net100),
    .A2(_2220_),
    .B1(_2222_),
    .B2(net160),
    .C1(_2198_),
    .X(_2223_));
 sky130_fd_sc_hd__o21a_1 _5345_ (.A1(_2214_),
    .A2(_2223_),
    .B1(_0575_),
    .X(_2224_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(net535),
    .A1(_2224_),
    .S(net106),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_1 _5347_ (.A(net109),
    .B(_2851_),
    .Y(_2225_));
 sky130_fd_sc_hd__a31o_1 _5348_ (.A1(net162),
    .A2(net109),
    .A3(_0692_),
    .B1(_2225_),
    .X(_0259_));
 sky130_fd_sc_hd__nand2_1 _5349_ (.A(_1350_),
    .B(_1366_),
    .Y(_2226_));
 sky130_fd_sc_hd__mux2_1 _5350_ (.A0(net135),
    .A1(_2226_),
    .S(net106),
    .X(_0260_));
 sky130_fd_sc_hd__mux2_1 _5351_ (.A0(net650),
    .A1(_1365_),
    .S(net106),
    .X(_0261_));
 sky130_fd_sc_hd__o31a_1 _5352_ (.A1(_0604_),
    .A2(_0608_),
    .A3(_0609_),
    .B1(net878),
    .X(_2227_));
 sky130_fd_sc_hd__or2_1 _5353_ (.A(_0611_),
    .B(_2227_),
    .X(_0262_));
 sky130_fd_sc_hd__or2_1 _5354_ (.A(_0612_),
    .B(_0616_),
    .X(_2228_));
 sky130_fd_sc_hd__a2bb2o_1 _5355_ (.A1_N(net139),
    .A2_N(_0629_),
    .B1(_2228_),
    .B2(net666),
    .X(_0263_));
 sky130_fd_sc_hd__a2bb2o_1 _5356_ (.A1_N(_2949_),
    .A2_N(_0629_),
    .B1(_2228_),
    .B2(net785),
    .X(_0264_));
 sky130_fd_sc_hd__o31ai_1 _5357_ (.A1(_2867_),
    .A2(_0452_),
    .A3(_1400_),
    .B1(_1401_),
    .Y(_2229_));
 sky130_fd_sc_hd__mux2_1 _5358_ (.A0(net133),
    .A1(_2229_),
    .S(net106),
    .X(_0265_));
 sky130_fd_sc_hd__or2_1 _5359_ (.A(_0388_),
    .B(_0487_),
    .X(_2230_));
 sky130_fd_sc_hd__and3b_1 _5360_ (.A_N(_0409_),
    .B(_0424_),
    .C(_0433_),
    .X(_2231_));
 sky130_fd_sc_hd__o21ai_1 _5361_ (.A1(net128),
    .A2(_0419_),
    .B1(_2231_),
    .Y(_2232_));
 sky130_fd_sc_hd__a22o_1 _5362_ (.A1(_0543_),
    .A2(_0632_),
    .B1(_2232_),
    .B2(net126),
    .X(_2233_));
 sky130_fd_sc_hd__a32o_1 _5363_ (.A1(net126),
    .A2(net101),
    .A3(_2230_),
    .B1(_2233_),
    .B2(net161),
    .X(_2234_));
 sky130_fd_sc_hd__nand2_4 _5364_ (.A(net116),
    .B(_2234_),
    .Y(_2235_));
 sky130_fd_sc_hd__and3_1 _5365_ (.A(net116),
    .B(\z80.tv80s.di_reg[0] ),
    .C(_1656_),
    .X(_2236_));
 sky130_fd_sc_hd__a21oi_2 _5366_ (.A1(_2831_),
    .A2(\z80.tv80s.i_tv80_core.SP[0] ),
    .B1(_2236_),
    .Y(_2237_));
 sky130_fd_sc_hd__inv_2 _5367_ (.A(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__o31ai_1 _5368_ (.A1(_2831_),
    .A2(\z80.tv80s.di_reg[0] ),
    .A3(_1656_),
    .B1(_2237_),
    .Y(_2239_));
 sky130_fd_sc_hd__and2_4 _5369_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(_2240_));
 sky130_fd_sc_hd__nand2_4 _5370_ (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .B(net115),
    .Y(_2241_));
 sky130_fd_sc_hd__nand2_1 _5371_ (.A(net92),
    .B(_2240_),
    .Y(_2242_));
 sky130_fd_sc_hd__and3_4 _5372_ (.A(_0598_),
    .B(_1550_),
    .C(_1555_),
    .X(_2243_));
 sky130_fd_sc_hd__mux2_1 _5373_ (.A0(net790),
    .A1(net9),
    .S(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__a2bb2o_1 _5374_ (.A1_N(_2239_),
    .A2_N(_2242_),
    .B1(_2244_),
    .B2(net96),
    .X(_2245_));
 sky130_fd_sc_hd__mux2_1 _5375_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_2245_),
    .S(_2235_),
    .X(_2246_));
 sky130_fd_sc_hd__or2_2 _5376_ (.A(_0599_),
    .B(_1660_),
    .X(_2247_));
 sky130_fd_sc_hd__and2_4 _5377_ (.A(_2241_),
    .B(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__a31o_1 _5378_ (.A1(net92),
    .A2(_2235_),
    .A3(_2248_),
    .B1(net119),
    .X(_2249_));
 sky130_fd_sc_hd__a22o_1 _5379_ (.A1(net107),
    .A2(_2246_),
    .B1(_2249_),
    .B2(net790),
    .X(_0266_));
 sky130_fd_sc_hd__or3_4 _5380_ (.A(net115),
    .B(_0870_),
    .C(_0872_),
    .X(_2250_));
 sky130_fd_sc_hd__or2_1 _5381_ (.A(_2831_),
    .B(\z80.tv80s.di_reg[1] ),
    .X(_2251_));
 sky130_fd_sc_hd__mux2_1 _5382_ (.A0(\z80.tv80s.i_tv80_core.SP[1] ),
    .A1(_1700_),
    .S(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(_2252_));
 sky130_fd_sc_hd__and3_1 _5383_ (.A(_2250_),
    .B(_2251_),
    .C(_2252_),
    .X(_2253_));
 sky130_fd_sc_hd__a21o_1 _5384_ (.A1(_2250_),
    .A2(_2251_),
    .B1(_2252_),
    .X(_2254_));
 sky130_fd_sc_hd__nand2b_1 _5385_ (.A_N(_2253_),
    .B(_2254_),
    .Y(_2255_));
 sky130_fd_sc_hd__xnor2_1 _5386_ (.A(_2237_),
    .B(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__inv_2 _5387_ (.A(_2256_),
    .Y(_2257_));
 sky130_fd_sc_hd__a22o_1 _5388_ (.A1(net796),
    .A2(_2248_),
    .B1(_2257_),
    .B2(_2240_),
    .X(_2258_));
 sky130_fd_sc_hd__mux2_1 _5389_ (.A0(net796),
    .A1(net8),
    .S(_2243_),
    .X(_2259_));
 sky130_fd_sc_hd__mux2_1 _5390_ (.A0(_2258_),
    .A1(_2259_),
    .S(net96),
    .X(_2260_));
 sky130_fd_sc_hd__mux2_1 _5391_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_2260_),
    .S(_2235_),
    .X(_2261_));
 sky130_fd_sc_hd__mux2_1 _5392_ (.A0(net796),
    .A1(_2261_),
    .S(net108),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _5393_ (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .B(_2853_),
    .Y(_2262_));
 sky130_fd_sc_hd__mux2_1 _5394_ (.A0(\z80.tv80s.i_tv80_core.SP[2] ),
    .A1(_1720_),
    .S(net116),
    .X(_2263_));
 sky130_fd_sc_hd__and3_1 _5395_ (.A(_2250_),
    .B(_2262_),
    .C(_2263_),
    .X(_2264_));
 sky130_fd_sc_hd__a21o_1 _5396_ (.A1(_2250_),
    .A2(_2262_),
    .B1(_2263_),
    .X(_2265_));
 sky130_fd_sc_hd__and2b_1 _5397_ (.A_N(_2264_),
    .B(_2265_),
    .X(_2266_));
 sky130_fd_sc_hd__a21o_1 _5398_ (.A1(_2238_),
    .A2(_2254_),
    .B1(_2253_),
    .X(_2267_));
 sky130_fd_sc_hd__xnor2_1 _5399_ (.A(_2266_),
    .B(_2267_),
    .Y(_2268_));
 sky130_fd_sc_hd__inv_2 _5400_ (.A(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__a22o_1 _5401_ (.A1(net802),
    .A2(_2248_),
    .B1(_2269_),
    .B2(_2240_),
    .X(_2270_));
 sky130_fd_sc_hd__mux2_1 _5402_ (.A0(net802),
    .A1(net6),
    .S(_2243_),
    .X(_2271_));
 sky130_fd_sc_hd__mux2_1 _5403_ (.A0(_2270_),
    .A1(_2271_),
    .S(net96),
    .X(_2272_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_2272_),
    .S(_2235_),
    .X(_2273_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(net802),
    .A1(_2273_),
    .S(net108),
    .X(_0268_));
 sky130_fd_sc_hd__or2_1 _5406_ (.A(_2831_),
    .B(\z80.tv80s.di_reg[3] ),
    .X(_2274_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(\z80.tv80s.i_tv80_core.SP[3] ),
    .A1(_1737_),
    .S(net116),
    .X(_2275_));
 sky130_fd_sc_hd__nand3_1 _5408_ (.A(_2250_),
    .B(_2274_),
    .C(_2275_),
    .Y(_2276_));
 sky130_fd_sc_hd__a21o_1 _5409_ (.A1(_2250_),
    .A2(_2274_),
    .B1(_2275_),
    .X(_2277_));
 sky130_fd_sc_hd__nand2_1 _5410_ (.A(_2276_),
    .B(_2277_),
    .Y(_2278_));
 sky130_fd_sc_hd__a21o_1 _5411_ (.A1(_2265_),
    .A2(_2267_),
    .B1(_2264_),
    .X(_2279_));
 sky130_fd_sc_hd__xor2_1 _5412_ (.A(_2278_),
    .B(_2279_),
    .X(_2280_));
 sky130_fd_sc_hd__nand2_1 _5413_ (.A(_2240_),
    .B(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__mux2_1 _5414_ (.A0(net150),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .S(_2247_),
    .X(_2282_));
 sky130_fd_sc_hd__o21a_1 _5415_ (.A1(_2240_),
    .A2(_2282_),
    .B1(net92),
    .X(_2283_));
 sky130_fd_sc_hd__mux2_1 _5416_ (.A0(net825),
    .A1(net3),
    .S(_2243_),
    .X(_2284_));
 sky130_fd_sc_hd__a22o_1 _5417_ (.A1(_2281_),
    .A2(_2283_),
    .B1(_2284_),
    .B2(net96),
    .X(_2285_));
 sky130_fd_sc_hd__mux2_1 _5418_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_2285_),
    .S(_2235_),
    .X(_2286_));
 sky130_fd_sc_hd__mux2_1 _5419_ (.A0(net825),
    .A1(_2286_),
    .S(net108),
    .X(_0269_));
 sky130_fd_sc_hd__or2_1 _5420_ (.A(_2831_),
    .B(\z80.tv80s.di_reg[4] ),
    .X(_2287_));
 sky130_fd_sc_hd__mux2_1 _5421_ (.A0(\z80.tv80s.i_tv80_core.SP[4] ),
    .A1(_1754_),
    .S(net115),
    .X(_2288_));
 sky130_fd_sc_hd__and3_1 _5422_ (.A(_2250_),
    .B(_2287_),
    .C(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__a21o_1 _5423_ (.A1(_2250_),
    .A2(_2287_),
    .B1(_2288_),
    .X(_2290_));
 sky130_fd_sc_hd__nand2b_1 _5424_ (.A_N(_2289_),
    .B(_2290_),
    .Y(_2291_));
 sky130_fd_sc_hd__a21bo_1 _5425_ (.A1(_2277_),
    .A2(_2279_),
    .B1_N(_2276_),
    .X(_2292_));
 sky130_fd_sc_hd__xor2_1 _5426_ (.A(_2291_),
    .B(_2292_),
    .X(_2293_));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(_2240_),
    .B(_2293_),
    .Y(_2294_));
 sky130_fd_sc_hd__mux2_1 _5428_ (.A0(net144),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .S(_2247_),
    .X(_2295_));
 sky130_fd_sc_hd__o21a_1 _5429_ (.A1(_2240_),
    .A2(_2295_),
    .B1(net92),
    .X(_2296_));
 sky130_fd_sc_hd__mux2_1 _5430_ (.A0(net823),
    .A1(net2),
    .S(_2243_),
    .X(_2297_));
 sky130_fd_sc_hd__a22o_1 _5431_ (.A1(_2294_),
    .A2(_2296_),
    .B1(_2297_),
    .B2(net97),
    .X(_2298_));
 sky130_fd_sc_hd__mux2_1 _5432_ (.A0(\z80.tv80s.di_reg[4] ),
    .A1(_2298_),
    .S(_2235_),
    .X(_2299_));
 sky130_fd_sc_hd__mux2_1 _5433_ (.A0(net823),
    .A1(_2299_),
    .S(net107),
    .X(_0270_));
 sky130_fd_sc_hd__or2_1 _5434_ (.A(_2831_),
    .B(\z80.tv80s.di_reg[5] ),
    .X(_2300_));
 sky130_fd_sc_hd__mux2_1 _5435_ (.A0(\z80.tv80s.i_tv80_core.SP[5] ),
    .A1(_1772_),
    .S(net115),
    .X(_2301_));
 sky130_fd_sc_hd__and3_1 _5436_ (.A(_2250_),
    .B(_2300_),
    .C(_2301_),
    .X(_2302_));
 sky130_fd_sc_hd__a21o_1 _5437_ (.A1(_2250_),
    .A2(_2300_),
    .B1(_2301_),
    .X(_2303_));
 sky130_fd_sc_hd__and2b_1 _5438_ (.A_N(_2302_),
    .B(_2303_),
    .X(_2304_));
 sky130_fd_sc_hd__a21o_1 _5439_ (.A1(_2290_),
    .A2(_2292_),
    .B1(_2289_),
    .X(_2305_));
 sky130_fd_sc_hd__xnor2_1 _5440_ (.A(_2304_),
    .B(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__nand2_1 _5441_ (.A(_2240_),
    .B(_2306_),
    .Y(_2307_));
 sky130_fd_sc_hd__mux2_1 _5442_ (.A0(net141),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(_2247_),
    .X(_2308_));
 sky130_fd_sc_hd__o21a_1 _5443_ (.A1(_2240_),
    .A2(_2308_),
    .B1(net92),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _5444_ (.A0(net809),
    .A1(net4),
    .S(_2243_),
    .X(_2310_));
 sky130_fd_sc_hd__a22o_1 _5445_ (.A1(_2307_),
    .A2(_2309_),
    .B1(_2310_),
    .B2(net97),
    .X(_2311_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_2311_),
    .S(_2235_),
    .X(_2312_));
 sky130_fd_sc_hd__mux2_1 _5447_ (.A0(net809),
    .A1(_2312_),
    .S(net108),
    .X(_0271_));
 sky130_fd_sc_hd__or2_1 _5448_ (.A(_2831_),
    .B(\z80.tv80s.di_reg[6] ),
    .X(_2313_));
 sky130_fd_sc_hd__mux2_1 _5449_ (.A0(\z80.tv80s.i_tv80_core.SP[6] ),
    .A1(_1790_),
    .S(net116),
    .X(_2314_));
 sky130_fd_sc_hd__and3_1 _5450_ (.A(_2250_),
    .B(_2313_),
    .C(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__a21o_1 _5451_ (.A1(_2250_),
    .A2(_2313_),
    .B1(_2314_),
    .X(_2316_));
 sky130_fd_sc_hd__and2b_1 _5452_ (.A_N(_2315_),
    .B(_2316_),
    .X(_2317_));
 sky130_fd_sc_hd__a21o_1 _5453_ (.A1(_2303_),
    .A2(_2305_),
    .B1(_2302_),
    .X(_2318_));
 sky130_fd_sc_hd__xnor2_1 _5454_ (.A(_2317_),
    .B(_2318_),
    .Y(_2319_));
 sky130_fd_sc_hd__o2bb2a_1 _5455_ (.A1_N(net818),
    .A2_N(_2248_),
    .B1(_2319_),
    .B2(_2241_),
    .X(_2320_));
 sky130_fd_sc_hd__mux2_1 _5456_ (.A0(net818),
    .A1(net5),
    .S(_2243_),
    .X(_2321_));
 sky130_fd_sc_hd__nand2_1 _5457_ (.A(net96),
    .B(_2321_),
    .Y(_2322_));
 sky130_fd_sc_hd__o21ai_1 _5458_ (.A1(net96),
    .A2(_2320_),
    .B1(_2322_),
    .Y(_2323_));
 sky130_fd_sc_hd__mux2_1 _5459_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_2323_),
    .S(_2235_),
    .X(_2324_));
 sky130_fd_sc_hd__mux2_1 _5460_ (.A0(net818),
    .A1(_2324_),
    .S(net107),
    .X(_0272_));
 sky130_fd_sc_hd__a21oi_2 _5461_ (.A1(_2316_),
    .A2(_2318_),
    .B1(_2315_),
    .Y(_2325_));
 sky130_fd_sc_hd__o21a_1 _5462_ (.A1(_2831_),
    .A2(\z80.tv80s.di_reg[7] ),
    .B1(_2250_),
    .X(_2326_));
 sky130_fd_sc_hd__mux2_1 _5463_ (.A0(\z80.tv80s.i_tv80_core.SP[7] ),
    .A1(_1807_),
    .S(net115),
    .X(_2327_));
 sky130_fd_sc_hd__nor2_1 _5464_ (.A(net65),
    .B(_2327_),
    .Y(_2328_));
 sky130_fd_sc_hd__nand2_1 _5465_ (.A(net65),
    .B(_2327_),
    .Y(_2329_));
 sky130_fd_sc_hd__nand2b_1 _5466_ (.A_N(_2328_),
    .B(_2329_),
    .Y(_2330_));
 sky130_fd_sc_hd__xnor2_1 _5467_ (.A(_2325_),
    .B(_2330_),
    .Y(_2331_));
 sky130_fd_sc_hd__o2bb2ai_1 _5468_ (.A1_N(net807),
    .A2_N(_2248_),
    .B1(_2331_),
    .B2(_2241_),
    .Y(_2332_));
 sky130_fd_sc_hd__mux2_1 _5469_ (.A0(net807),
    .A1(net7),
    .S(_2243_),
    .X(_2333_));
 sky130_fd_sc_hd__mux2_1 _5470_ (.A0(_2332_),
    .A1(_2333_),
    .S(net96),
    .X(_2334_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_2334_),
    .S(_2235_),
    .X(_2335_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(net807),
    .A1(_2335_),
    .S(net107),
    .X(_0273_));
 sky130_fd_sc_hd__o21ai_2 _5473_ (.A1(_2325_),
    .A2(_2328_),
    .B1(_2329_),
    .Y(_2336_));
 sky130_fd_sc_hd__mux2_1 _5474_ (.A0(\z80.tv80s.i_tv80_core.SP[8] ),
    .A1(_1826_),
    .S(net115),
    .X(_2337_));
 sky130_fd_sc_hd__and2_1 _5475_ (.A(_2326_),
    .B(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__nor2_1 _5476_ (.A(net65),
    .B(_2337_),
    .Y(_2339_));
 sky130_fd_sc_hd__nor2_1 _5477_ (.A(_2338_),
    .B(_2339_),
    .Y(_2340_));
 sky130_fd_sc_hd__xnor2_1 _5478_ (.A(_2336_),
    .B(_2340_),
    .Y(_2341_));
 sky130_fd_sc_hd__o21ai_1 _5479_ (.A1(net95),
    .A2(_2248_),
    .B1(net739),
    .Y(_2342_));
 sky130_fd_sc_hd__or4_1 _5480_ (.A(net111),
    .B(_2964_),
    .C(_2982_),
    .D(_0514_),
    .X(_2343_));
 sky130_fd_sc_hd__or4_1 _5481_ (.A(_0477_),
    .B(_0507_),
    .C(_0703_),
    .D(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__nor2_1 _5482_ (.A(_2205_),
    .B(_2344_),
    .Y(_2345_));
 sky130_fd_sc_hd__a2bb2o_2 _5483_ (.A1_N(_0514_),
    .A2_N(_0634_),
    .B1(_1663_),
    .B2(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__nand2_4 _5484_ (.A(net116),
    .B(_2346_),
    .Y(_2347_));
 sky130_fd_sc_hd__o311a_1 _5485_ (.A1(net95),
    .A2(_2241_),
    .A3(_2341_),
    .B1(_2342_),
    .C1(_2347_),
    .X(_2348_));
 sky130_fd_sc_hd__a31o_1 _5486_ (.A1(net116),
    .A2(_2852_),
    .A3(_2346_),
    .B1(net118),
    .X(_2349_));
 sky130_fd_sc_hd__a2bb2o_1 _5487_ (.A1_N(_2348_),
    .A2_N(_2349_),
    .B1(net118),
    .B2(net739),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5488_ (.A0(\z80.tv80s.i_tv80_core.SP[9] ),
    .A1(_1843_),
    .S(net115),
    .X(_2350_));
 sky130_fd_sc_hd__xnor2_1 _5489_ (.A(net65),
    .B(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__inv_2 _5490_ (.A(_2351_),
    .Y(_2352_));
 sky130_fd_sc_hd__a21oi_1 _5491_ (.A1(_2336_),
    .A2(_2340_),
    .B1(_2338_),
    .Y(_2353_));
 sky130_fd_sc_hd__xnor2_1 _5492_ (.A(_2351_),
    .B(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__o21ai_1 _5493_ (.A1(net94),
    .A2(_2248_),
    .B1(net600),
    .Y(_2355_));
 sky130_fd_sc_hd__o311a_1 _5494_ (.A1(net94),
    .A2(_2241_),
    .A3(_2354_),
    .B1(_2355_),
    .C1(_2347_),
    .X(_2356_));
 sky130_fd_sc_hd__o21ba_1 _5495_ (.A1(\z80.tv80s.di_reg[1] ),
    .A2(_2347_),
    .B1_N(_2356_),
    .X(_2357_));
 sky130_fd_sc_hd__mux2_1 _5496_ (.A0(net600),
    .A1(_2357_),
    .S(net104),
    .X(_0275_));
 sky130_fd_sc_hd__o21a_1 _5497_ (.A1(_2337_),
    .A2(_2350_),
    .B1(net65),
    .X(_2358_));
 sky130_fd_sc_hd__a31o_1 _5498_ (.A1(_2336_),
    .A2(_2340_),
    .A3(_2352_),
    .B1(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__mux2_1 _5499_ (.A0(\z80.tv80s.i_tv80_core.SP[10] ),
    .A1(_1862_),
    .S(net115),
    .X(_2360_));
 sky130_fd_sc_hd__and2_1 _5500_ (.A(net65),
    .B(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__nor2_1 _5501_ (.A(net65),
    .B(_2360_),
    .Y(_2362_));
 sky130_fd_sc_hd__nor2_1 _5502_ (.A(_2361_),
    .B(_2362_),
    .Y(_2363_));
 sky130_fd_sc_hd__xnor2_1 _5503_ (.A(_2359_),
    .B(_2363_),
    .Y(_2364_));
 sky130_fd_sc_hd__inv_2 _5504_ (.A(_2364_),
    .Y(_2365_));
 sky130_fd_sc_hd__a22o_1 _5505_ (.A1(net775),
    .A2(_2248_),
    .B1(_2365_),
    .B2(_2240_),
    .X(_2366_));
 sky130_fd_sc_hd__mux2_1 _5506_ (.A0(net775),
    .A1(_2366_),
    .S(net91),
    .X(_2367_));
 sky130_fd_sc_hd__mux2_1 _5507_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_2367_),
    .S(_2347_),
    .X(_2368_));
 sky130_fd_sc_hd__mux2_1 _5508_ (.A0(net775),
    .A1(_2368_),
    .S(net104),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5509_ (.A0(\z80.tv80s.i_tv80_core.SP[11] ),
    .A1(_1879_),
    .S(net115),
    .X(_2369_));
 sky130_fd_sc_hd__xor2_1 _5510_ (.A(net65),
    .B(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__a21o_1 _5511_ (.A1(_2359_),
    .A2(_2363_),
    .B1(_2361_),
    .X(_2371_));
 sky130_fd_sc_hd__xnor2_1 _5512_ (.A(_2370_),
    .B(_2371_),
    .Y(_2372_));
 sky130_fd_sc_hd__o2bb2a_1 _5513_ (.A1_N(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2_N(_2248_),
    .B1(_2372_),
    .B2(_2241_),
    .X(_2373_));
 sky130_fd_sc_hd__nand2_1 _5514_ (.A(net741),
    .B(net94),
    .Y(_2374_));
 sky130_fd_sc_hd__o211a_1 _5515_ (.A1(net94),
    .A2(_2373_),
    .B1(_2374_),
    .C1(_2347_),
    .X(_2375_));
 sky130_fd_sc_hd__o21ba_1 _5516_ (.A1(\z80.tv80s.di_reg[3] ),
    .A2(_2347_),
    .B1_N(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__mux2_1 _5517_ (.A0(net741),
    .A1(_2376_),
    .S(net104),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5518_ (.A0(\z80.tv80s.i_tv80_core.SP[12] ),
    .A1(_1898_),
    .S(net115),
    .X(_2377_));
 sky130_fd_sc_hd__and2_1 _5519_ (.A(net65),
    .B(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__or2_1 _5520_ (.A(net65),
    .B(_2377_),
    .X(_2379_));
 sky130_fd_sc_hd__nand2b_1 _5521_ (.A_N(_2378_),
    .B(_2379_),
    .Y(_2380_));
 sky130_fd_sc_hd__o21a_1 _5522_ (.A1(_2360_),
    .A2(_2369_),
    .B1(net65),
    .X(_2381_));
 sky130_fd_sc_hd__a31o_1 _5523_ (.A1(_2359_),
    .A2(_2363_),
    .A3(_2370_),
    .B1(_2381_),
    .X(_2382_));
 sky130_fd_sc_hd__xor2_1 _5524_ (.A(_2380_),
    .B(_2382_),
    .X(_2383_));
 sky130_fd_sc_hd__o2bb2a_1 _5525_ (.A1_N(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2_N(_2248_),
    .B1(_2383_),
    .B2(_2241_),
    .X(_2384_));
 sky130_fd_sc_hd__nand2_1 _5526_ (.A(net729),
    .B(net94),
    .Y(_2385_));
 sky130_fd_sc_hd__o211a_1 _5527_ (.A1(net94),
    .A2(_2384_),
    .B1(_2385_),
    .C1(_2347_),
    .X(_2386_));
 sky130_fd_sc_hd__o21ba_1 _5528_ (.A1(\z80.tv80s.di_reg[4] ),
    .A2(_2347_),
    .B1_N(_2386_),
    .X(_2387_));
 sky130_fd_sc_hd__mux2_1 _5529_ (.A0(net729),
    .A1(_2387_),
    .S(net104),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5530_ (.A0(\z80.tv80s.i_tv80_core.SP[13] ),
    .A1(_1917_),
    .S(net116),
    .X(_2388_));
 sky130_fd_sc_hd__and2_1 _5531_ (.A(net65),
    .B(_2388_),
    .X(_2389_));
 sky130_fd_sc_hd__or2_1 _5532_ (.A(net65),
    .B(_2388_),
    .X(_2390_));
 sky130_fd_sc_hd__and2b_1 _5533_ (.A_N(_2389_),
    .B(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__a21o_1 _5534_ (.A1(_2379_),
    .A2(_2382_),
    .B1(_2378_),
    .X(_2392_));
 sky130_fd_sc_hd__xnor2_1 _5535_ (.A(_2391_),
    .B(_2392_),
    .Y(_2393_));
 sky130_fd_sc_hd__inv_2 _5536_ (.A(_2393_),
    .Y(_2394_));
 sky130_fd_sc_hd__a22o_1 _5537_ (.A1(net794),
    .A2(_2248_),
    .B1(_2394_),
    .B2(_2240_),
    .X(_2395_));
 sky130_fd_sc_hd__mux2_1 _5538_ (.A0(net794),
    .A1(_2395_),
    .S(net91),
    .X(_2396_));
 sky130_fd_sc_hd__mux2_1 _5539_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_2396_),
    .S(_2347_),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _5540_ (.A0(net794),
    .A1(_2397_),
    .S(net104),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5541_ (.A0(\z80.tv80s.i_tv80_core.SP[14] ),
    .A1(_1934_),
    .S(net116),
    .X(_2398_));
 sky130_fd_sc_hd__and2_1 _5542_ (.A(net65),
    .B(_2398_),
    .X(_2399_));
 sky130_fd_sc_hd__or2_1 _5543_ (.A(net65),
    .B(_2398_),
    .X(_2400_));
 sky130_fd_sc_hd__nand2b_1 _5544_ (.A_N(_2399_),
    .B(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__a21o_1 _5545_ (.A1(_2390_),
    .A2(_2392_),
    .B1(_2389_),
    .X(_2402_));
 sky130_fd_sc_hd__xor2_1 _5546_ (.A(_2401_),
    .B(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__o2bb2a_1 _5547_ (.A1_N(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2_N(_2248_),
    .B1(_2403_),
    .B2(_2241_),
    .X(_2404_));
 sky130_fd_sc_hd__nand2_1 _5548_ (.A(net747),
    .B(net94),
    .Y(_2405_));
 sky130_fd_sc_hd__o211a_1 _5549_ (.A1(net94),
    .A2(_2404_),
    .B1(_2405_),
    .C1(_2347_),
    .X(_2406_));
 sky130_fd_sc_hd__o21ba_1 _5550_ (.A1(\z80.tv80s.di_reg[6] ),
    .A2(_2347_),
    .B1_N(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__mux2_1 _5551_ (.A0(net747),
    .A1(_2407_),
    .S(net104),
    .X(_0280_));
 sky130_fd_sc_hd__a21oi_1 _5552_ (.A1(_2400_),
    .A2(_2402_),
    .B1(_2399_),
    .Y(_2408_));
 sky130_fd_sc_hd__mux2_1 _5553_ (.A0(\z80.tv80s.i_tv80_core.SP[15] ),
    .A1(_1953_),
    .S(net116),
    .X(_2409_));
 sky130_fd_sc_hd__xor2_1 _5554_ (.A(net65),
    .B(_2409_),
    .X(_2410_));
 sky130_fd_sc_hd__xnor2_1 _5555_ (.A(_2408_),
    .B(_2410_),
    .Y(_2411_));
 sky130_fd_sc_hd__a22o_1 _5556_ (.A1(net743),
    .A2(_2248_),
    .B1(_2411_),
    .B2(_2240_),
    .X(_2412_));
 sky130_fd_sc_hd__mux2_1 _5557_ (.A0(net743),
    .A1(_2412_),
    .S(net91),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_1 _5558_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_2413_),
    .S(_2347_),
    .X(_2414_));
 sky130_fd_sc_hd__mux2_1 _5559_ (.A0(net743),
    .A1(_2414_),
    .S(net104),
    .X(_0281_));
 sky130_fd_sc_hd__or4_1 _5560_ (.A(net111),
    .B(net122),
    .C(_2937_),
    .D(net96),
    .X(_2415_));
 sky130_fd_sc_hd__xnor2_1 _5561_ (.A(net553),
    .B(_2415_),
    .Y(_0282_));
 sky130_fd_sc_hd__a21o_1 _5562_ (.A1(_0415_),
    .A2(_0483_),
    .B1(_0692_),
    .X(_2416_));
 sky130_fd_sc_hd__or3_1 _5563_ (.A(_0756_),
    .B(_1340_),
    .C(_1357_),
    .X(_2417_));
 sky130_fd_sc_hd__a211o_1 _5564_ (.A1(_2948_),
    .A2(_2416_),
    .B1(_2417_),
    .C1(_0753_),
    .X(_2418_));
 sky130_fd_sc_hd__a32o_1 _5565_ (.A1(net139),
    .A2(_2879_),
    .A3(_1344_),
    .B1(_3008_),
    .B2(net129),
    .X(_2419_));
 sky130_fd_sc_hd__a21oi_1 _5566_ (.A1(_2948_),
    .A2(_1345_),
    .B1(_2419_),
    .Y(_2420_));
 sky130_fd_sc_hd__o2bb2a_1 _5567_ (.A1_N(net160),
    .A2_N(_2418_),
    .B1(_2420_),
    .B2(_0383_),
    .X(_2421_));
 sky130_fd_sc_hd__nor2_2 _5568_ (.A(net123),
    .B(_2421_),
    .Y(_2422_));
 sky130_fd_sc_hd__inv_2 _5569_ (.A(_2422_),
    .Y(_2423_));
 sky130_fd_sc_hd__a31o_1 _5570_ (.A1(_1351_),
    .A2(_1365_),
    .A3(_2422_),
    .B1(net119),
    .X(_2424_));
 sky130_fd_sc_hd__inv_2 _5571_ (.A(_2424_),
    .Y(_2425_));
 sky130_fd_sc_hd__nor2_1 _5572_ (.A(_1365_),
    .B(_2423_),
    .Y(_2426_));
 sky130_fd_sc_hd__a31o_1 _5573_ (.A1(net159),
    .A2(_2940_),
    .A3(_1342_),
    .B1(_1334_),
    .X(_2427_));
 sky130_fd_sc_hd__nand2_1 _5574_ (.A(_2829_),
    .B(_1505_),
    .Y(_2428_));
 sky130_fd_sc_hd__a32o_1 _5575_ (.A1(_0659_),
    .A2(_1497_),
    .A3(_2428_),
    .B1(_1344_),
    .B2(net147),
    .X(_2429_));
 sky130_fd_sc_hd__a211o_1 _5576_ (.A1(_2944_),
    .A2(_1499_),
    .B1(_2429_),
    .C1(_2942_),
    .X(_2430_));
 sky130_fd_sc_hd__o211a_1 _5577_ (.A1(_0423_),
    .A2(_0469_),
    .B1(_1335_),
    .C1(_1354_),
    .X(_2431_));
 sky130_fd_sc_hd__nand2_1 _5578_ (.A(net129),
    .B(_2949_),
    .Y(_2432_));
 sky130_fd_sc_hd__a32o_1 _5579_ (.A1(_0395_),
    .A2(_0415_),
    .A3(_2432_),
    .B1(_1499_),
    .B2(_0511_),
    .X(_2433_));
 sky130_fd_sc_hd__a221o_1 _5580_ (.A1(net156),
    .A2(_2931_),
    .B1(_2935_),
    .B2(_0483_),
    .C1(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__a211o_1 _5581_ (.A1(net87),
    .A2(_0473_),
    .B1(_0662_),
    .C1(_2986_),
    .X(_2435_));
 sky130_fd_sc_hd__a2bb2o_1 _5582_ (.A1_N(_0514_),
    .A2_N(_2431_),
    .B1(_2435_),
    .B2(net130),
    .X(_2436_));
 sky130_fd_sc_hd__a211o_1 _5583_ (.A1(net124),
    .A2(_2977_),
    .B1(_2434_),
    .C1(_2436_),
    .X(_2437_));
 sky130_fd_sc_hd__a22o_1 _5584_ (.A1(net100),
    .A2(_2430_),
    .B1(_2437_),
    .B2(net160),
    .X(_2438_));
 sky130_fd_sc_hd__a22o_4 _5585_ (.A1(net156),
    .A2(_2427_),
    .B1(_2438_),
    .B2(_2819_),
    .X(_2439_));
 sky130_fd_sc_hd__inv_2 _5586_ (.A(_2439_),
    .Y(_2440_));
 sky130_fd_sc_hd__and3_2 _5587_ (.A(_1351_),
    .B(_2426_),
    .C(_2439_),
    .X(_2441_));
 sky130_fd_sc_hd__and3_2 _5588_ (.A(_1350_),
    .B(_2426_),
    .C(_2440_),
    .X(_2442_));
 sky130_fd_sc_hd__and4_2 _5589_ (.A(_1351_),
    .B(_1365_),
    .C(_2423_),
    .D(_2439_),
    .X(_2443_));
 sky130_fd_sc_hd__a221o_1 _5590_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .C1(net72),
    .X(_2444_));
 sky130_fd_sc_hd__a221o_1 _5591_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .C1(net71),
    .X(_2445_));
 sky130_fd_sc_hd__a221o_1 _5592_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .A2(net135),
    .B1(_0814_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .C1(net73),
    .X(_2446_));
 sky130_fd_sc_hd__a221o_1 _5593_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(_0814_),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .C1(_0817_),
    .X(_2447_));
 sky130_fd_sc_hd__a21oi_4 _5594_ (.A1(_1351_),
    .A2(_1365_),
    .B1(_2422_),
    .Y(_2448_));
 sky130_fd_sc_hd__and3_1 _5595_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(net84),
    .C(_2447_),
    .X(_2449_));
 sky130_fd_sc_hd__a221o_1 _5596_ (.A1(_1286_),
    .A2(_1416_),
    .B1(_2446_),
    .B2(_2449_),
    .C1(_2440_),
    .X(_2450_));
 sky130_fd_sc_hd__and3_1 _5597_ (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .B(net84),
    .C(_2445_),
    .X(_2451_));
 sky130_fd_sc_hd__a221o_1 _5598_ (.A1(_0818_),
    .A2(_1286_),
    .B1(_2444_),
    .B2(_2451_),
    .C1(_2439_),
    .X(_2452_));
 sky130_fd_sc_hd__nor2_1 _5599_ (.A(_1351_),
    .B(_2440_),
    .Y(_2453_));
 sky130_fd_sc_hd__and3_2 _5600_ (.A(_1365_),
    .B(_2422_),
    .C(_2453_),
    .X(_2454_));
 sky130_fd_sc_hd__nor2_1 _5601_ (.A(_1350_),
    .B(_2439_),
    .Y(_2455_));
 sky130_fd_sc_hd__and3_2 _5602_ (.A(_1365_),
    .B(_2423_),
    .C(_2455_),
    .X(_2456_));
 sky130_fd_sc_hd__and4_2 _5603_ (.A(_1350_),
    .B(_1365_),
    .C(_2422_),
    .D(_2440_),
    .X(_2457_));
 sky130_fd_sc_hd__a21o_1 _5604_ (.A1(\z80.tv80s.i_tv80_core.SP[8] ),
    .A2(_2453_),
    .B1(_2455_),
    .X(_2458_));
 sky130_fd_sc_hd__a32o_1 _5605_ (.A1(_2448_),
    .A2(_2450_),
    .A3(_2452_),
    .B1(_2442_),
    .B2(\z80.tv80s.i_tv80_core.SP[0] ),
    .X(_2459_));
 sky130_fd_sc_hd__a221o_1 _5606_ (.A1(net138),
    .A2(_2441_),
    .B1(_2443_),
    .B2(\z80.tv80s.i_tv80_core.ACC[0] ),
    .C1(_2459_),
    .X(_2460_));
 sky130_fd_sc_hd__a221o_1 _5607_ (.A1(\z80.tv80s.di_reg[0] ),
    .A2(_2456_),
    .B1(_2458_),
    .B2(_2426_),
    .C1(_2460_),
    .X(_2461_));
 sky130_fd_sc_hd__a221o_1 _5608_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(_2454_),
    .B1(_2457_),
    .B2(net709),
    .C1(_2461_),
    .X(_2462_));
 sky130_fd_sc_hd__a22o_1 _5609_ (.A1(net120),
    .A2(net713),
    .B1(_2425_),
    .B2(_2462_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_2 _5610_ (.A(_2426_),
    .B(_2453_),
    .X(_2463_));
 sky130_fd_sc_hd__a22o_1 _5611_ (.A1(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A2(_2443_),
    .B1(_2463_),
    .B2(\z80.tv80s.i_tv80_core.SP[9] ),
    .X(_2464_));
 sky130_fd_sc_hd__a221o_1 _5612_ (.A1(\z80.tv80s.i_tv80_core.SP[1] ),
    .A2(_2442_),
    .B1(_2457_),
    .B2(\z80.tv80s.i_tv80_core.PC[1] ),
    .C1(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__o221a_1 _5613_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .C1(net71),
    .X(_2466_));
 sky130_fd_sc_hd__o221a_1 _5614_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .C1(net72),
    .X(_2467_));
 sky130_fd_sc_hd__or2_1 _5615_ (.A(_2466_),
    .B(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__mux2_1 _5616_ (.A0(_2468_),
    .A1(_1017_),
    .S(_1286_),
    .X(_2469_));
 sky130_fd_sc_hd__mux2_1 _5617_ (.A0(_2469_),
    .A1(_1426_),
    .S(_2439_),
    .X(_2470_));
 sky130_fd_sc_hd__a22o_1 _5618_ (.A1(\z80.tv80s.i_tv80_core.F[1] ),
    .A2(_2441_),
    .B1(_2448_),
    .B2(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__a221o_1 _5619_ (.A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .A2(_2454_),
    .B1(_2456_),
    .B2(\z80.tv80s.di_reg[1] ),
    .C1(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__or2_1 _5620_ (.A(_2465_),
    .B(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__a22o_1 _5621_ (.A1(net120),
    .A2(net592),
    .B1(_2425_),
    .B2(_2473_),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_1 _5622_ (.A1(\z80.tv80s.di_reg[2] ),
    .A2(_2456_),
    .B1(_2457_),
    .B2(\z80.tv80s.i_tv80_core.PC[2] ),
    .X(_2474_));
 sky130_fd_sc_hd__a221o_1 _5623_ (.A1(\z80.tv80s.i_tv80_core.F[2] ),
    .A2(_2441_),
    .B1(_2454_),
    .B2(\z80.tv80s.i_tv80_core.PC[10] ),
    .C1(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__o221a_1 _5624_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .A2(net134),
    .B1(net76),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .C1(net71),
    .X(_2476_));
 sky130_fd_sc_hd__o221a_1 _5625_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .C1(net72),
    .X(_2477_));
 sky130_fd_sc_hd__or2_1 _5626_ (.A(_2476_),
    .B(_2477_),
    .X(_2478_));
 sky130_fd_sc_hd__mux2_1 _5627_ (.A0(_2478_),
    .A1(_1058_),
    .S(_1286_),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _5628_ (.A0(_2479_),
    .A1(_1438_),
    .S(_2439_),
    .X(_2480_));
 sky130_fd_sc_hd__a22o_1 _5629_ (.A1(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A2(_2443_),
    .B1(_2448_),
    .B2(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__a221o_1 _5630_ (.A1(\z80.tv80s.i_tv80_core.SP[2] ),
    .A2(_2442_),
    .B1(_2463_),
    .B2(\z80.tv80s.i_tv80_core.SP[10] ),
    .C1(_2481_),
    .X(_2482_));
 sky130_fd_sc_hd__or2_1 _5631_ (.A(_2475_),
    .B(_2482_),
    .X(_2483_));
 sky130_fd_sc_hd__a22o_1 _5632_ (.A1(net120),
    .A2(net582),
    .B1(_2425_),
    .B2(_2483_),
    .X(_0285_));
 sky130_fd_sc_hd__o221a_1 _5633_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .A2(net135),
    .B1(net77),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .C1(net71),
    .X(_2484_));
 sky130_fd_sc_hd__o221a_1 _5634_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .A2(net135),
    .B1(net77),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .C1(net73),
    .X(_2485_));
 sky130_fd_sc_hd__or2_1 _5635_ (.A(_2484_),
    .B(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__o221a_1 _5636_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .A2(net134),
    .B1(net76),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .C1(net71),
    .X(_2487_));
 sky130_fd_sc_hd__o221a_1 _5637_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .A2(net135),
    .B1(net76),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .C1(net73),
    .X(_2488_));
 sky130_fd_sc_hd__or2_1 _5638_ (.A(_2487_),
    .B(_2488_),
    .X(_2489_));
 sky130_fd_sc_hd__mux4_2 _5639_ (.A0(_2489_),
    .A1(_2486_),
    .A2(_1099_),
    .A3(_1447_),
    .S0(_2439_),
    .S1(_1286_),
    .X(_2490_));
 sky130_fd_sc_hd__a22o_1 _5640_ (.A1(\z80.tv80s.i_tv80_core.F[3] ),
    .A2(_2441_),
    .B1(_2456_),
    .B2(\z80.tv80s.di_reg[3] ),
    .X(_2491_));
 sky130_fd_sc_hd__a221o_1 _5641_ (.A1(\z80.tv80s.i_tv80_core.SP[3] ),
    .A2(_2442_),
    .B1(_2457_),
    .B2(net612),
    .C1(_2491_),
    .X(_2492_));
 sky130_fd_sc_hd__a22o_1 _5642_ (.A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .A2(_2454_),
    .B1(_2490_),
    .B2(_2448_),
    .X(_2493_));
 sky130_fd_sc_hd__a221o_1 _5643_ (.A1(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A2(_2443_),
    .B1(_2463_),
    .B2(net628),
    .C1(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__or2_1 _5644_ (.A(_2492_),
    .B(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__a22o_1 _5645_ (.A1(net120),
    .A2(net656),
    .B1(_2425_),
    .B2(_2495_),
    .X(_0286_));
 sky130_fd_sc_hd__o221a_1 _5646_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .C1(net71),
    .X(_2496_));
 sky130_fd_sc_hd__o221a_1 _5647_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .C1(net72),
    .X(_2497_));
 sky130_fd_sc_hd__or2_1 _5648_ (.A(_2496_),
    .B(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__o221a_1 _5649_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .A2(net135),
    .B1(net76),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .C1(net71),
    .X(_2499_));
 sky130_fd_sc_hd__o221a_1 _5650_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .A2(net135),
    .B1(net76),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .C1(net73),
    .X(_2500_));
 sky130_fd_sc_hd__or2_1 _5651_ (.A(_2499_),
    .B(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__mux4_1 _5652_ (.A0(_2501_),
    .A1(_2498_),
    .A2(_1145_),
    .A3(_1452_),
    .S0(_2439_),
    .S1(_1286_),
    .X(_2502_));
 sky130_fd_sc_hd__a22o_1 _5653_ (.A1(\z80.tv80s.i_tv80_core.F[4] ),
    .A2(_2441_),
    .B1(_2456_),
    .B2(\z80.tv80s.di_reg[4] ),
    .X(_2503_));
 sky130_fd_sc_hd__a221o_1 _5654_ (.A1(\z80.tv80s.i_tv80_core.SP[4] ),
    .A2(_2442_),
    .B1(_2457_),
    .B2(\z80.tv80s.i_tv80_core.PC[4] ),
    .C1(_2503_),
    .X(_2504_));
 sky130_fd_sc_hd__a22o_1 _5655_ (.A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .A2(_2454_),
    .B1(_2502_),
    .B2(_2448_),
    .X(_2505_));
 sky130_fd_sc_hd__a221o_1 _5656_ (.A1(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A2(_2443_),
    .B1(_2463_),
    .B2(net616),
    .C1(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__or2_1 _5657_ (.A(_2504_),
    .B(_2506_),
    .X(_2507_));
 sky130_fd_sc_hd__a22o_1 _5658_ (.A1(net120),
    .A2(net691),
    .B1(_2425_),
    .B2(_2507_),
    .X(_0287_));
 sky130_fd_sc_hd__o221a_1 _5659_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .C1(net71),
    .X(_2508_));
 sky130_fd_sc_hd__o221a_1 _5660_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .C1(net72),
    .X(_2509_));
 sky130_fd_sc_hd__or2_1 _5661_ (.A(_2508_),
    .B(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__o221a_1 _5662_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .A2(net135),
    .B1(net76),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .C1(net71),
    .X(_2511_));
 sky130_fd_sc_hd__o221a_1 _5663_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .A2(net135),
    .B1(net76),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .C1(net73),
    .X(_2512_));
 sky130_fd_sc_hd__or2_1 _5664_ (.A(_2511_),
    .B(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__mux4_1 _5665_ (.A0(_2513_),
    .A1(_2510_),
    .A2(_1192_),
    .A3(_1458_),
    .S0(_2439_),
    .S1(_1286_),
    .X(_2514_));
 sky130_fd_sc_hd__a22o_1 _5666_ (.A1(\z80.tv80s.i_tv80_core.F[5] ),
    .A2(_2441_),
    .B1(_2456_),
    .B2(\z80.tv80s.di_reg[5] ),
    .X(_2515_));
 sky130_fd_sc_hd__a221o_1 _5667_ (.A1(\z80.tv80s.i_tv80_core.SP[5] ),
    .A2(_2442_),
    .B1(_2457_),
    .B2(\z80.tv80s.i_tv80_core.PC[5] ),
    .C1(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__a22o_1 _5668_ (.A1(\z80.tv80s.i_tv80_core.PC[13] ),
    .A2(_2454_),
    .B1(_2514_),
    .B2(_2448_),
    .X(_2517_));
 sky130_fd_sc_hd__a221o_1 _5669_ (.A1(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A2(_2443_),
    .B1(_2463_),
    .B2(\z80.tv80s.i_tv80_core.SP[13] ),
    .C1(_2517_),
    .X(_2518_));
 sky130_fd_sc_hd__or2_1 _5670_ (.A(_2516_),
    .B(_2518_),
    .X(_2519_));
 sky130_fd_sc_hd__a22o_1 _5671_ (.A1(net120),
    .A2(net674),
    .B1(_2425_),
    .B2(_2519_),
    .X(_0288_));
 sky130_fd_sc_hd__o221a_1 _5672_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(net77),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .C1(_0817_),
    .X(_2520_));
 sky130_fd_sc_hd__o221a_1 _5673_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(net77),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .C1(net73),
    .X(_2521_));
 sky130_fd_sc_hd__or2_1 _5674_ (.A(_2520_),
    .B(_2521_),
    .X(_2522_));
 sky130_fd_sc_hd__o221a_1 _5675_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .C1(net71),
    .X(_2523_));
 sky130_fd_sc_hd__o221a_1 _5676_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .A2(net134),
    .B1(net75),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .C1(net72),
    .X(_2524_));
 sky130_fd_sc_hd__or2_1 _5677_ (.A(_2523_),
    .B(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__mux4_2 _5678_ (.A0(_2525_),
    .A1(_2522_),
    .A2(_1237_),
    .A3(_1465_),
    .S0(_2439_),
    .S1(_1286_),
    .X(_2526_));
 sky130_fd_sc_hd__a22o_1 _5679_ (.A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .A2(_2454_),
    .B1(_2456_),
    .B2(\z80.tv80s.di_reg[6] ),
    .X(_2527_));
 sky130_fd_sc_hd__a221o_1 _5680_ (.A1(\z80.tv80s.i_tv80_core.F[6] ),
    .A2(_2441_),
    .B1(_2463_),
    .B2(\z80.tv80s.i_tv80_core.SP[14] ),
    .C1(_2527_),
    .X(_2528_));
 sky130_fd_sc_hd__a22o_1 _5681_ (.A1(net631),
    .A2(_2442_),
    .B1(_2448_),
    .B2(_2526_),
    .X(_2529_));
 sky130_fd_sc_hd__a221o_1 _5682_ (.A1(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A2(_2443_),
    .B1(_2457_),
    .B2(\z80.tv80s.i_tv80_core.PC[6] ),
    .C1(_2529_),
    .X(_2530_));
 sky130_fd_sc_hd__or2_1 _5683_ (.A(_2528_),
    .B(_2530_),
    .X(_2531_));
 sky130_fd_sc_hd__a22o_1 _5684_ (.A1(net120),
    .A2(net642),
    .B1(_2425_),
    .B2(_2531_),
    .X(_0289_));
 sky130_fd_sc_hd__a22o_1 _5685_ (.A1(\z80.tv80s.i_tv80_core.F[7] ),
    .A2(_2441_),
    .B1(_2442_),
    .B2(\z80.tv80s.i_tv80_core.SP[7] ),
    .X(_2532_));
 sky130_fd_sc_hd__a22o_1 _5686_ (.A1(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A2(_2443_),
    .B1(_2463_),
    .B2(\z80.tv80s.i_tv80_core.SP[15] ),
    .X(_2533_));
 sky130_fd_sc_hd__o221a_1 _5687_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(net77),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .C1(_0817_),
    .X(_2534_));
 sky130_fd_sc_hd__o221a_1 _5688_ (.A1(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .A2(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .B1(net77),
    .B2(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .C1(_0816_),
    .X(_2535_));
 sky130_fd_sc_hd__or2_1 _5689_ (.A(_2534_),
    .B(_2535_),
    .X(_2536_));
 sky130_fd_sc_hd__mux2_1 _5690_ (.A0(_2536_),
    .A1(_1471_),
    .S(_1286_),
    .X(_2537_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(_1293_),
    .A1(_2537_),
    .S(_2439_),
    .X(_2538_));
 sky130_fd_sc_hd__a22o_1 _5692_ (.A1(\z80.tv80s.i_tv80_core.PC[7] ),
    .A2(_2457_),
    .B1(_2538_),
    .B2(_2448_),
    .X(_2539_));
 sky130_fd_sc_hd__a221o_1 _5693_ (.A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .A2(_2454_),
    .B1(_2456_),
    .B2(\z80.tv80s.di_reg[7] ),
    .C1(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__or3_1 _5694_ (.A(_2532_),
    .B(_2533_),
    .C(_2540_),
    .X(_2541_));
 sky130_fd_sc_hd__a22o_1 _5695_ (.A1(net120),
    .A2(net678),
    .B1(_2425_),
    .B2(_2541_),
    .X(_0290_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(_2864_),
    .A1(_0960_),
    .S(net106),
    .X(_2542_));
 sky130_fd_sc_hd__inv_2 _5697_ (.A(_2542_),
    .Y(_0291_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(_2865_),
    .A1(_0947_),
    .S(net106),
    .X(_2543_));
 sky130_fd_sc_hd__inv_2 _5699_ (.A(net571),
    .Y(_0292_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(net240),
    .A1(_0937_),
    .S(net104),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_1 _5701_ (.A0(net232),
    .A1(_0927_),
    .S(net104),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(net228),
    .A1(_0920_),
    .S(net104),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_1 _5703_ (.A0(net222),
    .A1(_0914_),
    .S(net104),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _5704_ (.A0(net220),
    .A1(_0907_),
    .S(net104),
    .X(_0297_));
 sky130_fd_sc_hd__mux2_1 _5705_ (.A0(net224),
    .A1(_0900_),
    .S(net104),
    .X(_0298_));
 sky130_fd_sc_hd__mux2_1 _5706_ (.A0(_2863_),
    .A1(_0893_),
    .S(net104),
    .X(_2544_));
 sky130_fd_sc_hd__inv_2 _5707_ (.A(_2544_),
    .Y(_0299_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(net230),
    .A1(_1011_),
    .S(net105),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _5709_ (.A0(net236),
    .A1(_1023_),
    .S(net104),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(net226),
    .A1(_1093_),
    .S(net105),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_1 _5711_ (.A0(net234),
    .A1(_1110_),
    .S(net105),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _5712_ (.A0(net244),
    .A1(_1185_),
    .S(net105),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _5713_ (.A0(net246),
    .A1(_1199_),
    .S(net105),
    .X(_0305_));
 sky130_fd_sc_hd__mux2_1 _5714_ (.A0(net242),
    .A1(_1244_),
    .S(net105),
    .X(_0306_));
 sky130_fd_sc_hd__or4b_4 _5715_ (.A(_2831_),
    .B(net121),
    .C(_2992_),
    .D_N(_1369_),
    .X(_2545_));
 sky130_fd_sc_hd__mux2_1 _5716_ (.A0(\z80.tv80s.i_tv80_core.ACC[0] ),
    .A1(net614),
    .S(_2545_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_1 _5717_ (.A0(\z80.tv80s.i_tv80_core.ACC[1] ),
    .A1(net594),
    .S(_2545_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_1 _5718_ (.A0(\z80.tv80s.i_tv80_core.ACC[2] ),
    .A1(net633),
    .S(_2545_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_1 _5719_ (.A0(\z80.tv80s.i_tv80_core.ACC[3] ),
    .A1(net701),
    .S(_2545_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_1 _5720_ (.A0(\z80.tv80s.i_tv80_core.ACC[4] ),
    .A1(net719),
    .S(_2545_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_1 _5721_ (.A0(\z80.tv80s.i_tv80_core.ACC[5] ),
    .A1(net751),
    .S(_2545_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_1 _5722_ (.A0(\z80.tv80s.i_tv80_core.ACC[6] ),
    .A1(net622),
    .S(_2545_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_1 _5723_ (.A0(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A1(net777),
    .S(_2545_),
    .X(_0314_));
 sky130_fd_sc_hd__mux2_1 _5724_ (.A0(\z80.tv80s.i_tv80_core.ACC[7] ),
    .A1(net374),
    .S(_1396_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _5725_ (.A(_1315_),
    .B(_1331_),
    .Y(_2546_));
 sky130_fd_sc_hd__mux2_1 _5726_ (.A0(net252),
    .A1(_2546_),
    .S(net106),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _5727_ (.A0(net238),
    .A1(_1330_),
    .S(net106),
    .X(_0317_));
 sky130_fd_sc_hd__or4_1 _5728_ (.A(net773),
    .B(_0473_),
    .C(_0747_),
    .D(_1652_),
    .X(_2547_));
 sky130_fd_sc_hd__a41o_2 _5729_ (.A1(net162),
    .A2(_0706_),
    .A3(_0867_),
    .A4(_1663_),
    .B1(_2547_),
    .X(_2548_));
 sky130_fd_sc_hd__a21oi_4 _5730_ (.A1(net97),
    .A2(_2548_),
    .B1(_0603_),
    .Y(_2549_));
 sky130_fd_sc_hd__a21o_2 _5731_ (.A1(net97),
    .A2(_2548_),
    .B1(_0603_),
    .X(_2550_));
 sky130_fd_sc_hd__o41a_1 _5732_ (.A1(_2888_),
    .A2(_2975_),
    .A3(_0404_),
    .A4(_0689_),
    .B1(net126),
    .X(_2551_));
 sky130_fd_sc_hd__or3b_1 _5733_ (.A(_2964_),
    .B(_2551_),
    .C_N(_2231_),
    .X(_2552_));
 sky130_fd_sc_hd__a32o_1 _5734_ (.A1(_2826_),
    .A2(_0541_),
    .A3(_0632_),
    .B1(_2552_),
    .B2(_0392_),
    .X(_2553_));
 sky130_fd_sc_hd__a31o_4 _5735_ (.A1(net162),
    .A2(_0513_),
    .A3(_0689_),
    .B1(net345),
    .X(_2554_));
 sky130_fd_sc_hd__o21a_1 _5736_ (.A1(net158),
    .A2(_2890_),
    .B1(net123),
    .X(_2555_));
 sky130_fd_sc_hd__a311o_1 _5737_ (.A1(net101),
    .A2(_0388_),
    .A3(_0392_),
    .B1(_2555_),
    .C1(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .X(_2556_));
 sky130_fd_sc_hd__a211o_1 _5738_ (.A1(net161),
    .A2(_2553_),
    .B1(_2554_),
    .C1(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__and2_1 _5739_ (.A(_0598_),
    .B(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__nor2_2 _5740_ (.A(net97),
    .B(_2558_),
    .Y(_2559_));
 sky130_fd_sc_hd__a21oi_4 _5741_ (.A1(net56),
    .A2(net59),
    .B1(_2550_),
    .Y(_2560_));
 sky130_fd_sc_hd__inv_2 _5742_ (.A(_2560_),
    .Y(_2561_));
 sky130_fd_sc_hd__o31a_1 _5743_ (.A1(net112),
    .A2(_2852_),
    .A3(_0690_),
    .B1(_2554_),
    .X(_2562_));
 sky130_fd_sc_hd__nand2b_1 _5744_ (.A_N(_2562_),
    .B(\z80.tv80s.i_tv80_core.PC[0] ),
    .Y(_2563_));
 sky130_fd_sc_hd__xnor2_1 _5745_ (.A(net709),
    .B(_2562_),
    .Y(_2564_));
 sky130_fd_sc_hd__or2_4 _5746_ (.A(_1980_),
    .B(_2558_),
    .X(_2565_));
 sky130_fd_sc_hd__inv_2 _5747_ (.A(_2565_),
    .Y(_2566_));
 sky130_fd_sc_hd__mux2_1 _5748_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A1(net709),
    .S(net90),
    .X(_2567_));
 sky130_fd_sc_hd__a221o_1 _5749_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(net63),
    .B1(net61),
    .B2(_2567_),
    .C1(_1398_),
    .X(_2568_));
 sky130_fd_sc_hd__a22o_1 _5750_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .A2(_1652_),
    .B1(_1657_),
    .B2(_2568_),
    .X(_2569_));
 sky130_fd_sc_hd__o22a_1 _5751_ (.A1(net59),
    .A2(_2564_),
    .B1(_2565_),
    .B2(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__o22a_1 _5752_ (.A1(net709),
    .A2(_2560_),
    .B1(_2570_),
    .B2(_2550_),
    .X(_0318_));
 sky130_fd_sc_hd__o31a_1 _5753_ (.A1(net112),
    .A2(\z80.tv80s.di_reg[1] ),
    .A3(_0690_),
    .B1(_2554_),
    .X(_2571_));
 sky130_fd_sc_hd__and2_1 _5754_ (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .B(_2571_),
    .X(_2572_));
 sky130_fd_sc_hd__xnor2_1 _5755_ (.A(net689),
    .B(_2571_),
    .Y(_2573_));
 sky130_fd_sc_hd__and2_1 _5756_ (.A(_2563_),
    .B(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__nor2_1 _5757_ (.A(_2563_),
    .B(_2573_),
    .Y(_2575_));
 sky130_fd_sc_hd__a21o_1 _5758_ (.A1(\z80.tv80s.i_tv80_core.PC[1] ),
    .A2(net90),
    .B1(_1697_),
    .X(_2576_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(_2576_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .S(net63),
    .X(_2577_));
 sky130_fd_sc_hd__nand2_1 _5760_ (.A(net79),
    .B(_2577_),
    .Y(_2578_));
 sky130_fd_sc_hd__a221o_1 _5761_ (.A1(_2861_),
    .A2(_1652_),
    .B1(_1714_),
    .B2(_2578_),
    .C1(_2565_),
    .X(_2579_));
 sky130_fd_sc_hd__o31ai_1 _5762_ (.A1(net59),
    .A2(_2574_),
    .A3(_2575_),
    .B1(_2579_),
    .Y(_2580_));
 sky130_fd_sc_hd__a22o_1 _5763_ (.A1(net689),
    .A2(_2561_),
    .B1(_2580_),
    .B2(_2549_),
    .X(_0319_));
 sky130_fd_sc_hd__o31a_1 _5764_ (.A1(net112),
    .A2(\z80.tv80s.di_reg[2] ),
    .A3(_0690_),
    .B1(_2554_),
    .X(_2581_));
 sky130_fd_sc_hd__and2_1 _5765_ (.A(net596),
    .B(_2581_),
    .X(_2582_));
 sky130_fd_sc_hd__nor2_1 _5766_ (.A(\z80.tv80s.i_tv80_core.PC[2] ),
    .B(_2581_),
    .Y(_2583_));
 sky130_fd_sc_hd__or2_1 _5767_ (.A(_2582_),
    .B(_2583_),
    .X(_2584_));
 sky130_fd_sc_hd__o21ba_1 _5768_ (.A1(_2572_),
    .A2(_2575_),
    .B1_N(_2584_),
    .X(_2585_));
 sky130_fd_sc_hd__or3b_1 _5769_ (.A(_2572_),
    .B(_2575_),
    .C_N(_2584_),
    .X(_2586_));
 sky130_fd_sc_hd__and2b_1 _5770_ (.A_N(_2585_),
    .B(_2586_),
    .X(_2587_));
 sky130_fd_sc_hd__a21o_1 _5771_ (.A1(\z80.tv80s.i_tv80_core.PC[2] ),
    .A2(net90),
    .B1(_1717_),
    .X(_2588_));
 sky130_fd_sc_hd__mux2_1 _5772_ (.A0(_2588_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .S(_1664_),
    .X(_2589_));
 sky130_fd_sc_hd__nand2_1 _5773_ (.A(net79),
    .B(_2589_),
    .Y(_2590_));
 sky130_fd_sc_hd__o2bb2a_1 _5774_ (.A1_N(_1732_),
    .A2_N(_2590_),
    .B1(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .B2(net67),
    .X(_2591_));
 sky130_fd_sc_hd__o22a_1 _5775_ (.A1(net59),
    .A2(_2587_),
    .B1(_2591_),
    .B2(_2565_),
    .X(_2592_));
 sky130_fd_sc_hd__o22a_1 _5776_ (.A1(net596),
    .A2(_2560_),
    .B1(_2592_),
    .B2(_2550_),
    .X(_0320_));
 sky130_fd_sc_hd__o31a_1 _5777_ (.A1(net112),
    .A2(\z80.tv80s.di_reg[3] ),
    .A3(_0690_),
    .B1(_2554_),
    .X(_2593_));
 sky130_fd_sc_hd__and2_1 _5778_ (.A(net612),
    .B(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__nor2_1 _5779_ (.A(\z80.tv80s.i_tv80_core.PC[3] ),
    .B(_2593_),
    .Y(_2595_));
 sky130_fd_sc_hd__or2_1 _5780_ (.A(_2594_),
    .B(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__o21ba_1 _5781_ (.A1(_2582_),
    .A2(_2585_),
    .B1_N(_2596_),
    .X(_2597_));
 sky130_fd_sc_hd__or3b_1 _5782_ (.A(_2582_),
    .B(_2585_),
    .C_N(_2596_),
    .X(_2598_));
 sky130_fd_sc_hd__and2b_1 _5783_ (.A_N(_2597_),
    .B(_2598_),
    .X(_2599_));
 sky130_fd_sc_hd__mux2_1 _5784_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A1(net612),
    .S(_1668_),
    .X(_2600_));
 sky130_fd_sc_hd__a22o_1 _5785_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(_1664_),
    .B1(net61),
    .B2(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__a21o_1 _5786_ (.A1(net79),
    .A2(_2601_),
    .B1(_1738_),
    .X(_2602_));
 sky130_fd_sc_hd__o21a_1 _5787_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .A2(net67),
    .B1(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__o22a_1 _5788_ (.A1(net59),
    .A2(_2599_),
    .B1(_2603_),
    .B2(_2565_),
    .X(_2604_));
 sky130_fd_sc_hd__o22a_1 _5789_ (.A1(net612),
    .A2(_2560_),
    .B1(_2604_),
    .B2(_2550_),
    .X(_0321_));
 sky130_fd_sc_hd__o31a_1 _5790_ (.A1(net112),
    .A2(\z80.tv80s.di_reg[4] ),
    .A3(_0690_),
    .B1(_2554_),
    .X(_2605_));
 sky130_fd_sc_hd__and2_1 _5791_ (.A(net711),
    .B(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__nor2_1 _5792_ (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .B(_2605_),
    .Y(_2607_));
 sky130_fd_sc_hd__or2_1 _5793_ (.A(_2606_),
    .B(_2607_),
    .X(_2608_));
 sky130_fd_sc_hd__o21ba_1 _5794_ (.A1(_2594_),
    .A2(_2597_),
    .B1_N(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__or3b_1 _5795_ (.A(_2594_),
    .B(_2597_),
    .C_N(_2608_),
    .X(_2610_));
 sky130_fd_sc_hd__and2b_1 _5796_ (.A_N(_2609_),
    .B(_2610_),
    .X(_2611_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A1(\z80.tv80s.i_tv80_core.PC[4] ),
    .S(net90),
    .X(_2612_));
 sky130_fd_sc_hd__a22o_1 _5798_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net63),
    .B1(net61),
    .B2(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__a21o_1 _5799_ (.A1(net79),
    .A2(_2613_),
    .B1(_1755_),
    .X(_2614_));
 sky130_fd_sc_hd__o21a_1 _5800_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .A2(net67),
    .B1(_2614_),
    .X(_2615_));
 sky130_fd_sc_hd__o22a_1 _5801_ (.A1(_2559_),
    .A2(_2611_),
    .B1(_2615_),
    .B2(_2565_),
    .X(_2616_));
 sky130_fd_sc_hd__o22a_1 _5802_ (.A1(net711),
    .A2(_2560_),
    .B1(_2616_),
    .B2(_2550_),
    .X(_0322_));
 sky130_fd_sc_hd__a21o_1 _5803_ (.A1(\z80.tv80s.i_tv80_core.PC[5] ),
    .A2(net90),
    .B1(_1774_),
    .X(_2617_));
 sky130_fd_sc_hd__mux2_1 _5804_ (.A0(_2617_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .S(net63),
    .X(_2618_));
 sky130_fd_sc_hd__a21bo_1 _5805_ (.A1(net79),
    .A2(_2618_),
    .B1_N(_1773_),
    .X(_2619_));
 sky130_fd_sc_hd__mux2_1 _5806_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .A1(_2619_),
    .S(net67),
    .X(_2620_));
 sky130_fd_sc_hd__mux2_1 _5807_ (.A0(_2620_),
    .A1(net769),
    .S(net56),
    .X(_2621_));
 sky130_fd_sc_hd__o31a_1 _5808_ (.A1(net112),
    .A2(\z80.tv80s.di_reg[5] ),
    .A3(_0690_),
    .B1(_2554_),
    .X(_2622_));
 sky130_fd_sc_hd__and2_1 _5809_ (.A(\z80.tv80s.i_tv80_core.PC[5] ),
    .B(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__nor2_1 _5810_ (.A(\z80.tv80s.i_tv80_core.PC[5] ),
    .B(_2622_),
    .Y(_2624_));
 sky130_fd_sc_hd__or2_1 _5811_ (.A(_2623_),
    .B(_2624_),
    .X(_2625_));
 sky130_fd_sc_hd__o21ba_1 _5812_ (.A1(_2606_),
    .A2(_2609_),
    .B1_N(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__or3b_1 _5813_ (.A(_2606_),
    .B(_2609_),
    .C_N(_2625_),
    .X(_2627_));
 sky130_fd_sc_hd__and2b_1 _5814_ (.A_N(_2626_),
    .B(_2627_),
    .X(_2628_));
 sky130_fd_sc_hd__mux2_1 _5815_ (.A0(_2628_),
    .A1(_2621_),
    .S(_2559_),
    .X(_2629_));
 sky130_fd_sc_hd__mux2_1 _5816_ (.A0(net769),
    .A1(_2629_),
    .S(_2549_),
    .X(_0323_));
 sky130_fd_sc_hd__o31a_1 _5817_ (.A1(net112),
    .A2(\z80.tv80s.di_reg[6] ),
    .A3(_0690_),
    .B1(_2554_),
    .X(_2630_));
 sky130_fd_sc_hd__and2_1 _5818_ (.A(\z80.tv80s.i_tv80_core.PC[6] ),
    .B(_2630_),
    .X(_2631_));
 sky130_fd_sc_hd__nor2_1 _5819_ (.A(\z80.tv80s.i_tv80_core.PC[6] ),
    .B(_2630_),
    .Y(_2632_));
 sky130_fd_sc_hd__or2_1 _5820_ (.A(_2631_),
    .B(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__nor2_1 _5821_ (.A(_2623_),
    .B(_2626_),
    .Y(_2634_));
 sky130_fd_sc_hd__o21ba_1 _5822_ (.A1(_2623_),
    .A2(_2626_),
    .B1_N(_2633_),
    .X(_2635_));
 sky130_fd_sc_hd__a21o_1 _5823_ (.A1(_2633_),
    .A2(_2634_),
    .B1(net59),
    .X(_2636_));
 sky130_fd_sc_hd__a21o_1 _5824_ (.A1(\z80.tv80s.i_tv80_core.PC[6] ),
    .A2(net90),
    .B1(_1792_),
    .X(_2637_));
 sky130_fd_sc_hd__mux2_1 _5825_ (.A0(_2637_),
    .A1(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .S(net63),
    .X(_2638_));
 sky130_fd_sc_hd__a21bo_1 _5826_ (.A1(net79),
    .A2(_2638_),
    .B1_N(_1791_),
    .X(_2639_));
 sky130_fd_sc_hd__mux2_1 _5827_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .A1(_2639_),
    .S(net67),
    .X(_2640_));
 sky130_fd_sc_hd__mux2_1 _5828_ (.A0(_2640_),
    .A1(net721),
    .S(net56),
    .X(_2641_));
 sky130_fd_sc_hd__a2bb2o_1 _5829_ (.A1_N(_2635_),
    .A2_N(_2636_),
    .B1(_2641_),
    .B2(net59),
    .X(_2642_));
 sky130_fd_sc_hd__mux2_1 _5830_ (.A0(net721),
    .A1(_2642_),
    .S(_2549_),
    .X(_0324_));
 sky130_fd_sc_hd__o31a_1 _5831_ (.A1(net112),
    .A2(\z80.tv80s.di_reg[7] ),
    .A3(_0690_),
    .B1(_2554_),
    .X(_2643_));
 sky130_fd_sc_hd__and2_1 _5832_ (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .B(net64),
    .X(_2644_));
 sky130_fd_sc_hd__nor2_1 _5833_ (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .B(_2643_),
    .Y(_2645_));
 sky130_fd_sc_hd__or2_1 _5834_ (.A(_2644_),
    .B(_2645_),
    .X(_2646_));
 sky130_fd_sc_hd__o21ba_1 _5835_ (.A1(_2631_),
    .A2(_2635_),
    .B1_N(_2646_),
    .X(_2647_));
 sky130_fd_sc_hd__or3b_1 _5836_ (.A(_2631_),
    .B(_2635_),
    .C_N(_2646_),
    .X(_2648_));
 sky130_fd_sc_hd__and2b_1 _5837_ (.A_N(_2647_),
    .B(_2648_),
    .X(_2649_));
 sky130_fd_sc_hd__mux2_1 _5838_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(\z80.tv80s.i_tv80_core.PC[7] ),
    .S(net90),
    .X(_2650_));
 sky130_fd_sc_hd__a22o_1 _5839_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A2(net63),
    .B1(net60),
    .B2(_2650_),
    .X(_2651_));
 sky130_fd_sc_hd__a21bo_1 _5840_ (.A1(net78),
    .A2(_2651_),
    .B1_N(_1808_),
    .X(_2652_));
 sky130_fd_sc_hd__mux2_1 _5841_ (.A0(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .A1(_2652_),
    .S(net66),
    .X(_2653_));
 sky130_fd_sc_hd__mux2_1 _5842_ (.A0(_2653_),
    .A1(net755),
    .S(net56),
    .X(_2654_));
 sky130_fd_sc_hd__mux2_1 _5843_ (.A0(_2649_),
    .A1(_2654_),
    .S(net59),
    .X(_2655_));
 sky130_fd_sc_hd__mux2_1 _5844_ (.A0(net755),
    .A1(_2655_),
    .S(_2549_),
    .X(_0325_));
 sky130_fd_sc_hd__xnor2_1 _5845_ (.A(net812),
    .B(net64),
    .Y(_2656_));
 sky130_fd_sc_hd__or2_1 _5846_ (.A(_2644_),
    .B(_2647_),
    .X(_2657_));
 sky130_fd_sc_hd__o21ba_1 _5847_ (.A1(_2644_),
    .A2(_2647_),
    .B1_N(_2656_),
    .X(_2658_));
 sky130_fd_sc_hd__xnor2_1 _5848_ (.A(_2656_),
    .B(_2657_),
    .Y(_2659_));
 sky130_fd_sc_hd__mux2_1 _5849_ (.A0(\z80.tv80s.i_tv80_core.I[0] ),
    .A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .S(net90),
    .X(_2660_));
 sky130_fd_sc_hd__a22o_1 _5850_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .A2(net62),
    .B1(net61),
    .B2(_2660_),
    .X(_2661_));
 sky130_fd_sc_hd__a21bo_1 _5851_ (.A1(net78),
    .A2(_2661_),
    .B1_N(_1827_),
    .X(_2662_));
 sky130_fd_sc_hd__mux2_1 _5852_ (.A0(\z80.tv80s.di_reg[0] ),
    .A1(_2662_),
    .S(net67),
    .X(_2663_));
 sky130_fd_sc_hd__mux2_1 _5853_ (.A0(_2663_),
    .A1(net812),
    .S(net56),
    .X(_2664_));
 sky130_fd_sc_hd__mux2_1 _5854_ (.A0(_2659_),
    .A1(_2664_),
    .S(net59),
    .X(_2665_));
 sky130_fd_sc_hd__mux2_1 _5855_ (.A0(net812),
    .A1(_2665_),
    .S(_2549_),
    .X(_0326_));
 sky130_fd_sc_hd__xor2_2 _5856_ (.A(net820),
    .B(net64),
    .X(_2666_));
 sky130_fd_sc_hd__a21o_1 _5857_ (.A1(net812),
    .A2(net64),
    .B1(_2658_),
    .X(_2667_));
 sky130_fd_sc_hd__xnor2_1 _5858_ (.A(_2666_),
    .B(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__mux2_1 _5859_ (.A0(\z80.tv80s.i_tv80_core.I[1] ),
    .A1(\z80.tv80s.i_tv80_core.PC[9] ),
    .S(net89),
    .X(_2669_));
 sky130_fd_sc_hd__a22o_1 _5860_ (.A1(net600),
    .A2(net62),
    .B1(net60),
    .B2(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__a21bo_1 _5861_ (.A1(net78),
    .A2(_2670_),
    .B1_N(_1844_),
    .X(_2671_));
 sky130_fd_sc_hd__mux2_1 _5862_ (.A0(\z80.tv80s.di_reg[1] ),
    .A1(_2671_),
    .S(net66),
    .X(_2672_));
 sky130_fd_sc_hd__a2bb2o_1 _5863_ (.A1_N(net59),
    .A2_N(_2668_),
    .B1(_2672_),
    .B2(_2566_),
    .X(_2673_));
 sky130_fd_sc_hd__a22o_1 _5864_ (.A1(net820),
    .A2(_2561_),
    .B1(_2673_),
    .B2(_2549_),
    .X(_0327_));
 sky130_fd_sc_hd__xnor2_1 _5865_ (.A(net800),
    .B(net64),
    .Y(_2674_));
 sky130_fd_sc_hd__o21a_1 _5866_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(\z80.tv80s.i_tv80_core.PC[9] ),
    .B1(net64),
    .X(_2675_));
 sky130_fd_sc_hd__a21o_1 _5867_ (.A1(_2658_),
    .A2(_2666_),
    .B1(_2675_),
    .X(_2676_));
 sky130_fd_sc_hd__and2b_1 _5868_ (.A_N(_2674_),
    .B(_2676_),
    .X(_2677_));
 sky130_fd_sc_hd__xnor2_1 _5869_ (.A(_2674_),
    .B(_2676_),
    .Y(_2678_));
 sky130_fd_sc_hd__mux2_1 _5870_ (.A0(\z80.tv80s.i_tv80_core.I[2] ),
    .A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .S(net89),
    .X(_2679_));
 sky130_fd_sc_hd__a22o_1 _5871_ (.A1(net775),
    .A2(net62),
    .B1(net60),
    .B2(_2679_),
    .X(_2680_));
 sky130_fd_sc_hd__a21bo_1 _5872_ (.A1(net78),
    .A2(_2680_),
    .B1_N(_1863_),
    .X(_2681_));
 sky130_fd_sc_hd__mux2_1 _5873_ (.A0(\z80.tv80s.di_reg[2] ),
    .A1(_2681_),
    .S(net66),
    .X(_2682_));
 sky130_fd_sc_hd__o22a_1 _5874_ (.A1(net59),
    .A2(_2678_),
    .B1(_2682_),
    .B2(_2565_),
    .X(_2683_));
 sky130_fd_sc_hd__o22a_1 _5875_ (.A1(net800),
    .A2(_2560_),
    .B1(_2683_),
    .B2(_2550_),
    .X(_0328_));
 sky130_fd_sc_hd__xnor2_1 _5876_ (.A(net792),
    .B(net64),
    .Y(_2684_));
 sky130_fd_sc_hd__a21o_1 _5877_ (.A1(\z80.tv80s.i_tv80_core.PC[10] ),
    .A2(net64),
    .B1(_2677_),
    .X(_2685_));
 sky130_fd_sc_hd__xnor2_1 _5878_ (.A(_2684_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__mux2_1 _5879_ (.A0(\z80.tv80s.i_tv80_core.I[3] ),
    .A1(\z80.tv80s.i_tv80_core.PC[11] ),
    .S(net89),
    .X(_2687_));
 sky130_fd_sc_hd__a22o_1 _5880_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .A2(net62),
    .B1(net60),
    .B2(_2687_),
    .X(_2688_));
 sky130_fd_sc_hd__a21bo_1 _5881_ (.A1(net78),
    .A2(_2688_),
    .B1_N(_1880_),
    .X(_2689_));
 sky130_fd_sc_hd__mux2_1 _5882_ (.A0(\z80.tv80s.di_reg[3] ),
    .A1(_2689_),
    .S(net66),
    .X(_2690_));
 sky130_fd_sc_hd__mux2_1 _5883_ (.A0(_2690_),
    .A1(net792),
    .S(net56),
    .X(_2691_));
 sky130_fd_sc_hd__mux2_1 _5884_ (.A0(_2686_),
    .A1(_2691_),
    .S(net59),
    .X(_2692_));
 sky130_fd_sc_hd__mux2_1 _5885_ (.A0(net792),
    .A1(_2692_),
    .S(_2549_),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _5886_ (.A(net764),
    .B(net64),
    .Y(_2693_));
 sky130_fd_sc_hd__or2_1 _5887_ (.A(net764),
    .B(net64),
    .X(_2694_));
 sky130_fd_sc_hd__nand2_1 _5888_ (.A(_2693_),
    .B(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__nor2_1 _5889_ (.A(_2674_),
    .B(_2684_),
    .Y(_2696_));
 sky130_fd_sc_hd__o41a_1 _5890_ (.A1(\z80.tv80s.i_tv80_core.PC[8] ),
    .A2(\z80.tv80s.i_tv80_core.PC[9] ),
    .A3(\z80.tv80s.i_tv80_core.PC[10] ),
    .A4(\z80.tv80s.i_tv80_core.PC[11] ),
    .B1(net64),
    .X(_2697_));
 sky130_fd_sc_hd__a31o_1 _5891_ (.A1(_2658_),
    .A2(_2666_),
    .A3(_2696_),
    .B1(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__xnor2_1 _5892_ (.A(_2695_),
    .B(_2698_),
    .Y(_2699_));
 sky130_fd_sc_hd__mux2_1 _5893_ (.A0(\z80.tv80s.i_tv80_core.I[4] ),
    .A1(\z80.tv80s.i_tv80_core.PC[12] ),
    .S(net89),
    .X(_2700_));
 sky130_fd_sc_hd__a22o_1 _5894_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .A2(net62),
    .B1(net60),
    .B2(_2700_),
    .X(_2701_));
 sky130_fd_sc_hd__a21bo_1 _5895_ (.A1(net78),
    .A2(_2701_),
    .B1_N(_1899_),
    .X(_2702_));
 sky130_fd_sc_hd__mux2_1 _5896_ (.A0(\z80.tv80s.di_reg[4] ),
    .A1(_2702_),
    .S(net66),
    .X(_2703_));
 sky130_fd_sc_hd__mux2_1 _5897_ (.A0(_2703_),
    .A1(net764),
    .S(net56),
    .X(_2704_));
 sky130_fd_sc_hd__mux2_1 _5898_ (.A0(_2699_),
    .A1(_2704_),
    .S(net59),
    .X(_2705_));
 sky130_fd_sc_hd__mux2_1 _5899_ (.A0(net764),
    .A1(_2705_),
    .S(_2549_),
    .X(_0330_));
 sky130_fd_sc_hd__mux2_1 _5900_ (.A0(\z80.tv80s.i_tv80_core.I[5] ),
    .A1(\z80.tv80s.i_tv80_core.PC[13] ),
    .S(net89),
    .X(_2706_));
 sky130_fd_sc_hd__a22o_1 _5901_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .A2(net62),
    .B1(net60),
    .B2(_2706_),
    .X(_2707_));
 sky130_fd_sc_hd__a21bo_1 _5902_ (.A1(net78),
    .A2(_2707_),
    .B1_N(_1918_),
    .X(_2708_));
 sky130_fd_sc_hd__mux2_1 _5903_ (.A0(\z80.tv80s.di_reg[5] ),
    .A1(_2708_),
    .S(net66),
    .X(_2709_));
 sky130_fd_sc_hd__nand2_1 _5904_ (.A(net727),
    .B(net64),
    .Y(_2710_));
 sky130_fd_sc_hd__nor2_1 _5905_ (.A(net727),
    .B(net64),
    .Y(_2711_));
 sky130_fd_sc_hd__inv_2 _5906_ (.A(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(_2710_),
    .B(_2712_),
    .Y(_2713_));
 sky130_fd_sc_hd__a21boi_2 _5908_ (.A1(_2694_),
    .A2(_2698_),
    .B1_N(_2693_),
    .Y(_2714_));
 sky130_fd_sc_hd__nor2_1 _5909_ (.A(_2713_),
    .B(_2714_),
    .Y(_2715_));
 sky130_fd_sc_hd__a21o_1 _5910_ (.A1(_2713_),
    .A2(_2714_),
    .B1(net59),
    .X(_2716_));
 sky130_fd_sc_hd__a2bb2o_1 _5911_ (.A1_N(_2715_),
    .A2_N(_2716_),
    .B1(_2566_),
    .B2(_2709_),
    .X(_2717_));
 sky130_fd_sc_hd__a22o_1 _5912_ (.A1(net727),
    .A2(_2561_),
    .B1(_2717_),
    .B2(_2549_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _5913_ (.A(net735),
    .B(net64),
    .Y(_2718_));
 sky130_fd_sc_hd__or2_1 _5914_ (.A(net735),
    .B(net64),
    .X(_2719_));
 sky130_fd_sc_hd__nand2_1 _5915_ (.A(_2718_),
    .B(_2719_),
    .Y(_2720_));
 sky130_fd_sc_hd__o21ai_1 _5916_ (.A1(_2711_),
    .A2(_2714_),
    .B1(_2710_),
    .Y(_2721_));
 sky130_fd_sc_hd__xnor2_1 _5917_ (.A(_2720_),
    .B(_2721_),
    .Y(_2722_));
 sky130_fd_sc_hd__mux2_1 _5918_ (.A0(\z80.tv80s.i_tv80_core.I[6] ),
    .A1(\z80.tv80s.i_tv80_core.PC[14] ),
    .S(net89),
    .X(_2723_));
 sky130_fd_sc_hd__a22o_1 _5919_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .A2(net62),
    .B1(net60),
    .B2(_2723_),
    .X(_2724_));
 sky130_fd_sc_hd__a21bo_1 _5920_ (.A1(net78),
    .A2(_2724_),
    .B1_N(_1935_),
    .X(_2725_));
 sky130_fd_sc_hd__mux2_1 _5921_ (.A0(\z80.tv80s.di_reg[6] ),
    .A1(_2725_),
    .S(net66),
    .X(_2726_));
 sky130_fd_sc_hd__o22a_1 _5922_ (.A1(net59),
    .A2(_2722_),
    .B1(_2726_),
    .B2(_2565_),
    .X(_2727_));
 sky130_fd_sc_hd__o22a_1 _5923_ (.A1(net735),
    .A2(_2560_),
    .B1(_2727_),
    .B2(_2550_),
    .X(_0332_));
 sky130_fd_sc_hd__a21bo_1 _5924_ (.A1(_2719_),
    .A2(_2721_),
    .B1_N(_2718_),
    .X(_2728_));
 sky130_fd_sc_hd__xor2_1 _5925_ (.A(net759),
    .B(_2728_),
    .X(_2729_));
 sky130_fd_sc_hd__xor2_1 _5926_ (.A(net64),
    .B(_2729_),
    .X(_2730_));
 sky130_fd_sc_hd__mux2_1 _5927_ (.A0(\z80.tv80s.i_tv80_core.I[7] ),
    .A1(\z80.tv80s.i_tv80_core.PC[15] ),
    .S(net89),
    .X(_2731_));
 sky130_fd_sc_hd__a22o_1 _5928_ (.A1(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .A2(net62),
    .B1(net60),
    .B2(_2731_),
    .X(_2732_));
 sky130_fd_sc_hd__a21bo_1 _5929_ (.A1(net78),
    .A2(_2732_),
    .B1_N(_1954_),
    .X(_2733_));
 sky130_fd_sc_hd__mux2_1 _5930_ (.A0(\z80.tv80s.di_reg[7] ),
    .A1(_2733_),
    .S(net66),
    .X(_2734_));
 sky130_fd_sc_hd__mux2_1 _5931_ (.A0(_2734_),
    .A1(net759),
    .S(net56),
    .X(_2735_));
 sky130_fd_sc_hd__mux2_1 _5932_ (.A0(_2730_),
    .A1(_2735_),
    .S(net59),
    .X(_2736_));
 sky130_fd_sc_hd__mux2_1 _5933_ (.A0(net759),
    .A1(_2736_),
    .S(_2549_),
    .X(_0333_));
 sky130_fd_sc_hd__and2_1 _5934_ (.A(net781),
    .B(_0035_),
    .X(_2737_));
 sky130_fd_sc_hd__and2_1 _5935_ (.A(net123),
    .B(net837),
    .X(_2738_));
 sky130_fd_sc_hd__nor2_1 _5936_ (.A(net781),
    .B(net855),
    .Y(_2739_));
 sky130_fd_sc_hd__nor2_1 _5937_ (.A(_2819_),
    .B(net837),
    .Y(_2740_));
 sky130_fd_sc_hd__a221o_1 _5938_ (.A1(net782),
    .A2(_2738_),
    .B1(_2739_),
    .B2(_2740_),
    .C1(_0729_),
    .X(_2741_));
 sky130_fd_sc_hd__a22o_1 _5939_ (.A1(net127),
    .A2(_0730_),
    .B1(_0732_),
    .B2(_2741_),
    .X(_0334_));
 sky130_fd_sc_hd__o31a_1 _5940_ (.A1(_2866_),
    .A2(net855),
    .A3(net837),
    .B1(net123),
    .X(_2742_));
 sky130_fd_sc_hd__nor2_1 _5941_ (.A(_2954_),
    .B(_2742_),
    .Y(_2743_));
 sky130_fd_sc_hd__a32o_1 _5942_ (.A1(_0728_),
    .A2(_0732_),
    .A3(_2743_),
    .B1(_0730_),
    .B2(net124),
    .X(_0335_));
 sky130_fd_sc_hd__a32o_1 _5943_ (.A1(_2866_),
    .A2(net855),
    .A3(_2740_),
    .B1(net124),
    .B2(_2819_),
    .X(_2744_));
 sky130_fd_sc_hd__a32o_1 _5944_ (.A1(_0728_),
    .A2(_0732_),
    .A3(net856),
    .B1(_0730_),
    .B2(net640),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _5945_ (.A1(_2819_),
    .A2(net640),
    .B1(net782),
    .B2(_2740_),
    .X(_2745_));
 sky130_fd_sc_hd__a32o_1 _5946_ (.A1(_0728_),
    .A2(_0732_),
    .A3(net783),
    .B1(_0730_),
    .B2(net761),
    .X(_0337_));
 sky130_fd_sc_hd__a22o_1 _5947_ (.A1(_2819_),
    .A2(net761),
    .B1(_2738_),
    .B2(_2739_),
    .X(_2746_));
 sky130_fd_sc_hd__a32o_1 _5948_ (.A1(_0728_),
    .A2(_0732_),
    .A3(net762),
    .B1(_0730_),
    .B2(net542),
    .X(_0338_));
 sky130_fd_sc_hd__and3b_1 _5949_ (.A_N(_0035_),
    .B(_2738_),
    .C(net781),
    .X(_2747_));
 sky130_fd_sc_hd__a31oi_1 _5950_ (.A1(_2819_),
    .A2(net542),
    .A3(_0727_),
    .B1(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__o2bb2a_1 _5951_ (.A1_N(_0732_),
    .A2_N(_2748_),
    .B1(net845),
    .B2(_0731_),
    .X(_0339_));
 sky130_fd_sc_hd__nor2_1 _5952_ (.A(_2819_),
    .B(_0731_),
    .Y(_2749_));
 sky130_fd_sc_hd__a31o_1 _5953_ (.A1(_2866_),
    .A2(_0035_),
    .A3(net837),
    .B1(_2819_),
    .X(_2750_));
 sky130_fd_sc_hd__a41o_1 _5954_ (.A1(_0594_),
    .A2(_0728_),
    .A3(_0732_),
    .A4(net838),
    .B1(_2749_),
    .X(_0340_));
 sky130_fd_sc_hd__a21bo_1 _5955_ (.A1(net648),
    .A2(_0733_),
    .B1_N(_0745_),
    .X(_0341_));
 sky130_fd_sc_hd__nor2_1 _5956_ (.A(_0574_),
    .B(_0578_),
    .Y(_2751_));
 sky130_fd_sc_hd__o21a_1 _5957_ (.A1(net121),
    .A2(_2751_),
    .B1(net567),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_1 _5958_ (.A1(\z80.tv80s.i_tv80_core.NMICycle ),
    .A2(_0733_),
    .B1(_0734_),
    .B2(net484),
    .X(_0343_));
 sky130_fd_sc_hd__or2_4 _5959_ (.A(_0888_),
    .B(_1414_),
    .X(_2752_));
 sky130_fd_sc_hd__mux2_1 _5960_ (.A0(_1419_),
    .A1(net519),
    .S(_2752_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_1 _5961_ (.A0(_1431_),
    .A1(net456),
    .S(_2752_),
    .X(_0345_));
 sky130_fd_sc_hd__mux2_1 _5962_ (.A0(_1442_),
    .A1(net347),
    .S(_2752_),
    .X(_0346_));
 sky130_fd_sc_hd__mux2_1 _5963_ (.A0(_1448_),
    .A1(net518),
    .S(_2752_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _5964_ (.A0(_1453_),
    .A1(net517),
    .S(_2752_),
    .X(_0348_));
 sky130_fd_sc_hd__mux2_1 _5965_ (.A0(_1459_),
    .A1(net508),
    .S(_2752_),
    .X(_0349_));
 sky130_fd_sc_hd__mux2_1 _5966_ (.A0(_1466_),
    .A1(net453),
    .S(_2752_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _5967_ (.A0(_1472_),
    .A1(net522),
    .S(_2752_),
    .X(_0351_));
 sky130_fd_sc_hd__mux2_1 _5968_ (.A0(net9),
    .A1(net854),
    .S(_0599_),
    .X(_0352_));
 sky130_fd_sc_hd__mux2_1 _5969_ (.A0(net8),
    .A1(net849),
    .S(_0599_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _5970_ (.A0(net6),
    .A1(net848),
    .S(_0599_),
    .X(_0354_));
 sky130_fd_sc_hd__mux2_1 _5971_ (.A0(net3),
    .A1(net858),
    .S(_0599_),
    .X(_0355_));
 sky130_fd_sc_hd__mux2_1 _5972_ (.A0(net2),
    .A1(net862),
    .S(_0599_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_1 _5973_ (.A0(net4),
    .A1(net859),
    .S(_0599_),
    .X(_0357_));
 sky130_fd_sc_hd__mux2_1 _5974_ (.A0(net5),
    .A1(net860),
    .S(_0599_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _5975_ (.A0(net7),
    .A1(net861),
    .S(_0599_),
    .X(_0359_));
 sky130_fd_sc_hd__a2bb2o_1 _5976_ (.A1_N(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .A2_N(_0714_),
    .B1(_0557_),
    .B2(_2834_),
    .X(_2753_));
 sky130_fd_sc_hd__mux2_1 _5977_ (.A0(net567),
    .A1(_2753_),
    .S(_0574_),
    .X(_2754_));
 sky130_fd_sc_hd__or2_4 _5978_ (.A(_0579_),
    .B(net568),
    .X(_2755_));
 sky130_fd_sc_hd__nor2_2 _5979_ (.A(_0575_),
    .B(_2755_),
    .Y(_2756_));
 sky130_fd_sc_hd__a22o_1 _5980_ (.A1(\z80.tv80s.i_tv80_core.ts[0] ),
    .A2(_2755_),
    .B1(_2756_),
    .B2(net523),
    .X(_0360_));
 sky130_fd_sc_hd__or2_1 _5981_ (.A(net635),
    .B(_0572_),
    .X(_2757_));
 sky130_fd_sc_hd__mux2_1 _5982_ (.A0(_2757_),
    .A1(net768),
    .S(_2755_),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_1 _5983_ (.A1(net117),
    .A2(_2755_),
    .B1(_2756_),
    .B2(net768),
    .X(_0362_));
 sky130_fd_sc_hd__a22o_1 _5984_ (.A1(net115),
    .A2(_2755_),
    .B1(_2756_),
    .B2(net117),
    .X(_0363_));
 sky130_fd_sc_hd__a22o_1 _5985_ (.A1(net486),
    .A2(_2755_),
    .B1(_2756_),
    .B2(net115),
    .X(_0364_));
 sky130_fd_sc_hd__a22o_1 _5986_ (.A1(net481),
    .A2(_2755_),
    .B1(_2756_),
    .B2(net486),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_1 _5987_ (.A1(net894),
    .A2(_2755_),
    .B1(_2756_),
    .B2(net481),
    .X(_0366_));
 sky130_fd_sc_hd__or3_1 _5988_ (.A(net511),
    .B(net525),
    .C(_2855_),
    .X(_2758_));
 sky130_fd_sc_hd__or4b_1 _5989_ (.A(net630),
    .B(_2856_),
    .C(_2758_),
    .D_N(_0788_),
    .X(_2759_));
 sky130_fd_sc_hd__a21o_1 _5990_ (.A1(net128),
    .A2(\z80.tv80s.i_tv80_core.ts[4] ),
    .B1(_0598_),
    .X(_2760_));
 sky130_fd_sc_hd__and2_4 _5991_ (.A(_0770_),
    .B(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__inv_2 _5992_ (.A(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__a21o_2 _5993_ (.A1(net81),
    .A2(_2762_),
    .B1(net95),
    .X(_2763_));
 sky130_fd_sc_hd__inv_2 _5994_ (.A(_2763_),
    .Y(_2764_));
 sky130_fd_sc_hd__a21oi_4 _5995_ (.A1(net74),
    .A2(_2763_),
    .B1(net118),
    .Y(_2765_));
 sky130_fd_sc_hd__o2bb2a_1 _5996_ (.A1_N(_2239_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1656_),
    .X(_2766_));
 sky130_fd_sc_hd__o21a_1 _5997_ (.A1(net96),
    .A2(_2766_),
    .B1(net74),
    .X(_2767_));
 sky130_fd_sc_hd__nor2_1 _5998_ (.A(_0863_),
    .B(net74),
    .Y(_2768_));
 sky130_fd_sc_hd__o32a_1 _5999_ (.A1(net119),
    .A2(_2767_),
    .A3(_2768_),
    .B1(net715),
    .B2(_2765_),
    .X(_0367_));
 sky130_fd_sc_hd__o22a_1 _6000_ (.A1(net81),
    .A2(_1700_),
    .B1(_2257_),
    .B2(_2762_),
    .X(_2769_));
 sky130_fd_sc_hd__o21a_1 _6001_ (.A1(net96),
    .A2(_2769_),
    .B1(net74),
    .X(_2770_));
 sky130_fd_sc_hd__nor2_1 _6002_ (.A(_1003_),
    .B(net74),
    .Y(_2771_));
 sky130_fd_sc_hd__o32a_1 _6003_ (.A1(net119),
    .A2(_2770_),
    .A3(_2771_),
    .B1(net654),
    .B2(_2765_),
    .X(_0368_));
 sky130_fd_sc_hd__o22a_1 _6004_ (.A1(_1397_),
    .A2(_1720_),
    .B1(_2269_),
    .B2(_2762_),
    .X(_2772_));
 sky130_fd_sc_hd__o21a_1 _6005_ (.A1(net96),
    .A2(_2772_),
    .B1(net74),
    .X(_2773_));
 sky130_fd_sc_hd__nor2_1 _6006_ (.A(_1053_),
    .B(net74),
    .Y(_2774_));
 sky130_fd_sc_hd__o32a_1 _6007_ (.A1(net119),
    .A2(_2773_),
    .A3(_2774_),
    .B1(net652),
    .B2(_2765_),
    .X(_0369_));
 sky130_fd_sc_hd__o2bb2a_1 _6008_ (.A1_N(_2280_),
    .A2_N(_2761_),
    .B1(_1397_),
    .B2(_1737_),
    .X(_2775_));
 sky130_fd_sc_hd__o21a_1 _6009_ (.A1(net96),
    .A2(_2775_),
    .B1(_2759_),
    .X(_2776_));
 sky130_fd_sc_hd__nor2_1 _6010_ (.A(_1086_),
    .B(net74),
    .Y(_2777_));
 sky130_fd_sc_hd__o32a_1 _6011_ (.A1(net118),
    .A2(_2776_),
    .A3(_2777_),
    .B1(net672),
    .B2(_2765_),
    .X(_0370_));
 sky130_fd_sc_hd__o2bb2a_1 _6012_ (.A1_N(_2293_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1754_),
    .X(_2778_));
 sky130_fd_sc_hd__o21a_1 _6013_ (.A1(net95),
    .A2(_2778_),
    .B1(net74),
    .X(_2779_));
 sky130_fd_sc_hd__nor2_1 _6014_ (.A(_1140_),
    .B(net74),
    .Y(_2780_));
 sky130_fd_sc_hd__o32a_1 _6015_ (.A1(net118),
    .A2(_2779_),
    .A3(_2780_),
    .B1(net779),
    .B2(_2765_),
    .X(_0371_));
 sky130_fd_sc_hd__o2bb2a_1 _6016_ (.A1_N(_2306_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1772_),
    .X(_2781_));
 sky130_fd_sc_hd__o21a_1 _6017_ (.A1(net94),
    .A2(_2781_),
    .B1(net74),
    .X(_2782_));
 sky130_fd_sc_hd__nor2_1 _6018_ (.A(_1177_),
    .B(net74),
    .Y(_2783_));
 sky130_fd_sc_hd__o32a_1 _6019_ (.A1(net118),
    .A2(_2782_),
    .A3(_2783_),
    .B1(net757),
    .B2(_2765_),
    .X(_0372_));
 sky130_fd_sc_hd__o2bb2a_1 _6020_ (.A1_N(_2319_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1790_),
    .X(_2784_));
 sky130_fd_sc_hd__o21a_1 _6021_ (.A1(net94),
    .A2(_2784_),
    .B1(net74),
    .X(_2785_));
 sky130_fd_sc_hd__nor2_1 _6022_ (.A(_1232_),
    .B(net74),
    .Y(_2786_));
 sky130_fd_sc_hd__o32a_1 _6023_ (.A1(net118),
    .A2(_2785_),
    .A3(_2786_),
    .B1(net631),
    .B2(_2765_),
    .X(_0373_));
 sky130_fd_sc_hd__o2bb2a_1 _6024_ (.A1_N(_2331_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1807_),
    .X(_2787_));
 sky130_fd_sc_hd__o21a_1 _6025_ (.A1(net94),
    .A2(_2787_),
    .B1(net74),
    .X(_2788_));
 sky130_fd_sc_hd__nor2_1 _6026_ (.A(_1281_),
    .B(net74),
    .Y(_2789_));
 sky130_fd_sc_hd__o32a_1 _6027_ (.A1(net118),
    .A2(_2788_),
    .A3(_2789_),
    .B1(net753),
    .B2(_2765_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_4 _6028_ (.A(_1968_),
    .B(_2758_),
    .X(_2790_));
 sky130_fd_sc_hd__a21oi_4 _6029_ (.A1(_2763_),
    .A2(_2790_),
    .B1(net118),
    .Y(_2791_));
 sky130_fd_sc_hd__o2bb2a_1 _6030_ (.A1_N(_2341_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1826_),
    .X(_2792_));
 sky130_fd_sc_hd__o21a_1 _6031_ (.A1(net95),
    .A2(_2792_),
    .B1(_2790_),
    .X(_2793_));
 sky130_fd_sc_hd__nor2_1 _6032_ (.A(_0863_),
    .B(_2790_),
    .Y(_2794_));
 sky130_fd_sc_hd__o32a_1 _6033_ (.A1(net118),
    .A2(_2793_),
    .A3(_2794_),
    .B1(net737),
    .B2(_2791_),
    .X(_0375_));
 sky130_fd_sc_hd__o2bb2a_1 _6034_ (.A1_N(_2354_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1843_),
    .X(_2795_));
 sky130_fd_sc_hd__o21a_1 _6035_ (.A1(net95),
    .A2(_2795_),
    .B1(_2790_),
    .X(_2796_));
 sky130_fd_sc_hd__nor2_1 _6036_ (.A(_1003_),
    .B(_2790_),
    .Y(_2797_));
 sky130_fd_sc_hd__o32a_1 _6037_ (.A1(net118),
    .A2(_2796_),
    .A3(_2797_),
    .B1(net604),
    .B2(_2791_),
    .X(_0376_));
 sky130_fd_sc_hd__o22a_1 _6038_ (.A1(net81),
    .A2(_1862_),
    .B1(_2365_),
    .B2(_2762_),
    .X(_2798_));
 sky130_fd_sc_hd__o21a_1 _6039_ (.A1(net94),
    .A2(_2798_),
    .B1(_2790_),
    .X(_2799_));
 sky130_fd_sc_hd__nor2_1 _6040_ (.A(_1053_),
    .B(_2790_),
    .Y(_2800_));
 sky130_fd_sc_hd__o32a_1 _6041_ (.A1(net118),
    .A2(_2799_),
    .A3(_2800_),
    .B1(net771),
    .B2(_2791_),
    .X(_0377_));
 sky130_fd_sc_hd__o2bb2a_1 _6042_ (.A1_N(_2372_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1879_),
    .X(_2801_));
 sky130_fd_sc_hd__o21a_1 _6043_ (.A1(net94),
    .A2(_2801_),
    .B1(_2790_),
    .X(_2802_));
 sky130_fd_sc_hd__nor2_1 _6044_ (.A(_1086_),
    .B(_2790_),
    .Y(_2803_));
 sky130_fd_sc_hd__o32a_1 _6045_ (.A1(net118),
    .A2(_2802_),
    .A3(_2803_),
    .B1(net628),
    .B2(_2791_),
    .X(_0378_));
 sky130_fd_sc_hd__o2bb2a_1 _6046_ (.A1_N(_2383_),
    .A2_N(_2761_),
    .B1(net81),
    .B2(_1898_),
    .X(_2804_));
 sky130_fd_sc_hd__o21a_1 _6047_ (.A1(net94),
    .A2(_2804_),
    .B1(_2790_),
    .X(_2805_));
 sky130_fd_sc_hd__nor2_1 _6048_ (.A(_1140_),
    .B(_2790_),
    .Y(_2806_));
 sky130_fd_sc_hd__o32a_1 _6049_ (.A1(net118),
    .A2(_2805_),
    .A3(_2806_),
    .B1(net616),
    .B2(_2791_),
    .X(_0379_));
 sky130_fd_sc_hd__o22a_1 _6050_ (.A1(net81),
    .A2(_1917_),
    .B1(_2394_),
    .B2(_2762_),
    .X(_2807_));
 sky130_fd_sc_hd__o21a_1 _6051_ (.A1(net94),
    .A2(_2807_),
    .B1(_2790_),
    .X(_2808_));
 sky130_fd_sc_hd__nor2_1 _6052_ (.A(_1177_),
    .B(_2790_),
    .Y(_2809_));
 sky130_fd_sc_hd__o32a_1 _6053_ (.A1(net118),
    .A2(_2808_),
    .A3(_2809_),
    .B1(net725),
    .B2(_2791_),
    .X(_0380_));
 sky130_fd_sc_hd__nor2_1 _6054_ (.A(net822),
    .B(_2761_),
    .Y(_2810_));
 sky130_fd_sc_hd__a31o_1 _6055_ (.A1(net91),
    .A2(_2403_),
    .A3(_2761_),
    .B1(_2810_),
    .X(_2811_));
 sky130_fd_sc_hd__nand2_1 _6056_ (.A(net81),
    .B(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__or3_1 _6057_ (.A(net94),
    .B(net81),
    .C(_1934_),
    .X(_2813_));
 sky130_fd_sc_hd__o211a_1 _6058_ (.A1(net822),
    .A2(net91),
    .B1(_2790_),
    .C1(_2813_),
    .X(_2814_));
 sky130_fd_sc_hd__a2bb2o_1 _6059_ (.A1_N(_1232_),
    .A2_N(_2790_),
    .B1(_2812_),
    .B2(_2814_),
    .X(_2815_));
 sky130_fd_sc_hd__mux2_1 _6060_ (.A0(net822),
    .A1(_2815_),
    .S(net104),
    .X(_0381_));
 sky130_fd_sc_hd__o22a_1 _6061_ (.A1(net81),
    .A2(_1953_),
    .B1(_2411_),
    .B2(_2762_),
    .X(_2816_));
 sky130_fd_sc_hd__o22a_1 _6062_ (.A1(net811),
    .A2(_2764_),
    .B1(_2816_),
    .B2(net95),
    .X(_2817_));
 sky130_fd_sc_hd__mux2_1 _6063_ (.A0(_1282_),
    .A1(_2817_),
    .S(_2790_),
    .X(_2818_));
 sky130_fd_sc_hd__mux2_1 _6064_ (.A0(net811),
    .A1(_2818_),
    .S(net105),
    .X(_0382_));
 sky130_fd_sc_hd__inv_2 _6065__2 (.A(clknet_leaf_21_wb_clk_i),
    .Y(net215));
 sky130_fd_sc_hd__inv_2 _6066__3 (.A(clknet_leaf_24_wb_clk_i),
    .Y(net216));
 sky130_fd_sc_hd__inv_2 _6067__4 (.A(clknet_leaf_24_wb_clk_i),
    .Y(net217));
 sky130_fd_sc_hd__dfxtp_1 _6068_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net516),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6069_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net423),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6070_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net393),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6071_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0044_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6072_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net442),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6073_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0046_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6074_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0047_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6075_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net419),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6076_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net219),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6077_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net539),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6078_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net724),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.R[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6079_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net579),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.R[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6080_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net625),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.R[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6081_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net541),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.R[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6082_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net611),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.R[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6083_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net587),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.R[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6084_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net609),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.R[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6085_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0058_),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6086_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net507),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.mcycles[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6087_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net467),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.mcycles[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6088_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net336),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.mcycles[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6089_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net319),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.mcycles[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6090_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net874),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6091_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net425),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6092_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net417),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6093_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net434),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6094_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net470),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6095_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0064_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6096_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net363),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6097_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net365),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6098_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net387),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6099_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net315),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6100_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net269),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6101_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net281),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6102_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net325),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6103_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net295),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6104_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net361),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6105_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net297),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6106_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net391),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6107_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(_0076_),
    .RESET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.PreserveC_r ));
 sky130_fd_sc_hd__dfxtp_1 _6108_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net356),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6109_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net344),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6110_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net327),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6111_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net381),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6112_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net338),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6113_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0082_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6114_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net317),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6115_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net352),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ));
 sky130_fd_sc_hd__dfstp_1 _6116_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net832),
    .SET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ISet[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6117_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0001_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ISet[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6118_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0002_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ISet[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6119_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0003_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ISet[3] ));
 sky130_fd_sc_hd__dfstp_1 _6120_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0020_),
    .SET_B(net176),
    .Q(\z80.normal_wr_n ));
 sky130_fd_sc_hd__dfstp_1 _6121_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0019_),
    .SET_B(net176),
    .Q(\z80.normal_rd_n ));
 sky130_fd_sc_hd__dfstp_1 _6122_ (.CLK(net214),
    .D(_0018_),
    .SET_B(net180),
    .Q(\z80.early_mreq_n ));
 sky130_fd_sc_hd__dfstp_1 _6123_ (.CLK(net215),
    .D(_0017_),
    .SET_B(net180),
    .Q(\z80.early_iorq_n ));
 sky130_fd_sc_hd__dfstp_1 _6124_ (.CLK(net216),
    .D(_0019_),
    .SET_B(net176),
    .Q(\z80.early_rd_n ));
 sky130_fd_sc_hd__dfstp_1 _6125_ (.CLK(net217),
    .D(_0020_),
    .SET_B(net176),
    .Q(\z80.early_wr_n ));
 sky130_fd_sc_hd__dfstp_1 _6126_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0018_),
    .SET_B(net180),
    .Q(\z80.normal_mreq_n ));
 sky130_fd_sc_hd__dfstp_1 _6127_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0017_),
    .SET_B(net180),
    .Q(\z80.normal_iorq_n ));
 sky130_fd_sc_hd__dfxtp_1 _6128_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net405),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6129_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net293),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6130_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net263),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6131_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net479),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6132_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net440),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6133_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0090_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6134_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net350),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6135_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net477),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6136_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net496),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6137_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net403),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6138_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net438),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6139_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net447),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6140_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net444),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6141_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0098_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6142_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_0099_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6143_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net383),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6144_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net309),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6145_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net472),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6146_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net273),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6147_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net277),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6148_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net279),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6149_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net267),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6150_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net354),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6151_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net283),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6152_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net451),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6153_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(net421),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6154_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net401),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6155_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0112_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6156_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(_0113_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6157_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net303),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6158_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0115_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6159_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net367),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6160_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net313),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6161_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net385),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6162_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net329),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6163_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0120_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6164_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0121_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6165_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(_0122_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6166_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net307),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6167_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0124_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6168_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net271),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6169_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net285),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6170_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net261),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6171_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net399),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6172_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net475),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6173_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net305),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6174_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net299),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6175_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net459),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6176_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net432),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6177_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net333),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6178_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net373),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6179_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net490),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6180_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net436),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6181_ (.CLK(clknet_leaf_51_wb_clk_i),
    .D(net428),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6182_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net411),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6183_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net494),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6184_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net323),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6185_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net492),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6186_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net257),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6187_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net259),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6188_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net311),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6189_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net359),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6190_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net377),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6191_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net289),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6192_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net510),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6193_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0150_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6194_ (.CLK(clknet_leaf_49_wb_clk_i),
    .D(net462),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6195_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0152_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6196_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(_0153_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6197_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(_0154_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6198_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(_0155_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6199_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net504),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6200_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net255),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6201_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net251),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6202_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net287),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6203_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net249),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6204_ (.CLK(clknet_leaf_14_wb_clk_i),
    .D(net389),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6205_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net265),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6206_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net409),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6207_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net342),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6208_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(net275),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6209_ (.CLK(clknet_leaf_12_wb_clk_i),
    .D(net291),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6210_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net379),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6211_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net395),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6212_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(net407),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6213_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net371),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6214_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(net369),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _6215_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net397),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6216_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0166_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6217_ (.CLK(clknet_leaf_50_wb_clk_i),
    .D(_0167_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6218_ (.CLK(clknet_leaf_47_wb_clk_i),
    .D(net449),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6219_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net430),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6220_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net321),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6221_ (.CLK(clknet_leaf_0_wb_clk_i),
    .D(net301),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6222_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net340),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _6223_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net577),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IStatus[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6224_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net413),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IStatus[2] ));
 sky130_fd_sc_hd__dfstp_1 _6225_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net704),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Ap[0] ));
 sky130_fd_sc_hd__dfstp_1 _6226_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net671),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Ap[1] ));
 sky130_fd_sc_hd__dfstp_1 _6227_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net669),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Ap[2] ));
 sky130_fd_sc_hd__dfstp_1 _6228_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net706),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Ap[3] ));
 sky130_fd_sc_hd__dfstp_1 _6229_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net694),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Ap[4] ));
 sky130_fd_sc_hd__dfstp_1 _6230_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net684),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Ap[5] ));
 sky130_fd_sc_hd__dfstp_1 _6231_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net661),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Ap[6] ));
 sky130_fd_sc_hd__dfstp_1 _6232_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net663),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.Ap[7] ));
 sky130_fd_sc_hd__dfstp_1 _6233_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net708),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Fp[0] ));
 sky130_fd_sc_hd__dfstp_1 _6234_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net746),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Fp[1] ));
 sky130_fd_sc_hd__dfstp_1 _6235_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net682),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Fp[2] ));
 sky130_fd_sc_hd__dfstp_1 _6236_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(net698),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Fp[3] ));
 sky130_fd_sc_hd__dfstp_1 _6237_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(net700),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Fp[4] ));
 sky130_fd_sc_hd__dfstp_1 _6238_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net696),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Fp[5] ));
 sky130_fd_sc_hd__dfstp_1 _6239_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net677),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Fp[6] ));
 sky130_fd_sc_hd__dfstp_1 _6240_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net686),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.Fp[7] ));
 sky130_fd_sc_hd__dfstp_1 _6241_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(_0033_),
    .SET_B(net166),
    .Q(net50));
 sky130_fd_sc_hd__dfxtp_4 _6242_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net647),
    .Q(\z80.tv80s.i_tv80_core.BusA[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6243_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net767),
    .Q(\z80.tv80s.i_tv80_core.BusA[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6244_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net659),
    .Q(\z80.tv80s.i_tv80_core.BusA[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6245_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net688),
    .Q(\z80.tv80s.i_tv80_core.BusA[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6246_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net638),
    .Q(\z80.tv80s.i_tv80_core.BusA[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6247_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(net718),
    .Q(\z80.tv80s.i_tv80_core.BusA[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6248_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net750),
    .Q(\z80.tv80s.i_tv80_core.BusA[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6249_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net534),
    .Q(\z80.tv80s.i_tv80_core.BusA[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6250_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net585),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.NMI_s ));
 sky130_fd_sc_hd__dfrtp_1 _6251_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net465),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IR[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6252_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net877),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IR[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6253_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0200_),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.IR[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6254_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0201_),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IR[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6255_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0202_),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IR[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6256_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net889),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IR[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6257_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net815),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IR[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6258_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net842),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.IR[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6259_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net528),
    .RESET_B(net177),
    .Q(net44));
 sky130_fd_sc_hd__dfrtp_1 _6260_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net530),
    .RESET_B(net177),
    .Q(net43));
 sky130_fd_sc_hd__dfrtp_1 _6261_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net546),
    .RESET_B(net177),
    .Q(net41));
 sky130_fd_sc_hd__dfrtp_1 _6262_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net566),
    .RESET_B(net177),
    .Q(net38));
 sky130_fd_sc_hd__dfrtp_1 _6263_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net562),
    .RESET_B(net177),
    .Q(net37));
 sky130_fd_sc_hd__dfrtp_1 _6264_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net573),
    .RESET_B(net177),
    .Q(net39));
 sky130_fd_sc_hd__dfrtp_1 _6265_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(net552),
    .RESET_B(net177),
    .Q(net40));
 sky130_fd_sc_hd__dfrtp_1 _6266_ (.CLK(clknet_leaf_22_wb_clk_i),
    .D(net550),
    .RESET_B(net177),
    .Q(net42));
 sky130_fd_sc_hd__dfstp_2 _6267_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0214_),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.ACC[0] ));
 sky130_fd_sc_hd__dfstp_4 _6268_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(net871),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.ACC[1] ));
 sky130_fd_sc_hd__dfstp_4 _6269_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0216_),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.ACC[2] ));
 sky130_fd_sc_hd__dfstp_4 _6270_ (.CLK(clknet_leaf_24_wb_clk_i),
    .D(_0217_),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.ACC[3] ));
 sky130_fd_sc_hd__dfstp_4 _6271_ (.CLK(clknet_leaf_33_wb_clk_i),
    .D(_0218_),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.ACC[4] ));
 sky130_fd_sc_hd__dfstp_4 _6272_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0219_),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.ACC[5] ));
 sky130_fd_sc_hd__dfstp_4 _6273_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(_0220_),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.ACC[6] ));
 sky130_fd_sc_hd__dfstp_2 _6274_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(_0221_),
    .SET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.ACC[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6275_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net548),
    .RESET_B(net166),
    .Q(net54));
 sky130_fd_sc_hd__dfrtp_1 _6276_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net591),
    .RESET_B(net169),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _6277_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net556),
    .RESET_B(net166),
    .Q(net53));
 sky130_fd_sc_hd__dfrtp_1 _6278_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net603),
    .RESET_B(net166),
    .Q(net52));
 sky130_fd_sc_hd__dfrtp_1 _6279_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net537),
    .RESET_B(net166),
    .Q(net51));
 sky130_fd_sc_hd__dfrtp_1 _6280_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net599),
    .RESET_B(net169),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _6281_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net589),
    .RESET_B(net169),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _6282_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net564),
    .RESET_B(net169),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_2 _6283_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net645),
    .RESET_B(net166),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_2 _6284_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net558),
    .RESET_B(net166),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_2 _6285_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net581),
    .RESET_B(net166),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_2 _6286_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net607),
    .RESET_B(net166),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_2 _6287_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net619),
    .RESET_B(net166),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_4 _6288_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net621),
    .RESET_B(net167),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_4 _6289_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net627),
    .RESET_B(net167),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_4 _6290_ (.CLK(clknet_leaf_36_wb_clk_i),
    .D(net665),
    .RESET_B(net167),
    .Q(net36));
 sky130_fd_sc_hd__dfstp_1 _6291_ (.CLK(clknet_leaf_23_wb_clk_i),
    .D(_0238_),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.F[0] ));
 sky130_fd_sc_hd__dfstp_4 _6292_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0239_),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.F[1] ));
 sky130_fd_sc_hd__dfstp_4 _6293_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net828),
    .SET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.F[2] ));
 sky130_fd_sc_hd__dfstp_2 _6294_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0241_),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.F[3] ));
 sky130_fd_sc_hd__dfstp_2 _6295_ (.CLK(clknet_leaf_25_wb_clk_i),
    .D(_0242_),
    .SET_B(net177),
    .Q(\z80.tv80s.i_tv80_core.F[4] ));
 sky130_fd_sc_hd__dfstp_2 _6296_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0243_),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.F[5] ));
 sky130_fd_sc_hd__dfstp_4 _6297_ (.CLK(clknet_leaf_26_wb_clk_i),
    .D(_0244_),
    .SET_B(net176),
    .Q(\z80.tv80s.i_tv80_core.F[6] ));
 sky130_fd_sc_hd__dfstp_2 _6298_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net835),
    .SET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.F[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6299_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net575),
    .Q(\z80.tv80s.i_tv80_core.IncDecZ ));
 sky130_fd_sc_hd__dfrtp_1 _6300_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net331),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.Z16_r ));
 sky130_fd_sc_hd__dfrtp_4 _6301_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(net853),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6302_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net851),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6303_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net844),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6304_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(_0251_),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6305_ (.CLK(clknet_leaf_19_wb_clk_i),
    .D(_0252_),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Save_ALU_r ));
 sky130_fd_sc_hd__dfrtp_1 _6306_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net346),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.BTR_r ));
 sky130_fd_sc_hd__dfrtp_1 _6307_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(_0254_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6308_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net512),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6309_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net526),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6310_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net532),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6311_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0258_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6312_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net799),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.Arith16_r ));
 sky130_fd_sc_hd__dfxtp_4 _6313_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net885),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ));
 sky130_fd_sc_hd__dfxtp_4 _6314_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net651),
    .Q(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6315_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(_0262_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.XY_Ind ));
 sky130_fd_sc_hd__dfrtp_1 _6316_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net667),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.XY_State[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6317_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net786),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.XY_State[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6318_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net881),
    .Q(\z80.tv80s.i_tv80_core.RegAddrC[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6319_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net791),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6320_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net797),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6321_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net803),
    .RESET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6322_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net826),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6323_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net824),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6324_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(net810),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6325_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net819),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6326_ (.CLK(clknet_leaf_29_wb_clk_i),
    .D(net808),
    .RESET_B(net175),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6327_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net740),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[8] ));
 sky130_fd_sc_hd__dfrtp_1 _6328_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net601),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6329_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net776),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6330_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net742),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[11] ));
 sky130_fd_sc_hd__dfrtp_4 _6331_ (.CLK(clknet_leaf_46_wb_clk_i),
    .D(net730),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[12] ));
 sky130_fd_sc_hd__dfrtp_4 _6332_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net795),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[13] ));
 sky130_fd_sc_hd__dfrtp_4 _6333_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net748),
    .RESET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[14] ));
 sky130_fd_sc_hd__dfrtp_2 _6334_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net744),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.TmpAddr[15] ));
 sky130_fd_sc_hd__dfrtp_2 _6335_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net554),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.Alternate ));
 sky130_fd_sc_hd__dfxtp_4 _6336_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net714),
    .Q(\z80.tv80s.i_tv80_core.BusB[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6337_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net593),
    .Q(\z80.tv80s.i_tv80_core.BusB[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6338_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net583),
    .Q(\z80.tv80s.i_tv80_core.BusB[2] ));
 sky130_fd_sc_hd__dfxtp_4 _6339_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net657),
    .Q(\z80.tv80s.i_tv80_core.BusB[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6340_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net692),
    .Q(\z80.tv80s.i_tv80_core.BusB[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6341_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net675),
    .Q(\z80.tv80s.i_tv80_core.BusB[5] ));
 sky130_fd_sc_hd__dfxtp_4 _6342_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net643),
    .Q(\z80.tv80s.i_tv80_core.BusB[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6343_ (.CLK(clknet_leaf_32_wb_clk_i),
    .D(net679),
    .Q(\z80.tv80s.i_tv80_core.BusB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6344_ (.CLK(clknet_leaf_11_wb_clk_i),
    .D(_0291_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6345_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(_0292_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6346_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net241),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6347_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net233),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6348_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net229),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6349_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net223),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6350_ (.CLK(clknet_leaf_6_wb_clk_i),
    .D(net221),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6351_ (.CLK(clknet_leaf_7_wb_clk_i),
    .D(net225),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6352_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(_0299_),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6353_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net231),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6354_ (.CLK(clknet_leaf_48_wb_clk_i),
    .D(net237),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6355_ (.CLK(clknet_leaf_44_wb_clk_i),
    .D(net227),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6356_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net235),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6357_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net245),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6358_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net247),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6359_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net243),
    .Q(\z80.tv80s.i_tv80_core.RegBusA_r[15] ));
 sky130_fd_sc_hd__dfrtp_1 _6360_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net615),
    .RESET_B(net166),
    .Q(\z80.tv80s.i_tv80_core.I[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6361_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net595),
    .RESET_B(net167),
    .Q(\z80.tv80s.i_tv80_core.I[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6362_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net634),
    .RESET_B(net167),
    .Q(\z80.tv80s.i_tv80_core.I[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6363_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net702),
    .RESET_B(net167),
    .Q(\z80.tv80s.i_tv80_core.I[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6364_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net720),
    .RESET_B(net166),
    .Q(\z80.tv80s.i_tv80_core.I[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6365_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net752),
    .RESET_B(net167),
    .Q(\z80.tv80s.i_tv80_core.I[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6366_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net623),
    .RESET_B(net166),
    .Q(\z80.tv80s.i_tv80_core.I[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6367_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net778),
    .RESET_B(net166),
    .Q(\z80.tv80s.i_tv80_core.I[7] ));
 sky130_fd_sc_hd__dfrtp_1 _6368_ (.CLK(clknet_leaf_34_wb_clk_i),
    .D(net375),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.R[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6369_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net253),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6370_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net239),
    .Q(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6371_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net710),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.PC[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6372_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net690),
    .RESET_B(net170),
    .Q(\z80.tv80s.i_tv80_core.PC[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6373_ (.CLK(clknet_leaf_30_wb_clk_i),
    .D(net597),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.PC[2] ));
 sky130_fd_sc_hd__dfrtp_1 _6374_ (.CLK(clknet_leaf_31_wb_clk_i),
    .D(net613),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.PC[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6375_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net712),
    .RESET_B(net169),
    .Q(\z80.tv80s.i_tv80_core.PC[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6376_ (.CLK(clknet_leaf_35_wb_clk_i),
    .D(net770),
    .RESET_B(net166),
    .Q(\z80.tv80s.i_tv80_core.PC[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6377_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net722),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.PC[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6378_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net756),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.PC[7] ));
 sky130_fd_sc_hd__dfrtp_4 _6379_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net813),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.PC[8] ));
 sky130_fd_sc_hd__dfrtp_4 _6380_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net821),
    .RESET_B(net167),
    .Q(\z80.tv80s.i_tv80_core.PC[9] ));
 sky130_fd_sc_hd__dfrtp_4 _6381_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net801),
    .RESET_B(net167),
    .Q(\z80.tv80s.i_tv80_core.PC[10] ));
 sky130_fd_sc_hd__dfrtp_4 _6382_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net793),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.PC[11] ));
 sky130_fd_sc_hd__dfrtp_2 _6383_ (.CLK(clknet_leaf_39_wb_clk_i),
    .D(net765),
    .RESET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.PC[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6384_ (.CLK(clknet_leaf_37_wb_clk_i),
    .D(net728),
    .RESET_B(net167),
    .Q(\z80.tv80s.i_tv80_core.PC[13] ));
 sky130_fd_sc_hd__dfrtp_4 _6385_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net736),
    .RESET_B(net167),
    .Q(\z80.tv80s.i_tv80_core.PC[14] ));
 sky130_fd_sc_hd__dfrtp_4 _6386_ (.CLK(clknet_leaf_38_wb_clk_i),
    .D(net760),
    .RESET_B(net166),
    .Q(\z80.tv80s.i_tv80_core.PC[15] ));
 sky130_fd_sc_hd__dfstp_1 _6387_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0334_),
    .SET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ));
 sky130_fd_sc_hd__dfrtp_1 _6388_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net868),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6389_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net857),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6390_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net784),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6391_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net763),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6392_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net846),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6393_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net839),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6394_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net774),
    .RESET_B(net179),
    .Q(\z80.tv80s.i_tv80_core.Halt_FF ));
 sky130_fd_sc_hd__dfrtp_1 _6395_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0029_),
    .RESET_B(net172),
    .Q(_0034_));
 sky130_fd_sc_hd__dfrtp_1 _6396_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(_0030_),
    .RESET_B(net173),
    .Q(_0035_));
 sky130_fd_sc_hd__dfrtp_1 _6397_ (.CLK(clknet_leaf_13_wb_clk_i),
    .D(net544),
    .RESET_B(net174),
    .Q(_0036_));
 sky130_fd_sc_hd__dfrtp_1 _6398_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(net734),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ));
 sky130_fd_sc_hd__dfrtp_1 _6399_ (.CLK(clknet_leaf_15_wb_clk_i),
    .D(net732),
    .RESET_B(net174),
    .Q(\z80.tv80s.i_tv80_core.No_BTR ));
 sky130_fd_sc_hd__dfrtp_1 _6400_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net649),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.IntCycle ));
 sky130_fd_sc_hd__dfrtp_1 _6401_ (.CLK(clknet_leaf_17_wb_clk_i),
    .D(_0022_),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ));
 sky130_fd_sc_hd__dfrtp_4 _6402_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0342_),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.BusAck ));
 sky130_fd_sc_hd__dfrtp_1 _6403_ (.CLK(clknet_leaf_18_wb_clk_i),
    .D(net10),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.Oldnmi_n ));
 sky130_fd_sc_hd__dfrtp_1 _6404_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(_0025_),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.INT_s ));
 sky130_fd_sc_hd__dfrtp_4 _6405_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net485),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.NMICycle ));
 sky130_fd_sc_hd__dfrtp_1 _6406_ (.CLK(clknet_leaf_21_wb_clk_i),
    .D(_0023_),
    .RESET_B(net180),
    .Q(\z80.tv80s.i_tv80_core.BusReq_s ));
 sky130_fd_sc_hd__dfxtp_1 _6407_ (.CLK(clknet_leaf_4_wb_clk_i),
    .D(net520),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _6408_ (.CLK(clknet_leaf_5_wb_clk_i),
    .D(net457),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _6409_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(net348),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _6410_ (.CLK(clknet_leaf_2_wb_clk_i),
    .D(_0347_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _6411_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0348_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _6412_ (.CLK(clknet_leaf_52_wb_clk_i),
    .D(_0349_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _6413_ (.CLK(clknet_leaf_1_wb_clk_i),
    .D(net454),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _6414_ (.CLK(clknet_leaf_3_wb_clk_i),
    .D(_0351_),
    .Q(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ));
 sky130_fd_sc_hd__dfstp_2 _6415_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(net636),
    .SET_B(net175),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_4 _6416_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0352_),
    .RESET_B(net175),
    .Q(\z80.tv80s.di_reg[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6417_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0353_),
    .RESET_B(net175),
    .Q(\z80.tv80s.di_reg[1] ));
 sky130_fd_sc_hd__dfrtp_4 _6418_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0354_),
    .RESET_B(net175),
    .Q(\z80.tv80s.di_reg[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6419_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0355_),
    .RESET_B(net175),
    .Q(\z80.tv80s.di_reg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _6420_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(_0356_),
    .RESET_B(net175),
    .Q(\z80.tv80s.di_reg[4] ));
 sky130_fd_sc_hd__dfrtp_4 _6421_ (.CLK(clknet_leaf_28_wb_clk_i),
    .D(_0357_),
    .RESET_B(net175),
    .Q(\z80.tv80s.di_reg[5] ));
 sky130_fd_sc_hd__dfrtp_4 _6422_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0358_),
    .RESET_B(net175),
    .Q(\z80.tv80s.di_reg[6] ));
 sky130_fd_sc_hd__dfrtp_4 _6423_ (.CLK(clknet_leaf_27_wb_clk_i),
    .D(_0359_),
    .RESET_B(net175),
    .Q(\z80.tv80s.di_reg[7] ));
 sky130_fd_sc_hd__dfstp_1 _6424_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net524),
    .SET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.ts[0] ));
 sky130_fd_sc_hd__dfrtp_4 _6425_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(_0361_),
    .RESET_B(net173),
    .Q(\z80.tv80s.i_tv80_core.ts[1] ));
 sky130_fd_sc_hd__dfrtp_1 _6426_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0362_),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.ts[2] ));
 sky130_fd_sc_hd__dfrtp_4 _6427_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(_0363_),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.ts[3] ));
 sky130_fd_sc_hd__dfrtp_1 _6428_ (.CLK(clknet_leaf_9_wb_clk_i),
    .D(net569),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.ts[4] ));
 sky130_fd_sc_hd__dfrtp_1 _6429_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net487),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.ts[5] ));
 sky130_fd_sc_hd__dfrtp_1 _6430_ (.CLK(clknet_leaf_10_wb_clk_i),
    .D(net482),
    .RESET_B(net172),
    .Q(\z80.tv80s.i_tv80_core.ts[6] ));
 sky130_fd_sc_hd__dfrtp_1 _6431_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net789),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.IntE ));
 sky130_fd_sc_hd__dfrtp_1 _6432_ (.CLK(clknet_leaf_16_wb_clk_i),
    .D(net806),
    .RESET_B(net178),
    .Q(\z80.tv80s.i_tv80_core.IntE_FF2 ));
 sky130_fd_sc_hd__dfstp_1 _6433_ (.CLK(clknet_leaf_8_wb_clk_i),
    .D(net716),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[0] ));
 sky130_fd_sc_hd__dfstp_1 _6434_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net655),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[1] ));
 sky130_fd_sc_hd__dfstp_1 _6435_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net653),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[2] ));
 sky130_fd_sc_hd__dfstp_1 _6436_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net673),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[3] ));
 sky130_fd_sc_hd__dfstp_1 _6437_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net780),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[4] ));
 sky130_fd_sc_hd__dfstp_2 _6438_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net758),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[5] ));
 sky130_fd_sc_hd__dfstp_1 _6439_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net632),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.SP[6] ));
 sky130_fd_sc_hd__dfstp_1 _6440_ (.CLK(clknet_leaf_42_wb_clk_i),
    .D(net754),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[7] ));
 sky130_fd_sc_hd__dfstp_1 _6441_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(net738),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[8] ));
 sky130_fd_sc_hd__dfstp_1 _6442_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net605),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[9] ));
 sky130_fd_sc_hd__dfstp_1 _6443_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net772),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[10] ));
 sky130_fd_sc_hd__dfstp_1 _6444_ (.CLK(clknet_leaf_45_wb_clk_i),
    .D(net629),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[11] ));
 sky130_fd_sc_hd__dfstp_1 _6445_ (.CLK(clknet_leaf_43_wb_clk_i),
    .D(net617),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[12] ));
 sky130_fd_sc_hd__dfstp_1 _6446_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(net726),
    .SET_B(net171),
    .Q(\z80.tv80s.i_tv80_core.SP[13] ));
 sky130_fd_sc_hd__dfstp_2 _6447_ (.CLK(clknet_leaf_40_wb_clk_i),
    .D(_0381_),
    .SET_B(net168),
    .Q(\z80.tv80s.i_tv80_core.SP[14] ));
 sky130_fd_sc_hd__dfstp_1 _6448_ (.CLK(clknet_leaf_41_wb_clk_i),
    .D(_0382_),
    .SET_B(net181),
    .Q(\z80.tv80s.i_tv80_core.SP[15] ));
 sky130_fd_sc_hd__buf_1 _6481_ (.A(net22),
    .X(net15));
 sky130_fd_sc_hd__buf_1 _6482_ (.A(net22),
    .X(net16));
 sky130_fd_sc_hd__buf_1 _6483_ (.A(net22),
    .X(net17));
 sky130_fd_sc_hd__buf_1 _6484_ (.A(net22),
    .X(net18));
 sky130_fd_sc_hd__buf_1 _6485_ (.A(net22),
    .X(net19));
 sky130_fd_sc_hd__buf_1 _6486_ (.A(net22),
    .X(net20));
 sky130_fd_sc_hd__buf_1 _6487_ (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__conb_1 ci2406_z80_182 (.LO(net182));
 sky130_fd_sc_hd__conb_1 ci2406_z80_183 (.LO(net183));
 sky130_fd_sc_hd__conb_1 ci2406_z80_184 (.LO(net184));
 sky130_fd_sc_hd__conb_1 ci2406_z80_185 (.LO(net185));
 sky130_fd_sc_hd__conb_1 ci2406_z80_186 (.LO(net186));
 sky130_fd_sc_hd__conb_1 ci2406_z80_187 (.LO(net187));
 sky130_fd_sc_hd__conb_1 ci2406_z80_188 (.LO(net188));
 sky130_fd_sc_hd__conb_1 ci2406_z80_189 (.LO(net189));
 sky130_fd_sc_hd__conb_1 ci2406_z80_190 (.LO(net190));
 sky130_fd_sc_hd__conb_1 ci2406_z80_191 (.LO(net191));
 sky130_fd_sc_hd__conb_1 ci2406_z80_192 (.LO(net192));
 sky130_fd_sc_hd__conb_1 ci2406_z80_193 (.LO(net193));
 sky130_fd_sc_hd__conb_1 ci2406_z80_194 (.LO(net194));
 sky130_fd_sc_hd__conb_1 ci2406_z80_195 (.LO(net195));
 sky130_fd_sc_hd__conb_1 ci2406_z80_196 (.LO(net196));
 sky130_fd_sc_hd__conb_1 ci2406_z80_197 (.LO(net197));
 sky130_fd_sc_hd__conb_1 ci2406_z80_198 (.LO(net198));
 sky130_fd_sc_hd__conb_1 ci2406_z80_199 (.LO(net199));
 sky130_fd_sc_hd__conb_1 ci2406_z80_200 (.LO(net200));
 sky130_fd_sc_hd__conb_1 ci2406_z80_201 (.LO(net201));
 sky130_fd_sc_hd__conb_1 ci2406_z80_202 (.LO(net202));
 sky130_fd_sc_hd__conb_1 ci2406_z80_203 (.LO(net203));
 sky130_fd_sc_hd__conb_1 ci2406_z80_204 (.LO(net204));
 sky130_fd_sc_hd__conb_1 ci2406_z80_205 (.LO(net205));
 sky130_fd_sc_hd__conb_1 ci2406_z80_206 (.LO(net206));
 sky130_fd_sc_hd__conb_1 ci2406_z80_207 (.LO(net207));
 sky130_fd_sc_hd__conb_1 ci2406_z80_208 (.LO(net208));
 sky130_fd_sc_hd__conb_1 ci2406_z80_209 (.LO(net209));
 sky130_fd_sc_hd__conb_1 ci2406_z80_210 (.HI(net210));
 sky130_fd_sc_hd__conb_1 ci2406_z80_211 (.HI(net211));
 sky130_fd_sc_hd__conb_1 ci2406_z80_212 (.HI(net212));
 sky130_fd_sc_hd__conb_1 ci2406_z80_213 (.HI(net213));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_10_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_11_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_12_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_13_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_14_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_15_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_16_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_17_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_18_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_19_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_1_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_21_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_22_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_23_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_24_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_25_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_26_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_27_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.A(clknet_2_3__leaf_wb_clk_i),
    .X(clknet_leaf_28_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_29_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_2_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_30_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_31_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_32_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_33_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_34_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_35_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_36_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_37_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_38_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.A(clknet_2_2__leaf_wb_clk_i),
    .X(clknet_leaf_39_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_3_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_40_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_41_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_42_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_43_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_44_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_45_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_46_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_47_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_48_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_49_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_4_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_50_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_51_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_52_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_5_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.A(clknet_2_0__leaf_wb_clk_i),
    .X(clknet_leaf_6_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_7_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_8_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.A(clknet_2_1__leaf_wb_clk_i),
    .X(clknet_leaf_9_wb_clk_i));
 sky130_fd_sc_hd__buf_2 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(_3031_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(_2941_),
    .X(net103));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(net110),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(net110),
    .X(net107));
 sky130_fd_sc_hd__buf_6 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout110 (.A(net23),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_8 fanout111 (.A(net112),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(_2827_),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_8 fanout113 (.A(_2826_),
    .X(net113));
 sky130_fd_sc_hd__buf_8 fanout114 (.A(_2822_),
    .X(net114));
 sky130_fd_sc_hd__buf_8 fanout115 (.A(net116),
    .X(net115));
 sky130_fd_sc_hd__buf_8 fanout116 (.A(\z80.tv80s.i_tv80_core.ts[3] ),
    .X(net116));
 sky130_fd_sc_hd__buf_8 fanout117 (.A(net639),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_8 fanout118 (.A(\z80.tv80s.i_tv80_core.BusAck ),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(net829),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(\z80.tv80s.i_tv80_core.BusAck ),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_8 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net829),
    .X(net122));
 sky130_fd_sc_hd__buf_4 fanout123 (.A(net804),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_8 fanout124 (.A(net126),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__buf_6 fanout126 (.A(net867),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net128),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net130),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_8 fanout129 (.A(net130),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net883),
    .X(net131));
 sky130_fd_sc_hd__buf_6 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__buf_6 fanout133 (.A(net880),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_8 fanout135 (.A(net884),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_8 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 fanout137 (.A(net850),
    .X(net137));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net872),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_8 fanout139 (.A(\z80.tv80s.i_tv80_core.IR[5] ),
    .X(net139));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(net888),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net145),
    .X(net142));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(net731),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_8 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_8 fanout147 (.A(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(net147));
 sky130_fd_sc_hd__buf_4 fanout148 (.A(net150),
    .X(net148));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(\z80.tv80s.i_tv80_core.IR[3] ),
    .X(net150));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(net153),
    .X(net151));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 fanout153 (.A(net891),
    .X(net153));
 sky130_fd_sc_hd__buf_6 fanout154 (.A(net876),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net876),
    .X(net155));
 sky130_fd_sc_hd__buf_6 fanout156 (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(net887),
    .X(net158));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(net831),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net831),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_8 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__buf_6 fanout164 (.A(net873),
    .X(net164));
 sky130_fd_sc_hd__buf_8 fanout165 (.A(net847),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_8 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__buf_4 fanout168 (.A(net181),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(net181),
    .X(net169));
 sky130_fd_sc_hd__buf_4 fanout170 (.A(net181),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_8 fanout171 (.A(net181),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_6 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_6 fanout174 (.A(net181),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_8 fanout175 (.A(net178),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_4 fanout178 (.A(net181),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_8 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__buf_4 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_8 fanout181 (.A(net14),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_8 fanout55 (.A(_1648_),
    .X(net55));
 sky130_fd_sc_hd__buf_8 fanout56 (.A(_0574_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_8 fanout57 (.A(_0494_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 fanout59 (.A(_2559_),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_4 fanout61 (.A(_1666_),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(_1664_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_8 fanout64 (.A(_2643_),
    .X(net64));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(_2326_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_8 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_4 fanout67 (.A(_1653_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_8 fanout68 (.A(_0874_),
    .X(net68));
 sky130_fd_sc_hd__buf_4 fanout69 (.A(_0819_),
    .X(net69));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(_1565_),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_8 fanout71 (.A(_0817_),
    .X(net71));
 sky130_fd_sc_hd__buf_6 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(_0816_),
    .X(net73));
 sky130_fd_sc_hd__buf_4 fanout74 (.A(_2759_),
    .X(net74));
 sky130_fd_sc_hd__buf_4 fanout75 (.A(_0814_),
    .X(net75));
 sky130_fd_sc_hd__buf_4 fanout76 (.A(_0814_),
    .X(net76));
 sky130_fd_sc_hd__buf_4 fanout77 (.A(_0814_),
    .X(net77));
 sky130_fd_sc_hd__buf_4 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_4 fanout79 (.A(_1399_),
    .X(net79));
 sky130_fd_sc_hd__buf_4 fanout80 (.A(_1398_),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_4 fanout81 (.A(_1397_),
    .X(net81));
 sky130_fd_sc_hd__buf_4 fanout82 (.A(_0783_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 fanout83 (.A(_0783_),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(_0781_),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_8 fanout85 (.A(_0780_),
    .X(net85));
 sky130_fd_sc_hd__buf_4 fanout86 (.A(_0780_),
    .X(net86));
 sky130_fd_sc_hd__buf_4 fanout88 (.A(_2884_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_8 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(_1668_),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_8 fanout91 (.A(net93),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_8 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_8 fanout93 (.A(_0602_),
    .X(net93));
 sky130_fd_sc_hd__buf_4 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_4 fanout95 (.A(_0601_),
    .X(net95));
 sky130_fd_sc_hd__buf_4 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_8 fanout97 (.A(_0601_),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(_0497_),
    .X(net98));
 sky130_fd_sc_hd__buf_6 fanout99 (.A(net101),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[2] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0302_),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0083_),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\z80.tv80s.i_tv80_core.mcycles[5] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0016_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][5] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0170_),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][0] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0141_),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][3] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0071_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][2] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[4] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0079_),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][2] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0119_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\z80.tv80s.i_tv80_core.Z16_r ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0247_),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][1] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0134_),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t1 ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\z80.tv80s.i_tv80_core.mcycles[4] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_0015_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0295_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][4] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_0081_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][7] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_0172_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][0] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_0157_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][1] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_0078_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\z80.tv80s.i_tv80_core.BTR_r ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_0253_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[9] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][2] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_0346_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][6] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_0091_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][7] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_0084_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][6] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_0107_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][0] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_0077_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0300_),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][6] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][5] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0146_),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][5] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0073_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][5] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0065_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][6] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0066_),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][7] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[3] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0116_),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][7] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0164_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][6] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_0163_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][2] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0135_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\z80.tv80s.i_tv80_core.R[7] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0315_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][6] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0294_),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0147_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][3] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0160_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][3] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0080_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][7] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0100_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][1] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0118_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][7] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[12] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0067_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[5] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0010_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][7] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0075_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][2] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0043_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][4] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0161_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][0] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0303_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0165_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][3] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0128_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][2] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0111_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][1] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0094_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][0] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0085_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][5] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[10] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_0162_),
    .X(net407));
 sky130_fd_sc_hd__buf_1 hold191 (.A(net900),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0012_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][6] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0139_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\z80.tv80s.i_tv80_core.IStatus[2] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0005_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][6] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][6] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][1] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0049_),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0301_),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0061_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][7] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0048_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][1] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0110_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][1] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0042_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][0] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0060_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][1] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[1] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][5] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_0138_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][4] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_0169_),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][0] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_0133_),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][2] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_0062_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][4] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_0137_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0317_),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][2] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_0095_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][4] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_0089_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][4] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_0045_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][4] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_0097_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][5] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][3] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[2] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0096_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][3] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0168_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][0] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0109_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][4] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][6] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(_0350_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][1] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][1] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0293_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0345_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][7] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_0132_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][6] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][2] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(_0151_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][5] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\z80.tv80s.i_tv80_core.IR[0] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0198_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\z80.tv80s.i_tv80_core.mcycles[2] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[15] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0014_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][5] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][3] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_0063_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][1] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_0102_),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\z80.tv80s.i_tv80_core.ISet[3] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][4] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0129_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][7] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0306_),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0092_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][3] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0088_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][5] ),
    .X(net480));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold264 (.A(\z80.tv80s.i_tv80_core.ts[5] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_0366_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][4] ),
    .X(net483));
 sky130_fd_sc_hd__buf_1 hold267 (.A(\z80.tv80s.i_tv80_core.NMI_s ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0343_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\z80.tv80s.i_tv80_core.ts[4] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[13] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0365_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][3] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][3] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_0136_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][1] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(_0142_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[3][7] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_0140_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][0] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_0093_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0304_),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][3] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][3] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[7][5] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][7] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][4] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][3] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][7] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(_0156_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][2] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\z80.tv80s.i_tv80_core.mcycles[1] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[14] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0013_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][5] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[2][0] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_0149_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[1] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_0255_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][5] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[6][4] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[3][0] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_0041_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[6] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0305_),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][4] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][3] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][0] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_0344_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\z80.tv80s.i_tv80_core.PreserveC_r ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[2][7] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\z80.tv80s.i_tv80_core.ts[6] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_0360_),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[2] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(_0256_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[4] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(net44),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(_0206_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(net43),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_0207_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[3] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(_0257_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\z80.tv80s.i_tv80_core.BusA[7] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(_0196_),
    .X(net534));
 sky130_fd_sc_hd__buf_1 hold318 (.A(net897),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(net51),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0009_),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0226_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[2] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0050_),
    .X(net539));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold323 (.A(\z80.tv80s.i_tv80_core.R[3] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0054_),
    .X(net541));
 sky130_fd_sc_hd__buf_1 hold325 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[4] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0593_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(_0031_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(net41),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(_0208_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[2] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(net54),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_0222_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(net42),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_0213_),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(net40),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(_0212_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\z80.tv80s.i_tv80_core.Alternate ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(_0282_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(net53),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(_0224_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0007_),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(net29),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(_0231_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[8] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[0] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(net37),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(_0210_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(net27),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(_0229_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(net38),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(_0209_),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\z80.tv80s.i_tv80_core.RegAddrA_r[0] ),
    .X(net252));
 sky130_fd_sc_hd__buf_2 hold350 (.A(net899),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(_2754_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0364_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[1] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_2543_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(net39),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_0211_),
    .X(net573));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold357 (.A(\z80.tv80s.i_tv80_core.IncDecZ ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0246_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\z80.tv80s.i_tv80_core.IStatus[1] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0316_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0004_),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_2 hold361 (.A(\z80.tv80s.i_tv80_core.R[1] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_0052_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(net30),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_0232_),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 hold365 (.A(\z80.tv80s.i_tv80_core.BusB[2] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0285_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\z80.tv80s.i_tv80_core.Oldnmi_n ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_0197_),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 hold369 (.A(\z80.tv80s.i_tv80_core.R[5] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[1] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0056_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(net26),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0228_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(net24),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0223_),
    .X(net591));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold375 (.A(\z80.tv80s.i_tv80_core.BusB[1] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0284_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\z80.tv80s.i_tv80_core.I[1] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_0308_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\z80.tv80s.i_tv80_core.PC[2] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0006_),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0320_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(net25),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_0227_),
    .X(net599));
 sky130_fd_sc_hd__buf_1 hold383 (.A(\z80.tv80s.i_tv80_core.TmpAddr[9] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_0275_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(net52),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0225_),
    .X(net603));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold387 (.A(\z80.tv80s.i_tv80_core.SP[9] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0376_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(net31),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][2] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_0233_),
    .X(net607));
 sky130_fd_sc_hd__buf_1 hold391 (.A(\z80.tv80s.i_tv80_core.R[6] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0057_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\z80.tv80s.i_tv80_core.R[4] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_0055_),
    .X(net611));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold395 (.A(\z80.tv80s.i_tv80_core.PC[3] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0321_),
    .X(net613));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold397 (.A(\z80.tv80s.i_tv80_core.I[0] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0307_),
    .X(net615));
 sky130_fd_sc_hd__buf_1 hold399 (.A(\z80.tv80s.i_tv80_core.SP[12] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0297_),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0143_),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0379_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(net32),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0234_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(net33),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0235_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\z80.tv80s.i_tv80_core.I[6] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_0313_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\z80.tv80s.i_tv80_core.R[2] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0053_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(net35),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][3] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0236_),
    .X(net627));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold411 (.A(\z80.tv80s.i_tv80_core.SP[11] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0378_),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_2 hold413 (.A(net898),
    .X(net630));
 sky130_fd_sc_hd__buf_1 hold414 (.A(\z80.tv80s.i_tv80_core.SP[6] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(_0373_),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\z80.tv80s.i_tv80_core.I[2] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(_0309_),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\z80.tv80s.i_tv80_core.ts[0] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(_0032_),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0144_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\z80.tv80s.i_tv80_core.BusA[4] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(_0193_),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_2 hold422 (.A(\z80.tv80s.i_tv80_core.ts[2] ),
    .X(net639));
 sky130_fd_sc_hd__buf_1 hold423 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[2] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0587_),
    .X(net641));
 sky130_fd_sc_hd__buf_1 hold425 (.A(\z80.tv80s.i_tv80_core.BusB[6] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0289_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(net28),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0230_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\z80.tv80s.i_tv80_core.BusA[0] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][2] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0189_),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_2 hold431 (.A(\z80.tv80s.i_tv80_core.IntCycle ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0341_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[1] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_0261_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\z80.tv80s.i_tv80_core.SP[2] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_0369_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\z80.tv80s.i_tv80_core.SP[1] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0368_),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_2 hold439 (.A(\z80.tv80s.i_tv80_core.BusB[3] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0127_),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0286_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\z80.tv80s.i_tv80_core.BusA[2] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0191_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\z80.tv80s.i_tv80_core.Ap[6] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0179_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\z80.tv80s.i_tv80_core.Ap[7] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_0180_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(net36),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0237_),
    .X(net665));
 sky130_fd_sc_hd__buf_1 hold449 (.A(\z80.tv80s.i_tv80_core.XY_State[0] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][2] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_0263_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\z80.tv80s.i_tv80_core.Ap[2] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_0175_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\z80.tv80s.i_tv80_core.Ap[1] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_0174_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\z80.tv80s.i_tv80_core.SP[3] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_0370_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\z80.tv80s.i_tv80_core.BusB[5] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0288_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\z80.tv80s.i_tv80_core.Fp[6] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0087_),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0187_),
    .X(net677));
 sky130_fd_sc_hd__buf_1 hold461 (.A(\z80.tv80s.i_tv80_core.BusB[7] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_0290_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\z80.tv80s.i_tv80_core.ISet[1] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\z80.tv80s.i_tv80_core.Fp[2] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(_0183_),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\z80.tv80s.i_tv80_core.Ap[5] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(_0178_),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\z80.tv80s.i_tv80_core.Fp[7] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(_0188_),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[6] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\z80.tv80s.i_tv80_core.BusA[3] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(_0192_),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\z80.tv80s.i_tv80_core.PC[1] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(_0319_),
    .X(net690));
 sky130_fd_sc_hd__buf_1 hold474 (.A(\z80.tv80s.i_tv80_core.BusB[4] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(_0287_),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\z80.tv80s.i_tv80_core.Ap[4] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(_0177_),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\z80.tv80s.i_tv80_core.Fp[5] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(_0186_),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0011_),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\z80.tv80s.i_tv80_core.Fp[3] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(_0184_),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\z80.tv80s.i_tv80_core.Fp[4] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(_0185_),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\z80.tv80s.i_tv80_core.I[3] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(_0310_),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\z80.tv80s.i_tv80_core.Ap[0] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(_0173_),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\z80.tv80s.i_tv80_core.Ap[3] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(_0176_),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][5] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\z80.tv80s.i_tv80_core.Fp[0] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(_0181_),
    .X(net708));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold492 (.A(\z80.tv80s.i_tv80_core.PC[0] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(_0318_),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\z80.tv80s.i_tv80_core.PC[4] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(_0322_),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_2 hold496 (.A(\z80.tv80s.i_tv80_core.BusB[0] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(_0283_),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\z80.tv80s.i_tv80_core.SP[0] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(_0367_),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[5] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0106_),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\z80.tv80s.i_tv80_core.BusA[5] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(_0194_),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\z80.tv80s.i_tv80_core.I[4] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(_0311_),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\z80.tv80s.i_tv80_core.PC[6] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(_0324_),
    .X(net722));
 sky130_fd_sc_hd__buf_1 hold506 (.A(\z80.tv80s.i_tv80_core.R[0] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(_0051_),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\z80.tv80s.i_tv80_core.SP[13] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(_0380_),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][1] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\z80.tv80s.i_tv80_core.PC[13] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(_0331_),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\z80.tv80s.i_tv80_core.TmpAddr[12] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(_0278_),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\z80.tv80s.i_tv80_core.IR[4] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(_0028_),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\z80.tv80s.i_tv80_core.Auto_Wait_t2 ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(_0021_),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\z80.tv80s.i_tv80_core.PC[14] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(_0332_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0069_),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\z80.tv80s.i_tv80_core.SP[8] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(_0375_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\z80.tv80s.i_tv80_core.TmpAddr[8] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(_0274_),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\z80.tv80s.i_tv80_core.TmpAddr[11] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(_0277_),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\z80.tv80s.i_tv80_core.TmpAddr[15] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(_0281_),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\z80.tv80s.i_tv80_core.Fp[1] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(_0182_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][0] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\z80.tv80s.i_tv80_core.TmpAddr[14] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(_0280_),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\z80.tv80s.i_tv80_core.BusA[6] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(_0195_),
    .X(net750));
 sky130_fd_sc_hd__buf_1 hold534 (.A(\z80.tv80s.i_tv80_core.I[5] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(_0312_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\z80.tv80s.i_tv80_core.SP[7] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(_0374_),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\z80.tv80s.i_tv80_core.PC[7] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(_0325_),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0125_),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\z80.tv80s.i_tv80_core.SP[5] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(_0372_),
    .X(net758));
 sky130_fd_sc_hd__buf_1 hold542 (.A(\z80.tv80s.i_tv80_core.PC[15] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(_0333_),
    .X(net760));
 sky130_fd_sc_hd__buf_1 hold544 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[3] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(_2746_),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0338_),
    .X(net763));
 sky130_fd_sc_hd__buf_1 hold547 (.A(\z80.tv80s.i_tv80_core.PC[12] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_0330_),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\z80.tv80s.i_tv80_core.BusA[1] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][2] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_0190_),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_2 hold551 (.A(\z80.tv80s.i_tv80_core.ts[1] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\z80.tv80s.i_tv80_core.PC[5] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(_0323_),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\z80.tv80s.i_tv80_core.SP[10] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(_0377_),
    .X(net772));
 sky130_fd_sc_hd__buf_1 hold556 (.A(\z80.tv80s.i_tv80_core.Halt_FF ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(_0024_),
    .X(net774));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold558 (.A(\z80.tv80s.i_tv80_core.TmpAddr[10] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(_0276_),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0103_),
    .X(net273));
 sky130_fd_sc_hd__buf_1 hold560 (.A(\z80.tv80s.i_tv80_core.I[7] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(_0314_),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\z80.tv80s.i_tv80_core.SP[4] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(_0371_),
    .X(net780));
 sky130_fd_sc_hd__buf_1 hold564 (.A(_0034_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(_2737_),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_2745_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(_0337_),
    .X(net784));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold568 (.A(\z80.tv80s.i_tv80_core.XY_State[1] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(_0264_),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][1] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\z80.tv80s.i_tv80_core.IntE ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(_0744_),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0026_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\z80.tv80s.i_tv80_core.TmpAddr[0] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0266_),
    .X(net791));
 sky130_fd_sc_hd__buf_1 hold575 (.A(\z80.tv80s.i_tv80_core.PC[11] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0329_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\z80.tv80s.i_tv80_core.TmpAddr[13] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0279_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\z80.tv80s.i_tv80_core.TmpAddr[1] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0158_),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0267_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\z80.tv80s.i_tv80_core.Arith16_r ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0259_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\z80.tv80s.i_tv80_core.PC[10] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0328_),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\z80.tv80s.i_tv80_core.TmpAddr[2] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0268_),
    .X(net803));
 sky130_fd_sc_hd__buf_1 hold587 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[6] ),
    .X(net804));
 sky130_fd_sc_hd__buf_1 hold588 (.A(\z80.tv80s.i_tv80_core.IntE_FF2 ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(_0027_),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][3] ),
    .X(net276));
 sky130_fd_sc_hd__buf_1 hold590 (.A(\z80.tv80s.i_tv80_core.TmpAddr[7] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(_0273_),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\z80.tv80s.i_tv80_core.TmpAddr[5] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(_0271_),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\z80.tv80s.i_tv80_core.SP[15] ),
    .X(net811));
 sky130_fd_sc_hd__buf_1 hold595 (.A(\z80.tv80s.i_tv80_core.PC[8] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0326_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\z80.tv80s.i_tv80_core.IR[6] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0204_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\z80.tv80s.i_tv80_core.F[3] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0296_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0104_),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\z80.tv80s.i_tv80_core.F[5] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\z80.tv80s.i_tv80_core.TmpAddr[6] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0272_),
    .X(net819));
 sky130_fd_sc_hd__buf_1 hold603 (.A(\z80.tv80s.i_tv80_core.PC[9] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0327_),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\z80.tv80s.i_tv80_core.SP[14] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\z80.tv80s.i_tv80_core.TmpAddr[4] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(_0270_),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\z80.tv80s.i_tv80_core.TmpAddr[3] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(_0269_),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][4] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\z80.tv80s.i_tv80_core.F[2] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(_0240_),
    .X(net828));
 sky130_fd_sc_hd__buf_1 hold612 (.A(\z80.tv80s.i_tv80_core.BusAck ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\z80.tv80s.i_tv80_core.F[4] ),
    .X(net830));
 sky130_fd_sc_hd__buf_1 hold614 (.A(\z80.tv80s.i_tv80_core.ISet[0] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(_0000_),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[3] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\z80.tv80s.i_tv80_core.F[7] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_0245_),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\z80.tv80s.i_tv80_core.ACC[7] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0105_),
    .X(net279));
 sky130_fd_sc_hd__buf_1 hold620 (.A(_0036_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(_2750_),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0340_),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_2 hold623 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net840));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold624 (.A(\z80.tv80s.i_tv80_core.IR[7] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(_0205_),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[2] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(_0250_),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_2 hold628 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[5] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(_0339_),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][2] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\z80.tv80s.i_tv80_core.RegAddrC[2] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\z80.tv80s.di_reg[2] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\z80.tv80s.di_reg[1] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[1] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_0249_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\z80.tv80s.i_tv80_core.ALU_Op_r[0] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_0248_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\z80.tv80s.di_reg[0] ),
    .X(net854));
 sky130_fd_sc_hd__buf_1 hold638 (.A(_0035_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(_2744_),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0070_),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_0336_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\z80.tv80s.di_reg[3] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\z80.tv80s.di_reg[5] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\z80.tv80s.di_reg[6] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\z80.tv80s.di_reg[7] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\z80.tv80s.di_reg[4] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\z80.tv80s.i_tv80_core.ACC[4] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\z80.tv80s.i_tv80_core.ACC[6] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\z80.tv80s.i_tv80_core.ACC[2] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\z80.tv80s.i_tv80_core.ACC[0] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][7] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[1] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(_0335_),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\z80.tv80s.i_tv80_core.F[6] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\z80.tv80s.i_tv80_core.ACC[1] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_0215_),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\z80.tv80s.i_tv80_core.F[0] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\z80.tv80s.i_tv80_core.RegAddrC[1] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(_0059_),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\z80.tv80s.i_tv80_core.ACC[5] ),
    .X(net875));
 sky130_fd_sc_hd__buf_1 hold659 (.A(\z80.tv80s.i_tv80_core.IR[1] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0108_),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_0199_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\z80.tv80s.i_tv80_core.XY_Ind ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\z80.tv80s.i_tv80_core.ACC[3] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\z80.tv80s.i_tv80_core.RegAddrC[0] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_0265_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\z80.tv80s.i_tv80_core.No_BTR ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\z80.tv80s.i_tv80_core.i_mcode.MCycle[0] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\z80.tv80s.i_tv80_core.RegAddrB_r[0] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_0260_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\z80.tv80s.i_tv80_core.F[1] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][1] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\z80.tv80s.i_tv80_core.ISet[2] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\z80.tv80s.i_tv80_core.IR[5] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_0203_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\z80.tv80s.i_tv80_core.NMICycle ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\z80.tv80s.i_tv80_core.IR[2] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\z80.tv80s.i_tv80_core.ts[6] ),
    .X(net894));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold678 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net895));
 sky130_fd_sc_hd__buf_1 hold679 (.A(\z80.tv80s.i_tv80_core.Save_ALU_r ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0126_),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[4] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\z80.tv80s.i_tv80_core.Read_To_Reg_r[0] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\z80.tv80s.i_tv80_core.BusReq_s ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[7] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\z80.tv80s.i_tv80_core.Pre_XY_F_M[3] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[7] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0008_),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][7] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0148_),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[7][2] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0159_),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[6][1] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0086_),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][4] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0072_),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][6] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0298_),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0074_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][6] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0131_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[0][6] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0171_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[1][5] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0114_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[1][5] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0130_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][6] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\z80.tv80s.i_tv80_core.RegBusA_r[11] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0123_),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[5][0] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0101_),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[4][4] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0145_),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsL[0][0] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0117_),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[5][0] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0068_),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\z80.tv80s.i_tv80_core.i_reg.RegsH[4][6] ),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(custom_settings[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(io_in[30]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(io_in[31]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(io_in[35]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 input13 (.A(io_in[4]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(rst_n),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(io_in[22]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(io_in[23]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(io_in[24]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(io_in[25]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(io_in[26]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(io_in[27]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(io_in[28]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(io_in[29]),
    .X(net9));
 sky130_fd_sc_hd__buf_4 max_cap58 (.A(_1671_),
    .X(net58));
 sky130_fd_sc_hd__buf_2 max_cap87 (.A(_2974_),
    .X(net87));
 sky130_fd_sc_hd__buf_12 output15 (.A(net15),
    .X(io_oeb[22]));
 sky130_fd_sc_hd__buf_12 output16 (.A(net16),
    .X(io_oeb[23]));
 sky130_fd_sc_hd__buf_12 output17 (.A(net17),
    .X(io_oeb[24]));
 sky130_fd_sc_hd__buf_12 output18 (.A(net18),
    .X(io_oeb[25]));
 sky130_fd_sc_hd__buf_12 output19 (.A(net19),
    .X(io_oeb[26]));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(io_oeb[27]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(io_oeb[28]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(io_oeb[29]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net110),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(io_out[10]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(io_out[11]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(io_out[12]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(io_out[13]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(io_out[14]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(io_out[15]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(io_out[16]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(io_out[17]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(io_out[18]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(io_out[19]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(io_out[20]));
 sky130_fd_sc_hd__buf_12 output36 (.A(net36),
    .X(io_out[21]));
 sky130_fd_sc_hd__buf_12 output37 (.A(net37),
    .X(io_out[22]));
 sky130_fd_sc_hd__buf_12 output38 (.A(net38),
    .X(io_out[23]));
 sky130_fd_sc_hd__buf_12 output39 (.A(net39),
    .X(io_out[24]));
 sky130_fd_sc_hd__buf_12 output40 (.A(net40),
    .X(io_out[25]));
 sky130_fd_sc_hd__buf_12 output41 (.A(net41),
    .X(io_out[26]));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(io_out[27]));
 sky130_fd_sc_hd__buf_12 output43 (.A(net43),
    .X(io_out[28]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net44),
    .X(io_out[29]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(io_out[32]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(io_out[33]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net48),
    .X(io_out[34]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net49),
    .X(io_out[3]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(io_out[5]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(io_out[6]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net52),
    .X(io_out[7]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net53),
    .X(io_out[8]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net54),
    .X(io_out[9]));
 assign io_oeb[0] = net182;
 assign io_oeb[10] = net191;
 assign io_oeb[11] = net192;
 assign io_oeb[12] = net193;
 assign io_oeb[13] = net194;
 assign io_oeb[14] = net195;
 assign io_oeb[15] = net196;
 assign io_oeb[16] = net197;
 assign io_oeb[17] = net198;
 assign io_oeb[18] = net199;
 assign io_oeb[19] = net200;
 assign io_oeb[1] = net183;
 assign io_oeb[20] = net201;
 assign io_oeb[21] = net202;
 assign io_oeb[2] = net184;
 assign io_oeb[30] = net211;
 assign io_oeb[31] = net212;
 assign io_oeb[32] = net203;
 assign io_oeb[33] = net204;
 assign io_oeb[34] = net205;
 assign io_oeb[35] = net213;
 assign io_oeb[3] = net185;
 assign io_oeb[4] = net210;
 assign io_oeb[5] = net186;
 assign io_oeb[6] = net187;
 assign io_oeb[7] = net188;
 assign io_oeb[8] = net189;
 assign io_oeb[9] = net190;
 assign io_out[30] = net207;
 assign io_out[31] = net208;
 assign io_out[35] = net209;
 assign io_out[4] = net206;
endmodule

