magic
tech sky130B
magscale 1 2
timestamp 1717259628
<< viali >>
rect 5273 32453 5307 32487
rect 10425 32453 10459 32487
rect 2881 32385 2915 32419
rect 4077 32385 4111 32419
rect 6193 32385 6227 32419
rect 8677 32385 8711 32419
rect 11161 32385 11195 32419
rect 13921 32385 13955 32419
rect 15301 32385 15335 32419
rect 17785 32385 17819 32419
rect 18337 32385 18371 32419
rect 19257 32385 19291 32419
rect 21833 32385 21867 32419
rect 23305 32385 23339 32419
rect 24409 32385 24443 32419
rect 26985 32385 27019 32419
rect 29561 32385 29595 32419
rect 32137 32385 32171 32419
rect 1593 32317 1627 32351
rect 2605 32317 2639 32351
rect 6745 32317 6779 32351
rect 8401 32317 8435 32351
rect 9873 32317 9907 32351
rect 11897 32317 11931 32351
rect 13461 32317 13495 32351
rect 14473 32317 14507 32351
rect 15577 32317 15611 32351
rect 17509 32317 17543 32351
rect 19717 32317 19751 32351
rect 21281 32317 21315 32351
rect 22293 32317 22327 32351
rect 24869 32317 24903 32351
rect 26433 32317 26467 32351
rect 27445 32317 27479 32351
rect 29009 32317 29043 32351
rect 30021 32317 30055 32351
rect 31585 32317 31619 32351
rect 32597 32317 32631 32351
rect 9229 32249 9263 32283
rect 25881 32249 25915 32283
rect 2145 32181 2179 32215
rect 4721 32181 4755 32215
rect 7297 32181 7331 32215
rect 12449 32181 12483 32215
rect 15025 32181 15059 32215
rect 16865 32181 16899 32215
rect 20729 32181 20763 32215
rect 23949 32181 23983 32215
rect 28457 32181 28491 32215
rect 31033 32181 31067 32215
rect 2973 31977 3007 32011
rect 3893 31909 3927 31943
rect 9321 31909 9355 31943
rect 9505 31909 9539 31943
rect 3525 31841 3559 31875
rect 4813 31841 4847 31875
rect 6561 31841 6595 31875
rect 7849 31841 7883 31875
rect 10609 31841 10643 31875
rect 12081 31841 12115 31875
rect 13001 31841 13035 31875
rect 15485 31841 15519 31875
rect 18521 31841 18555 31875
rect 20545 31841 20579 31875
rect 22845 31841 22879 31875
rect 25237 31841 25271 31875
rect 28181 31841 28215 31875
rect 30113 31841 30147 31875
rect 32045 31841 32079 31875
rect 1593 31773 1627 31807
rect 2605 31773 2639 31807
rect 4261 31773 4295 31807
rect 4353 31773 4387 31807
rect 7113 31773 7147 31807
rect 7481 31773 7515 31807
rect 9781 31773 9815 31807
rect 10885 31773 10919 31807
rect 12357 31773 12391 31807
rect 12541 31773 12575 31807
rect 14473 31773 14507 31807
rect 15025 31773 15059 31807
rect 15209 31773 15243 31807
rect 16865 31773 16899 31807
rect 19073 31773 19107 31807
rect 19993 31773 20027 31807
rect 20913 31773 20947 31807
rect 22293 31773 22327 31807
rect 23121 31773 23155 31807
rect 23305 31773 23339 31807
rect 23857 31773 23891 31807
rect 24685 31773 24719 31807
rect 26157 31773 26191 31807
rect 27629 31773 27663 31807
rect 29561 31773 29595 31807
rect 32321 31773 32355 31807
rect 32505 31773 32539 31807
rect 33057 31773 33091 31807
rect 9045 31705 9079 31739
rect 17233 31705 17267 31739
rect 26525 31705 26559 31739
rect 3801 31637 3835 31671
rect 18153 31637 18187 31671
rect 21281 31637 21315 31671
rect 25697 31637 25731 31671
rect 27169 31637 27203 31671
rect 28549 31637 28583 31671
rect 31217 31637 31251 31671
rect 1777 31433 1811 31467
rect 4261 31433 4295 31467
rect 8309 31433 8343 31467
rect 13185 31433 13219 31467
rect 15025 31433 15059 31467
rect 21005 31433 21039 31467
rect 26709 31433 26743 31467
rect 2780 31365 2814 31399
rect 6193 31365 6227 31399
rect 7972 31365 8006 31399
rect 31861 31365 31895 31399
rect 2513 31297 2547 31331
rect 5385 31297 5419 31331
rect 8217 31297 8251 31331
rect 9985 31297 10019 31331
rect 10241 31297 10275 31331
rect 12837 31297 12871 31331
rect 14309 31297 14343 31331
rect 14565 31297 14599 31331
rect 16149 31297 16183 31331
rect 16405 31297 16439 31331
rect 17805 31297 17839 31331
rect 18061 31297 18095 31331
rect 20013 31297 20047 31331
rect 20269 31297 20303 31331
rect 23222 31297 23256 31331
rect 23489 31297 23523 31331
rect 24797 31297 24831 31331
rect 25053 31297 25087 31331
rect 25329 31297 25363 31331
rect 25596 31297 25630 31331
rect 28109 31297 28143 31331
rect 28365 31297 28399 31331
rect 28549 31297 28583 31331
rect 29101 31297 29135 31331
rect 31042 31297 31076 31331
rect 31309 31297 31343 31331
rect 32229 31297 32263 31331
rect 2421 31229 2455 31263
rect 5641 31229 5675 31263
rect 8769 31229 8803 31263
rect 11345 31229 11379 31263
rect 13093 31229 13127 31263
rect 18705 31229 18739 31263
rect 20361 31229 20395 31263
rect 20821 31229 20855 31263
rect 21649 31229 21683 31263
rect 32505 31229 32539 31263
rect 3893 31161 3927 31195
rect 5917 31161 5951 31195
rect 8401 31161 8435 31195
rect 20545 31161 20579 31195
rect 31493 31161 31527 31195
rect 5733 31093 5767 31127
rect 6837 31093 6871 31127
rect 8861 31093 8895 31127
rect 10701 31093 10735 31127
rect 11713 31093 11747 31127
rect 16681 31093 16715 31127
rect 18153 31093 18187 31127
rect 18889 31093 18923 31127
rect 22109 31093 22143 31127
rect 23673 31093 23707 31127
rect 26985 31093 27019 31127
rect 29929 31093 29963 31127
rect 31401 31093 31435 31127
rect 12357 30889 12391 30923
rect 17141 30889 17175 30923
rect 21925 30889 21959 30923
rect 25881 30889 25915 30923
rect 33149 30889 33183 30923
rect 15577 30821 15611 30855
rect 21741 30821 21775 30855
rect 26065 30821 26099 30855
rect 5549 30753 5583 30787
rect 7481 30753 7515 30787
rect 9873 30753 9907 30787
rect 12265 30753 12299 30787
rect 16129 30753 16163 30787
rect 16589 30753 16623 30787
rect 17693 30753 17727 30787
rect 19257 30753 19291 30787
rect 20361 30753 20395 30787
rect 22477 30753 22511 30787
rect 22845 30753 22879 30787
rect 23673 30753 23707 30787
rect 27445 30753 27479 30787
rect 28365 30753 28399 30787
rect 30941 30753 30975 30787
rect 1777 30685 1811 30719
rect 5089 30685 5123 30719
rect 5816 30685 5850 30719
rect 8033 30685 8067 30719
rect 9413 30685 9447 30719
rect 11998 30685 12032 30719
rect 12909 30685 12943 30719
rect 13369 30685 13403 30719
rect 13921 30685 13955 30719
rect 14197 30685 14231 30719
rect 14565 30685 14599 30719
rect 17233 30685 17267 30719
rect 19901 30685 19935 30719
rect 23489 30685 23523 30719
rect 25789 30685 25823 30719
rect 27905 30685 27939 30719
rect 28089 30685 28123 30719
rect 32413 30685 32447 30719
rect 32505 30685 32539 30719
rect 2044 30617 2078 30651
rect 4721 30617 4755 30651
rect 20628 30617 20662 30651
rect 24593 30617 24627 30651
rect 26341 30617 26375 30651
rect 30674 30617 30708 30651
rect 32146 30617 32180 30651
rect 3157 30549 3191 30583
rect 6929 30549 6963 30583
rect 9137 30549 9171 30583
rect 10885 30549 10919 30583
rect 24225 30549 24259 30583
rect 29561 30549 29595 30583
rect 31033 30549 31067 30583
rect 6837 30345 6871 30379
rect 11345 30345 11379 30379
rect 13093 30345 13127 30379
rect 13737 30345 13771 30379
rect 14473 30345 14507 30379
rect 16313 30345 16347 30379
rect 18153 30345 18187 30379
rect 21189 30345 21223 30379
rect 22477 30345 22511 30379
rect 26525 30345 26559 30379
rect 2329 30277 2363 30311
rect 3065 30277 3099 30311
rect 4537 30277 4571 30311
rect 6377 30277 6411 30311
rect 9137 30277 9171 30311
rect 11897 30277 11931 30311
rect 24777 30277 24811 30311
rect 32382 30277 32416 30311
rect 2697 30209 2731 30243
rect 4261 30209 4295 30243
rect 5549 30209 5583 30243
rect 7021 30209 7055 30243
rect 9689 30209 9723 30243
rect 10425 30209 10459 30243
rect 10793 30209 10827 30243
rect 12449 30209 12483 30243
rect 12633 30209 12667 30243
rect 13461 30209 13495 30243
rect 18613 30209 18647 30243
rect 18981 30209 19015 30243
rect 21649 30209 21683 30243
rect 25421 30209 25455 30243
rect 29009 30209 29043 30243
rect 29745 30209 29779 30243
rect 30665 30209 30699 30243
rect 7665 30141 7699 30175
rect 8309 30141 8343 30175
rect 14289 30141 14323 30175
rect 14933 30141 14967 30175
rect 15853 30141 15887 30175
rect 22109 30141 22143 30175
rect 23397 30141 23431 30175
rect 23581 30141 23615 30175
rect 24225 30141 24259 30175
rect 24869 30141 24903 30175
rect 25973 30141 26007 30175
rect 26985 30141 27019 30175
rect 27445 30141 27479 30175
rect 28549 30141 28583 30175
rect 29193 30141 29227 30175
rect 30941 30141 30975 30175
rect 32137 30141 32171 30175
rect 6745 30073 6779 30107
rect 7757 30073 7791 30107
rect 9873 30073 9907 30107
rect 13001 30073 13035 30107
rect 14565 30073 14599 30107
rect 16221 30073 16255 30107
rect 18337 30073 18371 30107
rect 21373 30073 21407 30107
rect 22937 30073 22971 30107
rect 23121 30073 23155 30107
rect 23949 30073 23983 30107
rect 27169 30073 27203 30107
rect 15301 30005 15335 30039
rect 15761 30005 15795 30039
rect 24041 30005 24075 30039
rect 30113 30005 30147 30039
rect 33517 30005 33551 30039
rect 6009 29801 6043 29835
rect 7205 29801 7239 29835
rect 10333 29801 10367 29835
rect 11253 29801 11287 29835
rect 26249 29801 26283 29835
rect 27905 29801 27939 29835
rect 6193 29733 6227 29767
rect 7297 29733 7331 29767
rect 10517 29733 10551 29767
rect 29561 29733 29595 29767
rect 29745 29733 29779 29767
rect 4537 29665 4571 29699
rect 5273 29665 5307 29699
rect 6469 29665 6503 29699
rect 6653 29665 6687 29699
rect 7849 29665 7883 29699
rect 10793 29665 10827 29699
rect 11161 29665 11195 29699
rect 11805 29665 11839 29699
rect 24869 29665 24903 29699
rect 25421 29665 25455 29699
rect 30573 29665 30607 29699
rect 2697 29597 2731 29631
rect 2973 29597 3007 29631
rect 5089 29597 5123 29631
rect 23581 29597 23615 29631
rect 24225 29597 24259 29631
rect 25605 29597 25639 29631
rect 26893 29597 26927 29631
rect 27353 29597 27387 29631
rect 28089 29597 28123 29631
rect 30297 29597 30331 29631
rect 31677 29597 31711 29631
rect 2329 29529 2363 29563
rect 28641 29529 28675 29563
rect 30021 29529 30055 29563
rect 31922 29529 31956 29563
rect 3525 29461 3559 29495
rect 5917 29461 5951 29495
rect 26157 29461 26191 29495
rect 33057 29461 33091 29495
rect 7665 29257 7699 29291
rect 26065 29257 26099 29291
rect 29009 29257 29043 29291
rect 30297 29189 30331 29223
rect 2697 29121 2731 29155
rect 2881 29121 2915 29155
rect 4445 29121 4479 29155
rect 7021 29121 7055 29155
rect 27261 29121 27295 29155
rect 28457 29121 28491 29155
rect 29193 29121 29227 29155
rect 31953 29121 31987 29155
rect 32393 29121 32427 29155
rect 2145 29053 2179 29087
rect 3341 29053 3375 29087
rect 4813 29053 4847 29087
rect 25513 29053 25547 29087
rect 26801 29053 26835 29087
rect 27905 29053 27939 29087
rect 31493 29053 31527 29087
rect 32137 29053 32171 29087
rect 26157 28917 26191 28951
rect 28181 28917 28215 28951
rect 33517 28917 33551 28951
rect 29377 28713 29411 28747
rect 4445 28577 4479 28611
rect 5917 28577 5951 28611
rect 6009 28577 6043 28611
rect 25881 28577 25915 28611
rect 27353 28577 27387 28611
rect 30849 28577 30883 28611
rect 32505 28577 32539 28611
rect 2697 28509 2731 28543
rect 2973 28509 3007 28543
rect 3893 28509 3927 28543
rect 6653 28509 6687 28543
rect 7297 28509 7331 28543
rect 9597 28509 9631 28543
rect 26433 28509 26467 28543
rect 26525 28509 26559 28543
rect 27997 28509 28031 28543
rect 28733 28509 28767 28543
rect 30573 28509 30607 28543
rect 31861 28509 31895 28543
rect 32229 28509 32263 28543
rect 2329 28441 2363 28475
rect 28641 28441 28675 28475
rect 3525 28373 3559 28407
rect 5273 28373 5307 28407
rect 6745 28373 6779 28407
rect 8953 28373 8987 28407
rect 27169 28373 27203 28407
rect 27905 28373 27939 28407
rect 29929 28373 29963 28407
rect 5089 28169 5123 28203
rect 27537 28169 27571 28203
rect 29653 28169 29687 28203
rect 33517 28169 33551 28203
rect 3617 28101 3651 28135
rect 32382 28101 32416 28135
rect 2605 28033 2639 28067
rect 4169 28033 4203 28067
rect 5733 28033 5767 28067
rect 28825 28033 28859 28067
rect 30389 28033 30423 28067
rect 31953 28033 31987 28067
rect 1593 27965 1627 27999
rect 4445 27965 4479 27999
rect 26985 27965 27019 27999
rect 27445 27965 27479 27999
rect 28181 27965 28215 27999
rect 29101 27965 29135 27999
rect 31493 27965 31527 27999
rect 32137 27965 32171 27999
rect 27353 27897 27387 27931
rect 28273 27897 28307 27931
rect 4997 27829 5031 27863
rect 26801 27829 26835 27863
rect 29837 27829 29871 27863
rect 3157 27625 3191 27659
rect 3801 27625 3835 27659
rect 4537 27625 4571 27659
rect 5273 27625 5307 27659
rect 27905 27625 27939 27659
rect 30205 27625 30239 27659
rect 27169 27557 27203 27591
rect 27721 27557 27755 27591
rect 4445 27489 4479 27523
rect 5089 27489 5123 27523
rect 27353 27489 27387 27523
rect 28549 27489 28583 27523
rect 31861 27489 31895 27523
rect 32505 27489 32539 27523
rect 1777 27421 1811 27455
rect 5825 27421 5859 27455
rect 28733 27421 28767 27455
rect 29285 27421 29319 27455
rect 29561 27421 29595 27455
rect 30665 27421 30699 27455
rect 32229 27421 32263 27455
rect 2044 27353 2078 27387
rect 26893 27353 26927 27387
rect 27445 27353 27479 27387
rect 27997 27285 28031 27319
rect 4261 27081 4295 27115
rect 10425 27081 10459 27115
rect 28273 27081 28307 27115
rect 28365 27081 28399 27115
rect 29745 27081 29779 27115
rect 30481 27081 30515 27115
rect 5549 27013 5583 27047
rect 31769 27013 31803 27047
rect 2697 26945 2731 26979
rect 3148 26945 3182 26979
rect 4353 26945 4387 26979
rect 6469 26945 6503 26979
rect 7113 26945 7147 26979
rect 28917 26945 28951 26979
rect 29929 26945 29963 26979
rect 30757 26945 30791 26979
rect 32321 26945 32355 26979
rect 2421 26877 2455 26911
rect 2881 26877 2915 26911
rect 5089 26877 5123 26911
rect 11069 26877 11103 26911
rect 27537 26877 27571 26911
rect 27813 26877 27847 26911
rect 29101 26877 29135 26911
rect 33333 26877 33367 26911
rect 5181 26809 5215 26843
rect 28089 26809 28123 26843
rect 4997 26741 5031 26775
rect 3801 26537 3835 26571
rect 5273 26537 5307 26571
rect 29377 26537 29411 26571
rect 4537 26469 4571 26503
rect 5457 26469 5491 26503
rect 29193 26469 29227 26503
rect 30021 26469 30055 26503
rect 2329 26401 2363 26435
rect 4445 26401 4479 26435
rect 5733 26401 5767 26435
rect 28089 26401 28123 26435
rect 2605 26333 2639 26367
rect 2973 26333 3007 26367
rect 5089 26333 5123 26367
rect 18153 26333 18187 26367
rect 30205 26333 30239 26367
rect 30941 26333 30975 26367
rect 31677 26333 31711 26367
rect 28457 26265 28491 26299
rect 28917 26265 28951 26299
rect 29653 26265 29687 26299
rect 31922 26265 31956 26299
rect 3525 26197 3559 26231
rect 17601 26197 17635 26231
rect 28825 26197 28859 26231
rect 30113 26197 30147 26231
rect 30849 26197 30883 26231
rect 31585 26197 31619 26231
rect 33057 26197 33091 26231
rect 3249 25993 3283 26027
rect 3985 25993 4019 26027
rect 17417 25993 17451 26027
rect 29837 25993 29871 26027
rect 32597 25925 32631 25959
rect 1777 25857 1811 25891
rect 2044 25857 2078 25891
rect 30481 25857 30515 25891
rect 32229 25857 32263 25891
rect 3801 25789 3835 25823
rect 4537 25789 4571 25823
rect 4721 25789 4755 25823
rect 5181 25789 5215 25823
rect 16773 25789 16807 25823
rect 28825 25789 28859 25823
rect 29193 25789 29227 25823
rect 29285 25789 29319 25823
rect 30573 25789 30607 25823
rect 31217 25789 31251 25823
rect 31309 25789 31343 25823
rect 3157 25721 3191 25755
rect 4813 25721 4847 25755
rect 29653 25721 29687 25755
rect 29745 25653 29779 25687
rect 31953 25653 31987 25687
rect 1777 25449 1811 25483
rect 3801 25449 3835 25483
rect 29377 25449 29411 25483
rect 33057 25449 33091 25483
rect 30113 25313 30147 25347
rect 31677 25313 31711 25347
rect 3157 25245 3191 25279
rect 3617 25245 3651 25279
rect 4445 25245 4479 25279
rect 28733 25245 28767 25279
rect 31585 25245 31619 25279
rect 31933 25245 31967 25279
rect 2912 25177 2946 25211
rect 3249 25177 3283 25211
rect 3433 25177 3467 25211
rect 30665 25177 30699 25211
rect 31217 24905 31251 24939
rect 4077 24837 4111 24871
rect 32597 24837 32631 24871
rect 2605 24769 2639 24803
rect 13205 24769 13239 24803
rect 15577 24769 15611 24803
rect 15945 24769 15979 24803
rect 16221 24769 16255 24803
rect 30573 24769 30607 24803
rect 32229 24769 32263 24803
rect 1593 24701 1627 24735
rect 2973 24701 3007 24735
rect 13461 24701 13495 24735
rect 15117 24701 15151 24735
rect 31861 24701 31895 24735
rect 3801 24633 3835 24667
rect 15301 24633 15335 24667
rect 3525 24565 3559 24599
rect 3617 24565 3651 24599
rect 12081 24565 12115 24599
rect 15761 24565 15795 24599
rect 31309 24565 31343 24599
rect 2973 24361 3007 24395
rect 3801 24361 3835 24395
rect 15761 24361 15795 24395
rect 30757 24361 30791 24395
rect 31217 24293 31251 24327
rect 2421 24225 2455 24259
rect 3617 24225 3651 24259
rect 30849 24225 30883 24259
rect 2697 24157 2731 24191
rect 4353 24157 4387 24191
rect 31401 24157 31435 24191
rect 32321 24157 32355 24191
rect 33333 24089 33367 24123
rect 31309 24021 31343 24055
rect 32045 24021 32079 24055
rect 4261 23817 4295 23851
rect 8309 23817 8343 23851
rect 27629 23817 27663 23851
rect 31217 23817 31251 23851
rect 33517 23817 33551 23851
rect 3148 23749 3182 23783
rect 32382 23749 32416 23783
rect 2605 23681 2639 23715
rect 9597 23681 9631 23715
rect 28641 23681 28675 23715
rect 30389 23681 30423 23715
rect 32137 23681 32171 23715
rect 1593 23613 1627 23647
rect 2881 23613 2915 23647
rect 26985 23613 27019 23647
rect 30665 23613 30699 23647
rect 31953 23613 31987 23647
rect 28457 23545 28491 23579
rect 9873 23477 9907 23511
rect 31309 23477 31343 23511
rect 2973 23273 3007 23307
rect 4445 23273 4479 23307
rect 18153 23273 18187 23307
rect 27353 23273 27387 23307
rect 30757 23273 30791 23307
rect 4629 23205 4663 23239
rect 31217 23205 31251 23239
rect 2421 23137 2455 23171
rect 3525 23137 3559 23171
rect 30849 23137 30883 23171
rect 31953 23137 31987 23171
rect 32505 23137 32539 23171
rect 2697 23069 2731 23103
rect 3801 23069 3835 23103
rect 17509 23069 17543 23103
rect 32229 23069 32263 23103
rect 4997 23001 5031 23035
rect 26065 23001 26099 23035
rect 4537 22933 4571 22967
rect 25881 22933 25915 22967
rect 31309 22933 31343 22967
rect 31401 22933 31435 22967
rect 28549 22729 28583 22763
rect 1777 22593 1811 22627
rect 2044 22593 2078 22627
rect 31953 22593 31987 22627
rect 32229 22593 32263 22627
rect 3341 22525 3375 22559
rect 3985 22525 4019 22559
rect 4537 22525 4571 22559
rect 4721 22525 4755 22559
rect 5181 22525 5215 22559
rect 27905 22525 27939 22559
rect 31493 22525 31527 22559
rect 32505 22525 32539 22559
rect 3157 22457 3191 22491
rect 4813 22457 4847 22491
rect 3893 22389 3927 22423
rect 3801 22185 3835 22219
rect 31585 22185 31619 22219
rect 33057 22185 33091 22219
rect 1777 22049 1811 22083
rect 4353 22049 4387 22083
rect 31033 22049 31067 22083
rect 2044 21981 2078 22015
rect 31677 21981 31711 22015
rect 31922 21913 31956 21947
rect 3157 21845 3191 21879
rect 30665 21573 30699 21607
rect 30757 21573 30791 21607
rect 2605 21505 2639 21539
rect 32321 21505 32355 21539
rect 1593 21437 1627 21471
rect 2973 21437 3007 21471
rect 3617 21437 3651 21471
rect 4169 21437 4203 21471
rect 4813 21437 4847 21471
rect 31953 21437 31987 21471
rect 33333 21437 33367 21471
rect 4445 21369 4479 21403
rect 31125 21369 31159 21403
rect 3525 21301 3559 21335
rect 4353 21301 4387 21335
rect 31217 21301 31251 21335
rect 31309 21301 31343 21335
rect 3157 21097 3191 21131
rect 3801 21097 3835 21131
rect 25421 21097 25455 21131
rect 33057 21097 33091 21131
rect 1777 20961 1811 20995
rect 5273 20961 5307 20995
rect 31033 20961 31067 20995
rect 4445 20893 4479 20927
rect 24777 20893 24811 20927
rect 31677 20893 31711 20927
rect 2044 20825 2078 20859
rect 7021 20825 7055 20859
rect 31922 20825 31956 20859
rect 7389 20757 7423 20791
rect 31585 20757 31619 20791
rect 2329 20485 2363 20519
rect 32597 20485 32631 20519
rect 2697 20417 2731 20451
rect 2973 20417 3007 20451
rect 31953 20417 31987 20451
rect 32229 20417 32263 20451
rect 3617 20349 3651 20383
rect 31401 20349 31435 20383
rect 17233 20009 17267 20043
rect 31401 20009 31435 20043
rect 31861 19941 31895 19975
rect 1777 19873 1811 19907
rect 31585 19873 31619 19907
rect 4445 19805 4479 19839
rect 18613 19805 18647 19839
rect 32229 19805 32263 19839
rect 2044 19737 2078 19771
rect 18346 19737 18380 19771
rect 32597 19737 32631 19771
rect 3157 19669 3191 19703
rect 3801 19669 3835 19703
rect 18981 19669 19015 19703
rect 32045 19669 32079 19703
rect 4353 19465 4387 19499
rect 26801 19465 26835 19499
rect 27169 19465 27203 19499
rect 1593 19329 1627 19363
rect 2605 19329 2639 19363
rect 3525 19329 3559 19363
rect 25428 19329 25462 19363
rect 25677 19329 25711 19363
rect 32321 19329 32355 19363
rect 33333 19329 33367 19363
rect 2881 19261 2915 19295
rect 3709 19261 3743 19295
rect 4813 19261 4847 19295
rect 31309 19261 31343 19295
rect 4445 19193 4479 19227
rect 4261 19125 4295 19159
rect 31953 19125 31987 19159
rect 2881 18921 2915 18955
rect 4537 18921 4571 18955
rect 18061 18921 18095 18955
rect 1961 18853 1995 18887
rect 5365 18853 5399 18887
rect 18245 18853 18279 18887
rect 2421 18785 2455 18819
rect 3433 18785 3467 18819
rect 4353 18785 4387 18819
rect 5733 18785 5767 18819
rect 31677 18785 31711 18819
rect 2697 18717 2731 18751
rect 5089 18717 5123 18751
rect 31033 18717 31067 18751
rect 31944 18717 31978 18751
rect 18521 18649 18555 18683
rect 18889 18649 18923 18683
rect 3801 18581 3835 18615
rect 5273 18581 5307 18615
rect 31585 18581 31619 18615
rect 33057 18581 33091 18615
rect 30665 18377 30699 18411
rect 31033 18377 31067 18411
rect 31309 18377 31343 18411
rect 1777 18309 1811 18343
rect 2697 18241 2731 18275
rect 2881 18241 2915 18275
rect 31861 18241 31895 18275
rect 32229 18241 32263 18275
rect 2421 18173 2455 18207
rect 3341 18173 3375 18207
rect 4813 18173 4847 18207
rect 32505 18173 32539 18207
rect 4445 18105 4479 18139
rect 1685 18037 1719 18071
rect 4353 18037 4387 18071
rect 3157 17833 3191 17867
rect 22845 17833 22879 17867
rect 4629 17765 4663 17799
rect 24409 17765 24443 17799
rect 30665 17765 30699 17799
rect 1777 17697 1811 17731
rect 4997 17697 5031 17731
rect 30297 17697 30331 17731
rect 31033 17697 31067 17731
rect 33333 17697 33367 17731
rect 4445 17629 4479 17663
rect 17325 17629 17359 17663
rect 21465 17629 21499 17663
rect 23121 17629 23155 17663
rect 24961 17629 24995 17663
rect 30849 17629 30883 17663
rect 32045 17629 32079 17663
rect 32321 17629 32355 17663
rect 2044 17561 2078 17595
rect 19073 17561 19107 17595
rect 21710 17561 21744 17595
rect 3801 17493 3835 17527
rect 4537 17493 4571 17527
rect 30757 17493 30791 17527
rect 31401 17493 31435 17527
rect 3157 17289 3191 17323
rect 33517 17289 33551 17323
rect 32382 17221 32416 17255
rect 1777 17153 1811 17187
rect 2044 17153 2078 17187
rect 31953 17153 31987 17187
rect 3341 17085 3375 17119
rect 4537 17085 4571 17119
rect 31493 17085 31527 17119
rect 32137 17085 32171 17119
rect 3893 17017 3927 17051
rect 3985 16949 4019 16983
rect 3801 16745 3835 16779
rect 4537 16745 4571 16779
rect 4629 16677 4663 16711
rect 1777 16609 1811 16643
rect 19533 16609 19567 16643
rect 31953 16609 31987 16643
rect 32505 16609 32539 16643
rect 2044 16541 2078 16575
rect 4353 16541 4387 16575
rect 21465 16541 21499 16575
rect 32229 16541 32263 16575
rect 4997 16473 5031 16507
rect 20177 16473 20211 16507
rect 3157 16405 3191 16439
rect 5273 16405 5307 16439
rect 21649 16405 21683 16439
rect 31401 16405 31435 16439
rect 3525 16201 3559 16235
rect 30573 16201 30607 16235
rect 31953 16201 31987 16235
rect 2412 16133 2446 16167
rect 30757 16133 30791 16167
rect 1501 16065 1535 16099
rect 4905 16065 4939 16099
rect 31401 16065 31435 16099
rect 32321 16065 32355 16099
rect 2145 15997 2179 16031
rect 4353 15997 4387 16031
rect 33333 15997 33367 16031
rect 31125 15929 31159 15963
rect 2053 15861 2087 15895
rect 31217 15861 31251 15895
rect 6929 15657 6963 15691
rect 25053 15657 25087 15691
rect 24961 15589 24995 15623
rect 1593 15521 1627 15555
rect 30205 15521 30239 15555
rect 30941 15521 30975 15555
rect 2697 15453 2731 15487
rect 3617 15453 3651 15487
rect 3801 15453 3835 15487
rect 4445 15453 4479 15487
rect 5089 15453 5123 15487
rect 7573 15453 7607 15487
rect 30849 15453 30883 15487
rect 31677 15453 31711 15487
rect 31933 15453 31967 15487
rect 4537 15385 4571 15419
rect 24593 15385 24627 15419
rect 25329 15385 25363 15419
rect 2973 15317 3007 15351
rect 31585 15317 31619 15351
rect 33057 15317 33091 15351
rect 3341 15113 3375 15147
rect 20177 15113 20211 15147
rect 31309 15113 31343 15147
rect 18153 15045 18187 15079
rect 18981 15045 19015 15079
rect 19349 15045 19383 15079
rect 32597 15045 32631 15079
rect 2228 14977 2262 15011
rect 3617 14977 3651 15011
rect 3873 14977 3907 15011
rect 13993 14977 14027 15011
rect 32229 14977 32263 15011
rect 1961 14909 1995 14943
rect 13737 14909 13771 14943
rect 30021 14909 30055 14943
rect 30573 14909 30607 14943
rect 31953 14909 31987 14943
rect 18429 14841 18463 14875
rect 19717 14841 19751 14875
rect 30297 14841 30331 14875
rect 30481 14841 30515 14875
rect 4997 14773 5031 14807
rect 15117 14773 15151 14807
rect 18613 14773 18647 14807
rect 19809 14773 19843 14807
rect 29929 14773 29963 14807
rect 31217 14773 31251 14807
rect 3801 14569 3835 14603
rect 4353 14569 4387 14603
rect 11621 14569 11655 14603
rect 18521 14569 18555 14603
rect 19073 14569 19107 14603
rect 3985 14501 4019 14535
rect 4445 14501 4479 14535
rect 11437 14501 11471 14535
rect 18889 14501 18923 14535
rect 20637 14501 20671 14535
rect 1593 14433 1627 14467
rect 3433 14433 3467 14467
rect 31125 14433 31159 14467
rect 31677 14433 31711 14467
rect 2605 14365 2639 14399
rect 19257 14365 19291 14399
rect 31585 14365 31619 14399
rect 31933 14365 31967 14399
rect 4261 14297 4295 14331
rect 4813 14297 4847 14331
rect 5181 14297 5215 14331
rect 5549 14297 5583 14331
rect 11161 14297 11195 14331
rect 18613 14297 18647 14331
rect 19502 14297 19536 14331
rect 2881 14229 2915 14263
rect 11989 14229 12023 14263
rect 21005 14229 21039 14263
rect 33057 14229 33091 14263
rect 18889 14025 18923 14059
rect 30573 14025 30607 14059
rect 2329 13957 2363 13991
rect 20002 13957 20036 13991
rect 32597 13957 32631 13991
rect 2697 13889 2731 13923
rect 2881 13889 2915 13923
rect 20269 13889 20303 13923
rect 20637 13889 20671 13923
rect 31953 13889 31987 13923
rect 32229 13889 32263 13923
rect 3341 13821 3375 13855
rect 4813 13821 4847 13855
rect 29929 13821 29963 13855
rect 30021 13821 30055 13855
rect 31125 13821 31159 13855
rect 31309 13821 31343 13855
rect 4445 13753 4479 13787
rect 30389 13753 30423 13787
rect 4353 13685 4387 13719
rect 5089 13685 5123 13719
rect 30481 13685 30515 13719
rect 33057 13481 33091 13515
rect 10609 13413 10643 13447
rect 2421 13345 2455 13379
rect 4445 13345 4479 13379
rect 31033 13345 31067 13379
rect 2697 13277 2731 13311
rect 3525 13277 3559 13311
rect 19441 13277 19475 13311
rect 30297 13277 30331 13311
rect 31677 13277 31711 13311
rect 31933 13277 31967 13311
rect 10977 13209 11011 13243
rect 2881 13141 2915 13175
rect 3801 13141 3835 13175
rect 10517 13141 10551 13175
rect 11345 13141 11379 13175
rect 19993 13141 20027 13175
rect 30849 13141 30883 13175
rect 31585 13141 31619 13175
rect 4629 12937 4663 12971
rect 31217 12937 31251 12971
rect 2044 12869 2078 12903
rect 3341 12801 3375 12835
rect 3893 12801 3927 12835
rect 23489 12801 23523 12835
rect 31309 12801 31343 12835
rect 31861 12801 31895 12835
rect 32229 12801 32263 12835
rect 1777 12733 1811 12767
rect 3985 12733 4019 12767
rect 32505 12733 32539 12767
rect 3157 12597 3191 12631
rect 5089 12597 5123 12631
rect 23673 12597 23707 12631
rect 3525 12393 3559 12427
rect 30665 12393 30699 12427
rect 4629 12325 4663 12359
rect 31125 12325 31159 12359
rect 2973 12257 3007 12291
rect 5457 12257 5491 12291
rect 24409 12257 24443 12291
rect 30849 12257 30883 12291
rect 33333 12257 33367 12291
rect 2697 12189 2731 12223
rect 3801 12189 3835 12223
rect 9505 12189 9539 12223
rect 32045 12189 32079 12223
rect 32321 12189 32355 12223
rect 2329 12121 2363 12155
rect 4997 12121 5031 12155
rect 4445 12053 4479 12087
rect 4537 12053 4571 12087
rect 6009 12053 6043 12087
rect 8953 12053 8987 12087
rect 25053 12053 25087 12087
rect 31309 12053 31343 12087
rect 31401 12053 31435 12087
rect 33517 11849 33551 11883
rect 1593 11781 1627 11815
rect 12878 11781 12912 11815
rect 32382 11781 32416 11815
rect 2605 11713 2639 11747
rect 2881 11713 2915 11747
rect 4905 11713 4939 11747
rect 12633 11713 12667 11747
rect 19349 11713 19383 11747
rect 31953 11713 31987 11747
rect 3341 11645 3375 11679
rect 31493 11645 31527 11679
rect 32137 11645 32171 11679
rect 4353 11509 4387 11543
rect 14013 11509 14047 11543
rect 19993 11509 20027 11543
rect 3157 11305 3191 11339
rect 30573 11305 30607 11339
rect 4353 11169 4387 11203
rect 31953 11169 31987 11203
rect 32505 11169 32539 11203
rect 1777 11101 1811 11135
rect 2044 11101 2078 11135
rect 32229 11101 32263 11135
rect 3801 10965 3835 10999
rect 31401 10965 31435 10999
rect 9965 10761 9999 10795
rect 31953 10761 31987 10795
rect 2329 10693 2363 10727
rect 7849 10693 7883 10727
rect 30389 10693 30423 10727
rect 2697 10625 2731 10659
rect 28641 10625 28675 10659
rect 30757 10625 30791 10659
rect 31401 10625 31435 10659
rect 32321 10625 32355 10659
rect 3617 10557 3651 10591
rect 4169 10557 4203 10591
rect 9597 10557 9631 10591
rect 33333 10557 33367 10591
rect 3893 10489 3927 10523
rect 31125 10489 31159 10523
rect 2973 10421 3007 10455
rect 3709 10421 3743 10455
rect 4445 10421 4479 10455
rect 28457 10421 28491 10455
rect 31217 10421 31251 10455
rect 7389 10217 7423 10251
rect 25881 10217 25915 10251
rect 26525 10217 26559 10251
rect 5273 10081 5307 10115
rect 15485 10081 15519 10115
rect 30205 10081 30239 10115
rect 30941 10081 30975 10115
rect 31677 10081 31711 10115
rect 1777 10013 1811 10047
rect 4353 10013 4387 10047
rect 7021 10013 7055 10047
rect 27813 10013 27847 10047
rect 30849 10013 30883 10047
rect 31933 10013 31967 10047
rect 2044 9945 2078 9979
rect 3157 9877 3191 9911
rect 3801 9877 3835 9911
rect 16129 9877 16163 9911
rect 31585 9877 31619 9911
rect 33057 9877 33091 9911
rect 26985 9673 27019 9707
rect 31309 9673 31343 9707
rect 1593 9605 1627 9639
rect 32597 9605 32631 9639
rect 2605 9537 2639 9571
rect 3433 9537 3467 9571
rect 4077 9537 4111 9571
rect 24961 9537 24995 9571
rect 27537 9537 27571 9571
rect 32229 9537 32263 9571
rect 15209 9469 15243 9503
rect 30021 9469 30055 9503
rect 31125 9469 31159 9503
rect 31953 9469 31987 9503
rect 3801 9401 3835 9435
rect 30389 9401 30423 9435
rect 2881 9333 2915 9367
rect 3617 9333 3651 9367
rect 4445 9333 4479 9367
rect 14657 9333 14691 9367
rect 24317 9333 24351 9367
rect 29837 9333 29871 9367
rect 30481 9333 30515 9367
rect 30573 9333 30607 9367
rect 3525 9129 3559 9163
rect 6193 9129 6227 9163
rect 19717 9129 19751 9163
rect 2421 8993 2455 9027
rect 2881 8993 2915 9027
rect 5641 8993 5675 9027
rect 20269 8993 20303 9027
rect 31033 8993 31067 9027
rect 31677 8993 31711 9027
rect 2697 8925 2731 8959
rect 4353 8925 4387 8959
rect 31585 8925 31619 8959
rect 31922 8857 31956 8891
rect 3801 8789 3835 8823
rect 33057 8789 33091 8823
rect 30573 8585 30607 8619
rect 2044 8517 2078 8551
rect 32597 8517 32631 8551
rect 31953 8449 31987 8483
rect 32229 8449 32263 8483
rect 1777 8381 1811 8415
rect 3801 8381 3835 8415
rect 4445 8381 4479 8415
rect 30389 8381 30423 8415
rect 31217 8381 31251 8415
rect 31309 8381 31343 8415
rect 3157 8313 3191 8347
rect 3985 8313 4019 8347
rect 4169 8313 4203 8347
rect 29837 8313 29871 8347
rect 3249 8245 3283 8279
rect 4813 8245 4847 8279
rect 29469 8245 29503 8279
rect 3525 8041 3559 8075
rect 29377 8041 29411 8075
rect 4721 7973 4755 8007
rect 29285 7973 29319 8007
rect 30021 7973 30055 8007
rect 1593 7905 1627 7939
rect 2973 7905 3007 7939
rect 4537 7905 4571 7939
rect 30205 7905 30239 7939
rect 31677 7905 31711 7939
rect 2605 7837 2639 7871
rect 3801 7837 3835 7871
rect 30849 7837 30883 7871
rect 30941 7837 30975 7871
rect 31585 7837 31619 7871
rect 4997 7769 5031 7803
rect 5273 7769 5307 7803
rect 28917 7769 28951 7803
rect 29653 7769 29687 7803
rect 31922 7769 31956 7803
rect 4445 7701 4479 7735
rect 28733 7701 28767 7735
rect 30113 7701 30147 7735
rect 33057 7701 33091 7735
rect 2329 7429 2363 7463
rect 30481 7429 30515 7463
rect 2697 7361 2731 7395
rect 3994 7361 4028 7395
rect 4261 7361 4295 7395
rect 4445 7361 4479 7395
rect 17325 7361 17359 7395
rect 29009 7361 29043 7395
rect 29837 7361 29871 7395
rect 30757 7361 30791 7395
rect 32229 7361 32263 7395
rect 29653 7293 29687 7327
rect 31217 7293 31251 7327
rect 32505 7293 32539 7327
rect 2881 7157 2915 7191
rect 4997 7157 5031 7191
rect 16773 7157 16807 7191
rect 27997 7157 28031 7191
rect 28365 7157 28399 7191
rect 29101 7157 29135 7191
rect 3157 6953 3191 6987
rect 28733 6885 28767 6919
rect 1777 6817 1811 6851
rect 4445 6817 4479 6851
rect 28089 6817 28123 6851
rect 33333 6817 33367 6851
rect 2044 6749 2078 6783
rect 5089 6749 5123 6783
rect 28641 6749 28675 6783
rect 29377 6749 29411 6783
rect 30573 6749 30607 6783
rect 30757 6749 30791 6783
rect 31125 6749 31159 6783
rect 32321 6749 32355 6783
rect 27537 6681 27571 6715
rect 3801 6613 3835 6647
rect 4537 6613 4571 6647
rect 27629 6613 27663 6647
rect 29929 6613 29963 6647
rect 4721 6409 4755 6443
rect 27261 6409 27295 6443
rect 29009 6409 29043 6443
rect 33517 6409 33551 6443
rect 2044 6341 2078 6375
rect 26801 6341 26835 6375
rect 27169 6341 27203 6375
rect 32382 6341 32416 6375
rect 1777 6273 1811 6307
rect 3249 6273 3283 6307
rect 30481 6273 30515 6307
rect 31953 6273 31987 6307
rect 3709 6205 3743 6239
rect 5273 6205 5307 6239
rect 9597 6205 9631 6239
rect 27629 6205 27663 6239
rect 28457 6205 28491 6239
rect 30021 6205 30055 6239
rect 31493 6205 31527 6239
rect 32137 6205 32171 6239
rect 9873 6137 9907 6171
rect 3157 6069 3191 6103
rect 10057 6069 10091 6103
rect 10425 6069 10459 6103
rect 28273 6069 28307 6103
rect 3525 5865 3559 5899
rect 4445 5865 4479 5899
rect 10425 5865 10459 5899
rect 24961 5865 24995 5899
rect 27353 5865 27387 5899
rect 27445 5865 27479 5899
rect 11713 5797 11747 5831
rect 25237 5797 25271 5831
rect 25789 5797 25823 5831
rect 26617 5797 26651 5831
rect 29101 5797 29135 5831
rect 1593 5729 1627 5763
rect 2881 5729 2915 5763
rect 11529 5729 11563 5763
rect 26065 5729 26099 5763
rect 29377 5729 29411 5763
rect 29745 5729 29779 5763
rect 30481 5729 30515 5763
rect 31585 5729 31619 5763
rect 33149 5729 33183 5763
rect 2605 5661 2639 5695
rect 3801 5661 3835 5695
rect 10057 5661 10091 5695
rect 10241 5661 10275 5695
rect 26709 5661 26743 5695
rect 28089 5661 28123 5695
rect 28181 5661 28215 5695
rect 28825 5661 28859 5695
rect 32045 5661 32079 5695
rect 32873 5661 32907 5695
rect 8769 5593 8803 5627
rect 11989 5593 12023 5627
rect 9505 5525 9539 5559
rect 12357 5525 12391 5559
rect 28917 5525 28951 5559
rect 29929 5525 29963 5559
rect 3525 5321 3559 5355
rect 3617 5321 3651 5355
rect 10057 5321 10091 5355
rect 12357 5321 12391 5355
rect 26065 5321 26099 5355
rect 30113 5321 30147 5355
rect 33517 5321 33551 5355
rect 2329 5253 2363 5287
rect 8125 5253 8159 5287
rect 13553 5253 13587 5287
rect 14197 5253 14231 5287
rect 15209 5253 15243 5287
rect 15945 5253 15979 5287
rect 16313 5253 16347 5287
rect 23397 5253 23431 5287
rect 25605 5253 25639 5287
rect 32382 5253 32416 5287
rect 2697 5185 2731 5219
rect 2973 5185 3007 5219
rect 4077 5185 4111 5219
rect 11529 5185 11563 5219
rect 13921 5185 13955 5219
rect 14565 5185 14599 5219
rect 16773 5185 16807 5219
rect 24777 5185 24811 5219
rect 26249 5185 26283 5219
rect 26801 5185 26835 5219
rect 28989 5185 29023 5219
rect 31585 5185 31619 5219
rect 32137 5185 32171 5219
rect 9229 5117 9263 5151
rect 9505 5117 9539 5151
rect 10793 5117 10827 5151
rect 12081 5117 12115 5151
rect 12909 5117 12943 5151
rect 15669 5117 15703 5151
rect 24593 5117 24627 5151
rect 26985 5117 27019 5151
rect 27629 5117 27663 5151
rect 28273 5117 28307 5151
rect 28733 5117 28767 5151
rect 30389 5117 30423 5151
rect 3801 5049 3835 5083
rect 8401 5049 8435 5083
rect 10241 5049 10275 5083
rect 15577 5049 15611 5083
rect 25973 5049 26007 5083
rect 4445 4981 4479 5015
rect 8585 4981 8619 5015
rect 8677 4981 8711 5015
rect 17325 4981 17359 5015
rect 24041 4981 24075 5015
rect 25421 4981 25455 5015
rect 27721 4981 27755 5015
rect 8769 4777 8803 4811
rect 10517 4777 10551 4811
rect 10701 4777 10735 4811
rect 12081 4777 12115 4811
rect 24409 4777 24443 4811
rect 31585 4777 31619 4811
rect 7941 4709 7975 4743
rect 14381 4709 14415 4743
rect 15669 4709 15703 4743
rect 17049 4709 17083 4743
rect 22937 4709 22971 4743
rect 27629 4709 27663 4743
rect 2421 4641 2455 4675
rect 8217 4641 8251 4675
rect 9137 4641 9171 4675
rect 11345 4641 11379 4675
rect 12357 4641 12391 4675
rect 14105 4641 14139 4675
rect 14749 4641 14783 4675
rect 16129 4641 16163 4675
rect 23213 4641 23247 4675
rect 23673 4641 23707 4675
rect 26801 4641 26835 4675
rect 28917 4641 28951 4675
rect 30941 4641 30975 4675
rect 32505 4641 32539 4675
rect 2697 4573 2731 4607
rect 7481 4573 7515 4607
rect 7573 4573 7607 4607
rect 9393 4573 9427 4607
rect 11437 4573 11471 4607
rect 13737 4573 13771 4607
rect 15945 4573 15979 4607
rect 17325 4573 17359 4607
rect 17693 4573 17727 4607
rect 24961 4573 24995 4607
rect 25145 4573 25179 4607
rect 25881 4573 25915 4607
rect 29285 4573 29319 4607
rect 29561 4573 29595 4607
rect 30665 4573 30699 4607
rect 32229 4573 32263 4607
rect 26525 4505 26559 4539
rect 27905 4505 27939 4539
rect 31861 4505 31895 4539
rect 8033 4437 8067 4471
rect 13001 4437 13035 4471
rect 13093 4437 13127 4471
rect 14565 4437 14599 4471
rect 15393 4437 15427 4471
rect 15485 4437 15519 4471
rect 16773 4437 16807 4471
rect 16865 4437 16899 4471
rect 22753 4437 22787 4471
rect 24225 4437 24259 4471
rect 25789 4437 25823 4471
rect 27353 4437 27387 4471
rect 27445 4437 27479 4471
rect 30205 4437 30239 4471
rect 10701 4233 10735 4267
rect 13829 4233 13863 4267
rect 24777 4233 24811 4267
rect 27905 4233 27939 4267
rect 29561 4233 29595 4267
rect 2697 4097 2731 4131
rect 6561 4097 6595 4131
rect 7849 4097 7883 4131
rect 9321 4097 9355 4131
rect 9588 4097 9622 4131
rect 10885 4097 10919 4131
rect 11805 4097 11839 4131
rect 13001 4097 13035 4131
rect 15485 4097 15519 4131
rect 16773 4097 16807 4131
rect 18705 4097 18739 4131
rect 18889 4097 18923 4131
rect 23664 4097 23698 4131
rect 26249 4097 26283 4131
rect 29018 4097 29052 4131
rect 29285 4097 29319 4131
rect 30685 4097 30719 4131
rect 30941 4097 30975 4131
rect 32229 4097 32263 4131
rect 2421 4029 2455 4063
rect 6837 4029 6871 4063
rect 8309 4029 8343 4063
rect 12633 4029 12667 4063
rect 13185 4029 13219 4063
rect 14105 4029 14139 4063
rect 16037 4029 16071 4063
rect 17049 4029 17083 4063
rect 19533 4029 19567 4063
rect 22753 4029 22787 4063
rect 23397 4029 23431 4063
rect 25053 4029 25087 4063
rect 26801 4029 26835 4063
rect 27077 4029 27111 4063
rect 31585 4029 31619 4063
rect 32505 4029 32539 4063
rect 11253 3961 11287 3995
rect 26525 3961 26559 3995
rect 11345 3893 11379 3927
rect 14657 3893 14691 3927
rect 18153 3893 18187 3927
rect 23305 3893 23339 3927
rect 26341 3893 26375 3927
rect 27629 3893 27663 3927
rect 31033 3893 31067 3927
rect 11529 3689 11563 3723
rect 14105 3689 14139 3723
rect 19901 3689 19935 3723
rect 22109 3689 22143 3723
rect 24409 3689 24443 3723
rect 24961 3689 24995 3723
rect 32597 3689 32631 3723
rect 32873 3689 32907 3723
rect 18429 3621 18463 3655
rect 23581 3621 23615 3655
rect 24041 3621 24075 3655
rect 24501 3621 24535 3655
rect 1593 3553 1627 3587
rect 6653 3553 6687 3587
rect 10149 3553 10183 3587
rect 13645 3553 13679 3587
rect 19257 3553 19291 3587
rect 22201 3553 22235 3587
rect 26893 3553 26927 3587
rect 33425 3553 33459 3587
rect 2605 3485 2639 3519
rect 5733 3485 5767 3519
rect 7205 3485 7239 3519
rect 8677 3485 8711 3519
rect 9965 3485 9999 3519
rect 13001 3485 13035 3519
rect 15485 3485 15519 3519
rect 15577 3485 15611 3519
rect 17049 3485 17083 3519
rect 17305 3485 17339 3519
rect 20361 3485 20395 3519
rect 22468 3485 22502 3519
rect 24869 3485 24903 3519
rect 26085 3485 26119 3519
rect 26341 3485 26375 3519
rect 26433 3485 26467 3519
rect 27997 3485 28031 3519
rect 28549 3485 28583 3519
rect 30205 3485 30239 3519
rect 31769 3485 31803 3519
rect 32137 3485 32171 3519
rect 32781 3485 32815 3519
rect 5365 3417 5399 3451
rect 8309 3417 8343 3451
rect 10394 3417 10428 3451
rect 12734 3417 12768 3451
rect 15240 3417 15274 3451
rect 15844 3417 15878 3451
rect 20913 3417 20947 3451
rect 23673 3417 23707 3451
rect 29837 3417 29871 3451
rect 9413 3349 9447 3383
rect 11621 3349 11655 3383
rect 13093 3349 13127 3383
rect 16957 3349 16991 3383
rect 24133 3349 24167 3383
rect 29009 3349 29043 3383
rect 29377 3349 29411 3383
rect 30665 3349 30699 3383
rect 31309 3349 31343 3383
rect 9873 3145 9907 3179
rect 13185 3145 13219 3179
rect 16681 3145 16715 3179
rect 22293 3145 22327 3179
rect 26985 3145 27019 3179
rect 31401 3145 31435 3179
rect 33517 3145 33551 3179
rect 25890 3077 25924 3111
rect 31861 3077 31895 3111
rect 2697 3009 2731 3043
rect 6009 3009 6043 3043
rect 8309 3009 8343 3043
rect 8493 3009 8527 3043
rect 8760 3009 8794 3043
rect 9965 3009 9999 3043
rect 13001 3009 13035 3043
rect 14309 3009 14343 3043
rect 14565 3009 14599 3043
rect 16313 3009 16347 3043
rect 18153 3009 18187 3043
rect 19717 3009 19751 3043
rect 23121 3009 23155 3043
rect 23305 3009 23339 3043
rect 26157 3009 26191 3043
rect 28098 3009 28132 3043
rect 29837 3009 29871 3043
rect 29929 3009 29963 3043
rect 32137 3009 32171 3043
rect 32393 3009 32427 3043
rect 2421 2941 2455 2975
rect 4997 2941 5031 2975
rect 7941 2941 7975 2975
rect 10517 2941 10551 2975
rect 12541 2941 12575 2975
rect 15301 2941 15335 2975
rect 17325 2941 17359 2975
rect 17693 2941 17727 2975
rect 19993 2941 20027 2975
rect 22845 2941 22879 2975
rect 23765 2941 23799 2975
rect 26341 2941 26375 2975
rect 28365 2941 28399 2975
rect 28641 2941 28675 2975
rect 30389 2941 30423 2975
rect 24777 2873 24811 2907
rect 26709 2873 26743 2907
rect 31493 2873 31527 2907
rect 26801 2805 26835 2839
rect 12449 2601 12483 2635
rect 14381 2601 14415 2635
rect 17325 2601 17359 2635
rect 31677 2601 31711 2635
rect 2881 2533 2915 2567
rect 21557 2533 21591 2567
rect 23949 2533 23983 2567
rect 25513 2533 25547 2567
rect 28089 2533 28123 2567
rect 30573 2533 30607 2567
rect 1593 2465 1627 2499
rect 5825 2465 5859 2499
rect 8401 2465 8435 2499
rect 10885 2465 10919 2499
rect 11805 2465 11839 2499
rect 13277 2465 13311 2499
rect 14933 2465 14967 2499
rect 16037 2465 16071 2499
rect 16773 2465 16807 2499
rect 18153 2465 18187 2499
rect 19717 2465 19751 2499
rect 21649 2465 21683 2499
rect 22293 2465 22327 2499
rect 23305 2465 23339 2499
rect 25053 2465 25087 2499
rect 27353 2465 27387 2499
rect 30021 2465 30055 2499
rect 32597 2465 32631 2499
rect 2605 2397 2639 2431
rect 3157 2397 3191 2431
rect 3801 2397 3835 2431
rect 6101 2397 6135 2431
rect 8677 2397 8711 2431
rect 9229 2397 9263 2431
rect 9781 2397 9815 2431
rect 11345 2397 11379 2431
rect 12541 2397 12575 2431
rect 16497 2397 16531 2431
rect 17693 2397 17727 2431
rect 19349 2397 19383 2431
rect 21925 2397 21959 2431
rect 24501 2397 24535 2431
rect 25881 2397 25915 2431
rect 26433 2397 26467 2431
rect 27077 2397 27111 2431
rect 29009 2397 29043 2431
rect 29653 2397 29687 2431
rect 31033 2397 31067 2431
rect 32137 2397 32171 2431
rect 21097 2329 21131 2363
rect 21189 2329 21223 2363
rect 28457 2329 28491 2363
<< metal1 >>
rect 1104 32666 34016 32688
rect 1104 32614 9138 32666
rect 9190 32614 9202 32666
rect 9254 32614 9266 32666
rect 9318 32614 9330 32666
rect 9382 32614 9394 32666
rect 9446 32614 17326 32666
rect 17378 32614 17390 32666
rect 17442 32614 17454 32666
rect 17506 32614 17518 32666
rect 17570 32614 17582 32666
rect 17634 32614 25514 32666
rect 25566 32614 25578 32666
rect 25630 32614 25642 32666
rect 25694 32614 25706 32666
rect 25758 32614 25770 32666
rect 25822 32614 33702 32666
rect 33754 32614 33766 32666
rect 33818 32614 33830 32666
rect 33882 32614 33894 32666
rect 33946 32614 33958 32666
rect 34010 32614 34016 32666
rect 1104 32592 34016 32614
rect 5261 32487 5319 32493
rect 5261 32453 5273 32487
rect 5307 32484 5319 32487
rect 5718 32484 5724 32496
rect 5307 32456 5724 32484
rect 5307 32453 5319 32456
rect 5261 32447 5319 32453
rect 5718 32444 5724 32456
rect 5776 32444 5782 32496
rect 7006 32484 7012 32496
rect 5828 32456 7012 32484
rect 2866 32376 2872 32428
rect 2924 32376 2930 32428
rect 4065 32419 4123 32425
rect 4065 32385 4077 32419
rect 4111 32416 4123 32419
rect 5828 32416 5856 32456
rect 7006 32444 7012 32456
rect 7064 32444 7070 32496
rect 10410 32444 10416 32496
rect 10468 32444 10474 32496
rect 15194 32444 15200 32496
rect 15252 32444 15258 32496
rect 21358 32444 21364 32496
rect 21416 32484 21422 32496
rect 21416 32456 23428 32484
rect 21416 32444 21422 32456
rect 4111 32388 5856 32416
rect 6181 32419 6239 32425
rect 4111 32385 4123 32388
rect 4065 32379 4123 32385
rect 6181 32385 6193 32419
rect 6227 32416 6239 32419
rect 6227 32388 6592 32416
rect 6227 32385 6239 32388
rect 6181 32379 6239 32385
rect 1578 32308 1584 32360
rect 1636 32308 1642 32360
rect 2593 32351 2651 32357
rect 2593 32317 2605 32351
rect 2639 32348 2651 32351
rect 2639 32320 4384 32348
rect 2639 32317 2651 32320
rect 2593 32311 2651 32317
rect 4356 32224 4384 32320
rect 6564 32224 6592 32388
rect 8662 32376 8668 32428
rect 8720 32376 8726 32428
rect 11146 32376 11152 32428
rect 11204 32376 11210 32428
rect 13538 32376 13544 32428
rect 13596 32376 13602 32428
rect 13909 32419 13967 32425
rect 13909 32385 13921 32419
rect 13955 32416 13967 32419
rect 14274 32416 14280 32428
rect 13955 32388 14280 32416
rect 13955 32385 13967 32388
rect 13909 32379 13967 32385
rect 14274 32376 14280 32388
rect 14332 32376 14338 32428
rect 6730 32308 6736 32360
rect 6788 32308 6794 32360
rect 8386 32308 8392 32360
rect 8444 32308 8450 32360
rect 9858 32308 9864 32360
rect 9916 32308 9922 32360
rect 11885 32351 11943 32357
rect 11885 32317 11897 32351
rect 11931 32348 11943 32351
rect 12526 32348 12532 32360
rect 11931 32320 12532 32348
rect 11931 32317 11943 32320
rect 11885 32311 11943 32317
rect 12526 32308 12532 32320
rect 12584 32308 12590 32360
rect 13449 32351 13507 32357
rect 13449 32317 13461 32351
rect 13495 32348 13507 32351
rect 13556 32348 13584 32376
rect 13495 32320 13584 32348
rect 13495 32317 13507 32320
rect 13449 32311 13507 32317
rect 14458 32308 14464 32360
rect 14516 32308 14522 32360
rect 15212 32348 15240 32444
rect 15286 32376 15292 32428
rect 15344 32376 15350 32428
rect 17126 32376 17132 32428
rect 17184 32416 17190 32428
rect 17773 32419 17831 32425
rect 17773 32416 17785 32419
rect 17184 32388 17785 32416
rect 17184 32376 17190 32388
rect 17773 32385 17785 32388
rect 17819 32385 17831 32419
rect 17773 32379 17831 32385
rect 18325 32419 18383 32425
rect 18325 32385 18337 32419
rect 18371 32416 18383 32419
rect 19245 32419 19303 32425
rect 19245 32416 19257 32419
rect 18371 32388 19257 32416
rect 18371 32385 18383 32388
rect 18325 32379 18383 32385
rect 19245 32385 19257 32388
rect 19291 32385 19303 32419
rect 19245 32379 19303 32385
rect 21818 32376 21824 32428
rect 21876 32376 21882 32428
rect 23293 32419 23351 32425
rect 23293 32416 23305 32419
rect 22020 32388 23305 32416
rect 22020 32360 22048 32388
rect 23293 32385 23305 32388
rect 23339 32385 23351 32419
rect 23293 32379 23351 32385
rect 15565 32351 15623 32357
rect 15565 32348 15577 32351
rect 15212 32320 15577 32348
rect 15565 32317 15577 32320
rect 15611 32317 15623 32351
rect 15565 32311 15623 32317
rect 17497 32351 17555 32357
rect 17497 32317 17509 32351
rect 17543 32348 17555 32351
rect 17678 32348 17684 32360
rect 17543 32320 17684 32348
rect 17543 32317 17555 32320
rect 17497 32311 17555 32317
rect 17678 32308 17684 32320
rect 17736 32308 17742 32360
rect 18506 32308 18512 32360
rect 18564 32348 18570 32360
rect 19705 32351 19763 32357
rect 19705 32348 19717 32351
rect 18564 32320 19717 32348
rect 18564 32308 18570 32320
rect 19705 32317 19717 32320
rect 19751 32317 19763 32351
rect 19705 32311 19763 32317
rect 20898 32308 20904 32360
rect 20956 32348 20962 32360
rect 21269 32351 21327 32357
rect 21269 32348 21281 32351
rect 20956 32320 21281 32348
rect 20956 32308 20962 32320
rect 21269 32317 21281 32320
rect 21315 32317 21327 32351
rect 21269 32311 21327 32317
rect 22002 32308 22008 32360
rect 22060 32308 22066 32360
rect 22281 32351 22339 32357
rect 22281 32317 22293 32351
rect 22327 32317 22339 32351
rect 22281 32311 22339 32317
rect 9217 32283 9275 32289
rect 9217 32249 9229 32283
rect 9263 32280 9275 32283
rect 9398 32280 9404 32292
rect 9263 32252 9404 32280
rect 9263 32249 9275 32252
rect 9217 32243 9275 32249
rect 9398 32240 9404 32252
rect 9456 32280 9462 32292
rect 12894 32280 12900 32292
rect 9456 32252 12900 32280
rect 9456 32240 9462 32252
rect 12894 32240 12900 32252
rect 12952 32240 12958 32292
rect 20162 32240 20168 32292
rect 20220 32280 20226 32292
rect 22296 32280 22324 32311
rect 20220 32252 22324 32280
rect 23308 32280 23336 32379
rect 23400 32348 23428 32456
rect 29178 32444 29184 32496
rect 29236 32484 29242 32496
rect 29236 32456 31754 32484
rect 29236 32444 29242 32456
rect 24394 32376 24400 32428
rect 24452 32376 24458 32428
rect 25038 32376 25044 32428
rect 25096 32416 25102 32428
rect 25096 32388 26556 32416
rect 25096 32376 25102 32388
rect 24857 32351 24915 32357
rect 24857 32348 24869 32351
rect 23400 32320 24869 32348
rect 24857 32317 24869 32320
rect 24903 32317 24915 32351
rect 24857 32311 24915 32317
rect 26050 32308 26056 32360
rect 26108 32308 26114 32360
rect 26418 32308 26424 32360
rect 26476 32308 26482 32360
rect 26528 32348 26556 32388
rect 26970 32376 26976 32428
rect 27028 32376 27034 32428
rect 28166 32376 28172 32428
rect 28224 32416 28230 32428
rect 29549 32419 29607 32425
rect 29549 32416 29561 32419
rect 28224 32388 29561 32416
rect 28224 32376 28230 32388
rect 29549 32385 29561 32388
rect 29595 32385 29607 32419
rect 29549 32379 29607 32385
rect 27433 32351 27491 32357
rect 27433 32348 27445 32351
rect 26528 32320 27445 32348
rect 27433 32317 27445 32320
rect 27479 32317 27491 32351
rect 27433 32311 27491 32317
rect 28994 32308 29000 32360
rect 29052 32308 29058 32360
rect 30009 32351 30067 32357
rect 30009 32317 30021 32351
rect 30055 32317 30067 32351
rect 30009 32311 30067 32317
rect 25869 32283 25927 32289
rect 25869 32280 25881 32283
rect 23308 32252 25881 32280
rect 20220 32240 20226 32252
rect 25869 32249 25881 32252
rect 25915 32249 25927 32283
rect 26068 32280 26096 32308
rect 30024 32280 30052 32311
rect 30374 32308 30380 32360
rect 30432 32348 30438 32360
rect 31573 32351 31631 32357
rect 31573 32348 31585 32351
rect 30432 32320 31585 32348
rect 30432 32308 30438 32320
rect 31573 32317 31585 32320
rect 31619 32317 31631 32351
rect 31726 32348 31754 32456
rect 32122 32376 32128 32428
rect 32180 32376 32186 32428
rect 32585 32351 32643 32357
rect 32585 32348 32597 32351
rect 31726 32320 32597 32348
rect 31573 32311 31631 32317
rect 32585 32317 32597 32320
rect 32631 32317 32643 32351
rect 32585 32311 32643 32317
rect 26068 32252 30052 32280
rect 25869 32243 25927 32249
rect 2130 32172 2136 32224
rect 2188 32172 2194 32224
rect 4338 32172 4344 32224
rect 4396 32172 4402 32224
rect 4709 32215 4767 32221
rect 4709 32181 4721 32215
rect 4755 32212 4767 32215
rect 6270 32212 6276 32224
rect 4755 32184 6276 32212
rect 4755 32181 4767 32184
rect 4709 32175 4767 32181
rect 6270 32172 6276 32184
rect 6328 32172 6334 32224
rect 6546 32172 6552 32224
rect 6604 32172 6610 32224
rect 7285 32215 7343 32221
rect 7285 32181 7297 32215
rect 7331 32212 7343 32215
rect 8294 32212 8300 32224
rect 7331 32184 8300 32212
rect 7331 32181 7343 32184
rect 7285 32175 7343 32181
rect 8294 32172 8300 32184
rect 8352 32172 8358 32224
rect 12437 32215 12495 32221
rect 12437 32181 12449 32215
rect 12483 32212 12495 32215
rect 13630 32212 13636 32224
rect 12483 32184 13636 32212
rect 12483 32181 12495 32184
rect 12437 32175 12495 32181
rect 13630 32172 13636 32184
rect 13688 32172 13694 32224
rect 15013 32215 15071 32221
rect 15013 32181 15025 32215
rect 15059 32212 15071 32215
rect 16114 32212 16120 32224
rect 15059 32184 16120 32212
rect 15059 32181 15071 32184
rect 15013 32175 15071 32181
rect 16114 32172 16120 32184
rect 16172 32172 16178 32224
rect 16850 32172 16856 32224
rect 16908 32172 16914 32224
rect 18506 32172 18512 32224
rect 18564 32212 18570 32224
rect 20717 32215 20775 32221
rect 20717 32212 20729 32215
rect 18564 32184 20729 32212
rect 18564 32172 18570 32184
rect 20717 32181 20729 32184
rect 20763 32181 20775 32215
rect 20717 32175 20775 32181
rect 23937 32215 23995 32221
rect 23937 32181 23949 32215
rect 23983 32212 23995 32215
rect 26142 32212 26148 32224
rect 23983 32184 26148 32212
rect 23983 32181 23995 32184
rect 23937 32175 23995 32181
rect 26142 32172 26148 32184
rect 26200 32172 26206 32224
rect 26878 32172 26884 32224
rect 26936 32212 26942 32224
rect 28445 32215 28503 32221
rect 28445 32212 28457 32215
rect 26936 32184 28457 32212
rect 26936 32172 26942 32184
rect 28445 32181 28457 32184
rect 28491 32181 28503 32215
rect 28445 32175 28503 32181
rect 31018 32172 31024 32224
rect 31076 32172 31082 32224
rect 1104 32122 33856 32144
rect 1104 32070 5044 32122
rect 5096 32070 5108 32122
rect 5160 32070 5172 32122
rect 5224 32070 5236 32122
rect 5288 32070 5300 32122
rect 5352 32070 13232 32122
rect 13284 32070 13296 32122
rect 13348 32070 13360 32122
rect 13412 32070 13424 32122
rect 13476 32070 13488 32122
rect 13540 32070 21420 32122
rect 21472 32070 21484 32122
rect 21536 32070 21548 32122
rect 21600 32070 21612 32122
rect 21664 32070 21676 32122
rect 21728 32070 29608 32122
rect 29660 32070 29672 32122
rect 29724 32070 29736 32122
rect 29788 32070 29800 32122
rect 29852 32070 29864 32122
rect 29916 32070 33856 32122
rect 1104 32048 33856 32070
rect 2130 31968 2136 32020
rect 2188 31968 2194 32020
rect 2866 31968 2872 32020
rect 2924 32008 2930 32020
rect 2961 32011 3019 32017
rect 2961 32008 2973 32011
rect 2924 31980 2973 32008
rect 2924 31968 2930 31980
rect 2961 31977 2973 31980
rect 3007 31977 3019 32011
rect 2961 31971 3019 31977
rect 6730 31968 6736 32020
rect 6788 32008 6794 32020
rect 9398 32008 9404 32020
rect 6788 31980 9260 32008
rect 6788 31968 6794 31980
rect 2148 31872 2176 31968
rect 3881 31943 3939 31949
rect 3881 31940 3893 31943
rect 3528 31912 3893 31940
rect 3528 31881 3556 31912
rect 3881 31909 3893 31912
rect 3927 31909 3939 31943
rect 3881 31903 3939 31909
rect 3513 31875 3571 31881
rect 3513 31872 3525 31875
rect 2148 31844 3525 31872
rect 3513 31841 3525 31844
rect 3559 31841 3571 31875
rect 3513 31835 3571 31841
rect 4154 31832 4160 31884
rect 4212 31872 4218 31884
rect 4801 31875 4859 31881
rect 4801 31872 4813 31875
rect 4212 31844 4813 31872
rect 4212 31832 4218 31844
rect 4801 31841 4813 31844
rect 4847 31841 4859 31875
rect 4801 31835 4859 31841
rect 6546 31832 6552 31884
rect 6604 31832 6610 31884
rect 7282 31832 7288 31884
rect 7340 31872 7346 31884
rect 7837 31875 7895 31881
rect 7837 31872 7849 31875
rect 7340 31844 7849 31872
rect 7340 31832 7346 31844
rect 7837 31841 7849 31844
rect 7883 31841 7895 31875
rect 9232 31872 9260 31980
rect 9324 31980 9404 32008
rect 9324 31949 9352 31980
rect 9398 31968 9404 31980
rect 9456 31968 9462 32020
rect 11146 31968 11152 32020
rect 11204 31968 11210 32020
rect 15286 31968 15292 32020
rect 15344 31968 15350 32020
rect 16850 31968 16856 32020
rect 16908 31968 16914 32020
rect 21818 31968 21824 32020
rect 21876 31968 21882 32020
rect 24394 31968 24400 32020
rect 24452 31968 24458 32020
rect 27614 31968 27620 32020
rect 27672 32008 27678 32020
rect 27672 31980 30144 32008
rect 27672 31968 27678 31980
rect 9309 31943 9367 31949
rect 9309 31909 9321 31943
rect 9355 31909 9367 31943
rect 9309 31903 9367 31909
rect 9493 31943 9551 31949
rect 9493 31909 9505 31943
rect 9539 31940 9551 31943
rect 11054 31940 11060 31952
rect 9539 31912 11060 31940
rect 9539 31909 9551 31912
rect 9493 31903 9551 31909
rect 11054 31900 11060 31912
rect 11112 31900 11118 31952
rect 9674 31872 9680 31884
rect 9232 31844 9680 31872
rect 7837 31835 7895 31841
rect 9674 31832 9680 31844
rect 9732 31832 9738 31884
rect 10597 31875 10655 31881
rect 10597 31841 10609 31875
rect 10643 31872 10655 31875
rect 11164 31872 11192 31968
rect 10643 31844 11192 31872
rect 12069 31875 12127 31881
rect 10643 31841 10655 31844
rect 10597 31835 10655 31841
rect 12069 31841 12081 31875
rect 12115 31872 12127 31875
rect 12989 31875 13047 31881
rect 12115 31844 12572 31872
rect 12115 31841 12127 31844
rect 12069 31835 12127 31841
rect 1394 31764 1400 31816
rect 1452 31804 1458 31816
rect 1581 31807 1639 31813
rect 1581 31804 1593 31807
rect 1452 31776 1593 31804
rect 1452 31764 1458 31776
rect 1581 31773 1593 31776
rect 1627 31773 1639 31807
rect 1581 31767 1639 31773
rect 2590 31764 2596 31816
rect 2648 31764 2654 31816
rect 4249 31807 4307 31813
rect 4249 31773 4261 31807
rect 4295 31773 4307 31807
rect 4249 31767 4307 31773
rect 4264 31736 4292 31767
rect 4338 31764 4344 31816
rect 4396 31764 4402 31816
rect 6178 31804 6184 31816
rect 4448 31776 6184 31804
rect 4448 31736 4476 31776
rect 6178 31764 6184 31776
rect 6236 31764 6242 31816
rect 7098 31764 7104 31816
rect 7156 31764 7162 31816
rect 7466 31764 7472 31816
rect 7524 31764 7530 31816
rect 9769 31807 9827 31813
rect 9769 31804 9781 31807
rect 9048 31776 9781 31804
rect 9048 31745 9076 31776
rect 9769 31773 9781 31776
rect 9815 31773 9827 31807
rect 9769 31767 9827 31773
rect 10873 31807 10931 31813
rect 10873 31773 10885 31807
rect 10919 31804 10931 31807
rect 10962 31804 10968 31816
rect 10919 31776 10968 31804
rect 10919 31773 10931 31776
rect 10873 31767 10931 31773
rect 10962 31764 10968 31776
rect 11020 31764 11026 31816
rect 12342 31764 12348 31816
rect 12400 31764 12406 31816
rect 12544 31813 12572 31844
rect 12989 31841 13001 31875
rect 13035 31841 13047 31875
rect 15304 31872 15332 31968
rect 15473 31875 15531 31881
rect 15473 31872 15485 31875
rect 15304 31844 15485 31872
rect 12989 31835 13047 31841
rect 15473 31841 15485 31844
rect 15519 31841 15531 31875
rect 15473 31835 15531 31841
rect 12529 31807 12587 31813
rect 12529 31773 12541 31807
rect 12575 31773 12587 31807
rect 12529 31767 12587 31773
rect 9033 31739 9091 31745
rect 9033 31736 9045 31739
rect 4264 31708 4476 31736
rect 8956 31708 9045 31736
rect 8956 31680 8984 31708
rect 9033 31705 9045 31708
rect 9079 31705 9091 31739
rect 9033 31699 9091 31705
rect 11974 31696 11980 31748
rect 12032 31736 12038 31748
rect 13004 31736 13032 31835
rect 14461 31807 14519 31813
rect 14461 31773 14473 31807
rect 14507 31804 14519 31807
rect 14550 31804 14556 31816
rect 14507 31776 14556 31804
rect 14507 31773 14519 31776
rect 14461 31767 14519 31773
rect 14550 31764 14556 31776
rect 14608 31764 14614 31816
rect 16868 31813 16896 31968
rect 18506 31832 18512 31884
rect 18564 31832 18570 31884
rect 20533 31875 20591 31881
rect 20533 31841 20545 31875
rect 20579 31872 20591 31875
rect 21836 31872 21864 31968
rect 20579 31844 21864 31872
rect 22833 31875 22891 31881
rect 20579 31841 20591 31844
rect 20533 31835 20591 31841
rect 22833 31841 22845 31875
rect 22879 31872 22891 31875
rect 24412 31872 24440 31968
rect 22879 31844 24440 31872
rect 25225 31875 25283 31881
rect 22879 31841 22891 31844
rect 22833 31835 22891 31841
rect 25225 31841 25237 31875
rect 25271 31872 25283 31875
rect 26970 31872 26976 31884
rect 25271 31844 26976 31872
rect 25271 31841 25283 31844
rect 25225 31835 25283 31841
rect 26970 31832 26976 31844
rect 27028 31832 27034 31884
rect 28166 31832 28172 31884
rect 28224 31832 28230 31884
rect 30116 31881 30144 31980
rect 30101 31875 30159 31881
rect 30101 31841 30113 31875
rect 30147 31841 30159 31875
rect 30101 31835 30159 31841
rect 32033 31875 32091 31881
rect 32033 31841 32045 31875
rect 32079 31872 32091 31875
rect 32122 31872 32128 31884
rect 32079 31844 32128 31872
rect 32079 31841 32091 31844
rect 32033 31835 32091 31841
rect 32122 31832 32128 31844
rect 32180 31832 32186 31884
rect 15013 31807 15071 31813
rect 15013 31773 15025 31807
rect 15059 31804 15071 31807
rect 15197 31807 15255 31813
rect 15197 31804 15209 31807
rect 15059 31776 15209 31804
rect 15059 31773 15071 31776
rect 15013 31767 15071 31773
rect 15197 31773 15209 31776
rect 15243 31773 15255 31807
rect 15197 31767 15255 31773
rect 16853 31807 16911 31813
rect 16853 31773 16865 31807
rect 16899 31773 16911 31807
rect 16853 31767 16911 31773
rect 19061 31807 19119 31813
rect 19061 31773 19073 31807
rect 19107 31804 19119 31807
rect 19981 31807 20039 31813
rect 19981 31804 19993 31807
rect 19107 31776 19993 31804
rect 19107 31773 19119 31776
rect 19061 31767 19119 31773
rect 19981 31773 19993 31776
rect 20027 31773 20039 31807
rect 20901 31807 20959 31813
rect 20901 31804 20913 31807
rect 19981 31767 20039 31773
rect 20272 31776 20913 31804
rect 12032 31708 13032 31736
rect 12032 31696 12038 31708
rect 17218 31696 17224 31748
rect 17276 31696 17282 31748
rect 20272 31680 20300 31776
rect 20901 31773 20913 31776
rect 20947 31804 20959 31807
rect 22281 31807 22339 31813
rect 22281 31804 22293 31807
rect 20947 31776 22293 31804
rect 20947 31773 20959 31776
rect 20901 31767 20959 31773
rect 22281 31773 22293 31776
rect 22327 31804 22339 31807
rect 22370 31804 22376 31816
rect 22327 31776 22376 31804
rect 22327 31773 22339 31776
rect 22281 31767 22339 31773
rect 22370 31764 22376 31776
rect 22428 31764 22434 31816
rect 23109 31807 23167 31813
rect 23109 31773 23121 31807
rect 23155 31804 23167 31807
rect 23293 31807 23351 31813
rect 23293 31804 23305 31807
rect 23155 31776 23305 31804
rect 23155 31773 23167 31776
rect 23109 31767 23167 31773
rect 23293 31773 23305 31776
rect 23339 31773 23351 31807
rect 23293 31767 23351 31773
rect 23382 31764 23388 31816
rect 23440 31804 23446 31816
rect 23845 31807 23903 31813
rect 23845 31804 23857 31807
rect 23440 31776 23857 31804
rect 23440 31764 23446 31776
rect 23845 31773 23857 31776
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 24670 31764 24676 31816
rect 24728 31764 24734 31816
rect 26142 31764 26148 31816
rect 26200 31764 26206 31816
rect 27614 31764 27620 31816
rect 27672 31764 27678 31816
rect 29086 31764 29092 31816
rect 29144 31804 29150 31816
rect 29549 31807 29607 31813
rect 29549 31804 29561 31807
rect 29144 31776 29561 31804
rect 29144 31764 29150 31776
rect 29549 31773 29561 31776
rect 29595 31773 29607 31807
rect 29549 31767 29607 31773
rect 32309 31807 32367 31813
rect 32309 31773 32321 31807
rect 32355 31804 32367 31807
rect 32493 31807 32551 31813
rect 32493 31804 32505 31807
rect 32355 31776 32505 31804
rect 32355 31773 32367 31776
rect 32309 31767 32367 31773
rect 32493 31773 32505 31776
rect 32539 31773 32551 31807
rect 32493 31767 32551 31773
rect 33042 31764 33048 31816
rect 33100 31764 33106 31816
rect 26510 31696 26516 31748
rect 26568 31696 26574 31748
rect 26988 31708 27292 31736
rect 3786 31628 3792 31680
rect 3844 31628 3850 31680
rect 8938 31628 8944 31680
rect 8996 31628 9002 31680
rect 18138 31628 18144 31680
rect 18196 31628 18202 31680
rect 20254 31628 20260 31680
rect 20312 31628 20318 31680
rect 21266 31628 21272 31680
rect 21324 31628 21330 31680
rect 25406 31628 25412 31680
rect 25464 31668 25470 31680
rect 25685 31671 25743 31677
rect 25685 31668 25697 31671
rect 25464 31640 25697 31668
rect 25464 31628 25470 31640
rect 25685 31637 25697 31640
rect 25731 31668 25743 31671
rect 26988 31668 27016 31708
rect 25731 31640 27016 31668
rect 25731 31637 25743 31640
rect 25685 31631 25743 31637
rect 27154 31628 27160 31680
rect 27212 31628 27218 31680
rect 27264 31668 27292 31708
rect 28534 31668 28540 31680
rect 27264 31640 28540 31668
rect 28534 31628 28540 31640
rect 28592 31628 28598 31680
rect 30190 31628 30196 31680
rect 30248 31668 30254 31680
rect 31205 31671 31263 31677
rect 31205 31668 31217 31671
rect 30248 31640 31217 31668
rect 30248 31628 30254 31640
rect 31205 31637 31217 31640
rect 31251 31668 31263 31671
rect 31846 31668 31852 31680
rect 31251 31640 31852 31668
rect 31251 31637 31263 31640
rect 31205 31631 31263 31637
rect 31846 31628 31852 31640
rect 31904 31628 31910 31680
rect 1104 31578 34016 31600
rect 1104 31526 9138 31578
rect 9190 31526 9202 31578
rect 9254 31526 9266 31578
rect 9318 31526 9330 31578
rect 9382 31526 9394 31578
rect 9446 31526 17326 31578
rect 17378 31526 17390 31578
rect 17442 31526 17454 31578
rect 17506 31526 17518 31578
rect 17570 31526 17582 31578
rect 17634 31526 25514 31578
rect 25566 31526 25578 31578
rect 25630 31526 25642 31578
rect 25694 31526 25706 31578
rect 25758 31526 25770 31578
rect 25822 31526 33702 31578
rect 33754 31526 33766 31578
rect 33818 31526 33830 31578
rect 33882 31526 33894 31578
rect 33946 31526 33958 31578
rect 34010 31526 34016 31578
rect 1104 31504 34016 31526
rect 1578 31424 1584 31476
rect 1636 31464 1642 31476
rect 1765 31467 1823 31473
rect 1765 31464 1777 31467
rect 1636 31436 1777 31464
rect 1636 31424 1642 31436
rect 1765 31433 1777 31436
rect 1811 31433 1823 31467
rect 4249 31467 4307 31473
rect 4249 31464 4261 31467
rect 1765 31427 1823 31433
rect 2608 31436 4261 31464
rect 2501 31331 2559 31337
rect 2501 31328 2513 31331
rect 1780 31300 2513 31328
rect 1780 31272 1808 31300
rect 2501 31297 2513 31300
rect 2547 31297 2559 31331
rect 2501 31291 2559 31297
rect 1762 31220 1768 31272
rect 1820 31220 1826 31272
rect 2409 31263 2467 31269
rect 2409 31229 2421 31263
rect 2455 31260 2467 31263
rect 2608 31260 2636 31436
rect 4249 31433 4261 31436
rect 4295 31433 4307 31467
rect 8297 31467 8355 31473
rect 8297 31464 8309 31467
rect 4249 31427 4307 31433
rect 8128 31436 8309 31464
rect 2768 31399 2826 31405
rect 2768 31365 2780 31399
rect 2814 31396 2826 31399
rect 3786 31396 3792 31408
rect 2814 31368 3792 31396
rect 2814 31365 2826 31368
rect 2768 31359 2826 31365
rect 3786 31356 3792 31368
rect 3844 31356 3850 31408
rect 5994 31396 6000 31408
rect 3896 31368 6000 31396
rect 2455 31232 2636 31260
rect 2455 31229 2467 31232
rect 2409 31223 2467 31229
rect 3896 31201 3924 31368
rect 5994 31356 6000 31368
rect 6052 31356 6058 31408
rect 6178 31356 6184 31408
rect 6236 31356 6242 31408
rect 7960 31399 8018 31405
rect 7960 31365 7972 31399
rect 8006 31396 8018 31399
rect 8128 31396 8156 31436
rect 8297 31433 8309 31436
rect 8343 31433 8355 31467
rect 8297 31427 8355 31433
rect 12526 31424 12532 31476
rect 12584 31464 12590 31476
rect 13173 31467 13231 31473
rect 13173 31464 13185 31467
rect 12584 31436 13185 31464
rect 12584 31424 12590 31436
rect 13173 31433 13185 31436
rect 13219 31433 13231 31467
rect 13173 31427 13231 31433
rect 14458 31424 14464 31476
rect 14516 31464 14522 31476
rect 15013 31467 15071 31473
rect 15013 31464 15025 31467
rect 14516 31436 15025 31464
rect 14516 31424 14522 31436
rect 15013 31433 15025 31436
rect 15059 31433 15071 31467
rect 15013 31427 15071 31433
rect 20993 31467 21051 31473
rect 20993 31433 21005 31467
rect 21039 31464 21051 31467
rect 23382 31464 23388 31476
rect 21039 31436 23388 31464
rect 21039 31433 21051 31436
rect 20993 31427 21051 31433
rect 8006 31368 8156 31396
rect 8220 31368 16436 31396
rect 8006 31365 8018 31368
rect 7960 31359 8018 31365
rect 5373 31331 5431 31337
rect 5373 31297 5385 31331
rect 5419 31328 5431 31331
rect 6822 31328 6828 31340
rect 5419 31300 6828 31328
rect 5419 31297 5431 31300
rect 5373 31291 5431 31297
rect 6822 31288 6828 31300
rect 6880 31288 6886 31340
rect 8220 31337 8248 31368
rect 8205 31331 8263 31337
rect 8205 31297 8217 31331
rect 8251 31297 8263 31331
rect 8205 31291 8263 31297
rect 9973 31331 10031 31337
rect 9973 31297 9985 31331
rect 10019 31328 10031 31331
rect 10134 31328 10140 31340
rect 10019 31300 10140 31328
rect 10019 31297 10031 31300
rect 9973 31291 10031 31297
rect 10134 31288 10140 31300
rect 10192 31288 10198 31340
rect 10244 31337 10272 31368
rect 10229 31331 10287 31337
rect 10229 31297 10241 31331
rect 10275 31297 10287 31331
rect 10229 31291 10287 31297
rect 12825 31331 12883 31337
rect 12825 31297 12837 31331
rect 12871 31328 12883 31331
rect 12986 31328 12992 31340
rect 12871 31300 12992 31328
rect 12871 31297 12883 31300
rect 12825 31291 12883 31297
rect 12986 31288 12992 31300
rect 13044 31288 13050 31340
rect 13096 31272 13124 31368
rect 14297 31331 14355 31337
rect 14297 31297 14309 31331
rect 14343 31328 14355 31331
rect 14458 31328 14464 31340
rect 14343 31300 14464 31328
rect 14343 31297 14355 31300
rect 14297 31291 14355 31297
rect 14458 31288 14464 31300
rect 14516 31288 14522 31340
rect 14568 31337 14596 31368
rect 14553 31331 14611 31337
rect 14553 31297 14565 31331
rect 14599 31297 14611 31331
rect 14553 31291 14611 31297
rect 16137 31331 16195 31337
rect 16137 31297 16149 31331
rect 16183 31328 16195 31331
rect 16298 31328 16304 31340
rect 16183 31300 16304 31328
rect 16183 31297 16195 31300
rect 16137 31291 16195 31297
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 16408 31337 16436 31368
rect 18156 31368 20300 31396
rect 18156 31340 18184 31368
rect 20272 31340 20300 31368
rect 16393 31331 16451 31337
rect 16393 31297 16405 31331
rect 16439 31297 16451 31331
rect 16393 31291 16451 31297
rect 17793 31331 17851 31337
rect 17793 31297 17805 31331
rect 17839 31328 17851 31331
rect 17954 31328 17960 31340
rect 17839 31300 17960 31328
rect 17839 31297 17851 31300
rect 17793 31291 17851 31297
rect 17954 31288 17960 31300
rect 18012 31288 18018 31340
rect 18049 31331 18107 31337
rect 18049 31297 18061 31331
rect 18095 31328 18107 31331
rect 18138 31328 18144 31340
rect 18095 31300 18144 31328
rect 18095 31297 18107 31300
rect 18049 31291 18107 31297
rect 18138 31288 18144 31300
rect 18196 31288 18202 31340
rect 20001 31331 20059 31337
rect 20001 31297 20013 31331
rect 20047 31328 20059 31331
rect 20047 31300 20208 31328
rect 20047 31297 20059 31300
rect 20001 31291 20059 31297
rect 5629 31263 5687 31269
rect 5629 31229 5641 31263
rect 5675 31229 5687 31263
rect 5629 31223 5687 31229
rect 8757 31263 8815 31269
rect 8757 31229 8769 31263
rect 8803 31260 8815 31263
rect 8938 31260 8944 31272
rect 8803 31232 8944 31260
rect 8803 31229 8815 31232
rect 8757 31223 8815 31229
rect 3881 31195 3939 31201
rect 3881 31161 3893 31195
rect 3927 31161 3939 31195
rect 3881 31155 3939 31161
rect 5442 31084 5448 31136
rect 5500 31124 5506 31136
rect 5644 31124 5672 31223
rect 8938 31220 8944 31232
rect 8996 31220 9002 31272
rect 11330 31220 11336 31272
rect 11388 31220 11394 31272
rect 13078 31220 13084 31272
rect 13136 31220 13142 31272
rect 18690 31220 18696 31272
rect 18748 31220 18754 31272
rect 20180 31260 20208 31300
rect 20254 31288 20260 31340
rect 20312 31288 20318 31340
rect 21008 31328 21036 31427
rect 23382 31424 23388 31436
rect 23440 31424 23446 31476
rect 26697 31467 26755 31473
rect 26697 31433 26709 31467
rect 26743 31464 26755 31467
rect 28994 31464 29000 31476
rect 26743 31436 29000 31464
rect 26743 31433 26755 31436
rect 26697 31427 26755 31433
rect 28994 31424 29000 31436
rect 29052 31424 29058 31476
rect 30926 31396 30932 31408
rect 23492 31368 25084 31396
rect 20732 31300 21036 31328
rect 20349 31263 20407 31269
rect 20349 31260 20361 31263
rect 20180 31232 20361 31260
rect 20349 31229 20361 31232
rect 20395 31229 20407 31263
rect 20349 31223 20407 31229
rect 5905 31195 5963 31201
rect 5905 31161 5917 31195
rect 5951 31192 5963 31195
rect 6270 31192 6276 31204
rect 5951 31164 6276 31192
rect 5951 31161 5963 31164
rect 5905 31155 5963 31161
rect 6270 31152 6276 31164
rect 6328 31152 6334 31204
rect 8294 31152 8300 31204
rect 8352 31192 8358 31204
rect 8389 31195 8447 31201
rect 8389 31192 8401 31195
rect 8352 31164 8401 31192
rect 8352 31152 8358 31164
rect 8389 31161 8401 31164
rect 8435 31161 8447 31195
rect 8389 31155 8447 31161
rect 20533 31195 20591 31201
rect 20533 31161 20545 31195
rect 20579 31192 20591 31195
rect 20732 31192 20760 31300
rect 22922 31288 22928 31340
rect 22980 31328 22986 31340
rect 23210 31331 23268 31337
rect 23210 31328 23222 31331
rect 22980 31300 23222 31328
rect 22980 31288 22986 31300
rect 23210 31297 23222 31300
rect 23256 31297 23268 31331
rect 23210 31291 23268 31297
rect 23382 31288 23388 31340
rect 23440 31328 23446 31340
rect 23492 31337 23520 31368
rect 23477 31331 23535 31337
rect 23477 31328 23489 31331
rect 23440 31300 23489 31328
rect 23440 31288 23446 31300
rect 23477 31297 23489 31300
rect 23523 31297 23535 31331
rect 23477 31291 23535 31297
rect 24785 31331 24843 31337
rect 24785 31297 24797 31331
rect 24831 31328 24843 31331
rect 24946 31328 24952 31340
rect 24831 31300 24952 31328
rect 24831 31297 24843 31300
rect 24785 31291 24843 31297
rect 24946 31288 24952 31300
rect 25004 31288 25010 31340
rect 25056 31337 25084 31368
rect 28368 31368 30932 31396
rect 25041 31331 25099 31337
rect 25041 31297 25053 31331
rect 25087 31328 25099 31331
rect 25317 31331 25375 31337
rect 25317 31328 25329 31331
rect 25087 31300 25329 31328
rect 25087 31297 25099 31300
rect 25041 31291 25099 31297
rect 25317 31297 25329 31300
rect 25363 31328 25375 31331
rect 25406 31328 25412 31340
rect 25363 31300 25412 31328
rect 25363 31297 25375 31300
rect 25317 31291 25375 31297
rect 25406 31288 25412 31300
rect 25464 31288 25470 31340
rect 25584 31331 25642 31337
rect 25584 31297 25596 31331
rect 25630 31328 25642 31331
rect 26326 31328 26332 31340
rect 25630 31300 26332 31328
rect 25630 31297 25642 31300
rect 25584 31291 25642 31297
rect 26326 31288 26332 31300
rect 26384 31288 26390 31340
rect 28097 31331 28155 31337
rect 28097 31297 28109 31331
rect 28143 31328 28155 31331
rect 28258 31328 28264 31340
rect 28143 31300 28264 31328
rect 28143 31297 28155 31300
rect 28097 31291 28155 31297
rect 28258 31288 28264 31300
rect 28316 31288 28322 31340
rect 28368 31337 28396 31368
rect 30926 31356 30932 31368
rect 30984 31396 30990 31408
rect 30984 31368 31340 31396
rect 30984 31356 30990 31368
rect 28353 31331 28411 31337
rect 28353 31297 28365 31331
rect 28399 31297 28411 31331
rect 28353 31291 28411 31297
rect 28442 31288 28448 31340
rect 28500 31328 28506 31340
rect 28537 31331 28595 31337
rect 28537 31328 28549 31331
rect 28500 31300 28549 31328
rect 28500 31288 28506 31300
rect 28537 31297 28549 31300
rect 28583 31297 28595 31331
rect 28537 31291 28595 31297
rect 29086 31288 29092 31340
rect 29144 31288 29150 31340
rect 29270 31288 29276 31340
rect 29328 31328 29334 31340
rect 31312 31337 31340 31368
rect 31846 31356 31852 31408
rect 31904 31356 31910 31408
rect 31030 31331 31088 31337
rect 31030 31328 31042 31331
rect 29328 31300 31042 31328
rect 29328 31288 29334 31300
rect 31030 31297 31042 31300
rect 31076 31297 31088 31331
rect 31030 31291 31088 31297
rect 31297 31331 31355 31337
rect 31297 31297 31309 31331
rect 31343 31297 31355 31331
rect 31297 31291 31355 31297
rect 31570 31288 31576 31340
rect 31628 31328 31634 31340
rect 32217 31331 32275 31337
rect 32217 31328 32229 31331
rect 31628 31300 32229 31328
rect 31628 31288 31634 31300
rect 32217 31297 32229 31300
rect 32263 31297 32275 31331
rect 32217 31291 32275 31297
rect 20809 31263 20867 31269
rect 20809 31229 20821 31263
rect 20855 31229 20867 31263
rect 20809 31223 20867 31229
rect 20579 31164 20760 31192
rect 20824 31192 20852 31223
rect 21266 31220 21272 31272
rect 21324 31220 21330 31272
rect 21637 31263 21695 31269
rect 21637 31229 21649 31263
rect 21683 31260 21695 31263
rect 21910 31260 21916 31272
rect 21683 31232 21916 31260
rect 21683 31229 21695 31232
rect 21637 31223 21695 31229
rect 21910 31220 21916 31232
rect 21968 31220 21974 31272
rect 31846 31220 31852 31272
rect 31904 31260 31910 31272
rect 32493 31263 32551 31269
rect 32493 31260 32505 31263
rect 31904 31232 32505 31260
rect 31904 31220 31910 31232
rect 32493 31229 32505 31232
rect 32539 31229 32551 31263
rect 32493 31223 32551 31229
rect 21284 31192 21312 31220
rect 20824 31164 21312 31192
rect 20579 31161 20591 31164
rect 20533 31155 20591 31161
rect 31478 31152 31484 31204
rect 31536 31152 31542 31204
rect 5500 31096 5672 31124
rect 5500 31084 5506 31096
rect 5718 31084 5724 31136
rect 5776 31084 5782 31136
rect 6825 31127 6883 31133
rect 6825 31093 6837 31127
rect 6871 31124 6883 31127
rect 7834 31124 7840 31136
rect 6871 31096 7840 31124
rect 6871 31093 6883 31096
rect 6825 31087 6883 31093
rect 7834 31084 7840 31096
rect 7892 31084 7898 31136
rect 8849 31127 8907 31133
rect 8849 31093 8861 31127
rect 8895 31124 8907 31127
rect 10410 31124 10416 31136
rect 8895 31096 10416 31124
rect 8895 31093 8907 31096
rect 8849 31087 8907 31093
rect 10410 31084 10416 31096
rect 10468 31084 10474 31136
rect 10686 31084 10692 31136
rect 10744 31084 10750 31136
rect 11701 31127 11759 31133
rect 11701 31093 11713 31127
rect 11747 31124 11759 31127
rect 12434 31124 12440 31136
rect 11747 31096 12440 31124
rect 11747 31093 11759 31096
rect 11701 31087 11759 31093
rect 12434 31084 12440 31096
rect 12492 31084 12498 31136
rect 16666 31084 16672 31136
rect 16724 31084 16730 31136
rect 17678 31084 17684 31136
rect 17736 31124 17742 31136
rect 18141 31127 18199 31133
rect 18141 31124 18153 31127
rect 17736 31096 18153 31124
rect 17736 31084 17742 31096
rect 18141 31093 18153 31096
rect 18187 31093 18199 31127
rect 18141 31087 18199 31093
rect 18874 31084 18880 31136
rect 18932 31084 18938 31136
rect 22094 31084 22100 31136
rect 22152 31084 22158 31136
rect 23658 31084 23664 31136
rect 23716 31084 23722 31136
rect 26970 31084 26976 31136
rect 27028 31084 27034 31136
rect 29086 31084 29092 31136
rect 29144 31124 29150 31136
rect 29917 31127 29975 31133
rect 29917 31124 29929 31127
rect 29144 31096 29929 31124
rect 29144 31084 29150 31096
rect 29917 31093 29929 31096
rect 29963 31093 29975 31127
rect 29917 31087 29975 31093
rect 31389 31127 31447 31133
rect 31389 31093 31401 31127
rect 31435 31124 31447 31127
rect 32122 31124 32128 31136
rect 31435 31096 32128 31124
rect 31435 31093 31447 31096
rect 31389 31087 31447 31093
rect 32122 31084 32128 31096
rect 32180 31084 32186 31136
rect 1104 31034 33856 31056
rect 1104 30982 5044 31034
rect 5096 30982 5108 31034
rect 5160 30982 5172 31034
rect 5224 30982 5236 31034
rect 5288 30982 5300 31034
rect 5352 30982 13232 31034
rect 13284 30982 13296 31034
rect 13348 30982 13360 31034
rect 13412 30982 13424 31034
rect 13476 30982 13488 31034
rect 13540 30982 21420 31034
rect 21472 30982 21484 31034
rect 21536 30982 21548 31034
rect 21600 30982 21612 31034
rect 21664 30982 21676 31034
rect 21728 30982 29608 31034
rect 29660 30982 29672 31034
rect 29724 30982 29736 31034
rect 29788 30982 29800 31034
rect 29852 30982 29864 31034
rect 29916 30982 33856 31034
rect 1104 30960 33856 30982
rect 12342 30880 12348 30932
rect 12400 30880 12406 30932
rect 16666 30880 16672 30932
rect 16724 30880 16730 30932
rect 17129 30923 17187 30929
rect 17129 30889 17141 30923
rect 17175 30920 17187 30923
rect 18690 30920 18696 30932
rect 17175 30892 18696 30920
rect 17175 30889 17187 30892
rect 17129 30883 17187 30889
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 18874 30880 18880 30932
rect 18932 30880 18938 30932
rect 20254 30880 20260 30932
rect 20312 30880 20318 30932
rect 21910 30880 21916 30932
rect 21968 30880 21974 30932
rect 22094 30880 22100 30932
rect 22152 30920 22158 30932
rect 22152 30892 22876 30920
rect 22152 30880 22158 30892
rect 14550 30812 14556 30864
rect 14608 30852 14614 30864
rect 15565 30855 15623 30861
rect 15565 30852 15577 30855
rect 14608 30824 15577 30852
rect 14608 30812 14614 30824
rect 15565 30821 15577 30824
rect 15611 30821 15623 30855
rect 15565 30815 15623 30821
rect 5442 30784 5448 30796
rect 3160 30756 5448 30784
rect 1762 30676 1768 30728
rect 1820 30716 1826 30728
rect 3160 30716 3188 30756
rect 5442 30744 5448 30756
rect 5500 30784 5506 30796
rect 5537 30787 5595 30793
rect 5537 30784 5549 30787
rect 5500 30756 5549 30784
rect 5500 30744 5506 30756
rect 5537 30753 5549 30756
rect 5583 30753 5595 30787
rect 5537 30747 5595 30753
rect 7466 30744 7472 30796
rect 7524 30744 7530 30796
rect 8846 30744 8852 30796
rect 8904 30784 8910 30796
rect 9861 30787 9919 30793
rect 9861 30784 9873 30787
rect 8904 30756 9873 30784
rect 8904 30744 8910 30756
rect 9861 30753 9873 30756
rect 9907 30753 9919 30787
rect 9861 30747 9919 30753
rect 12253 30787 12311 30793
rect 12253 30753 12265 30787
rect 12299 30784 12311 30787
rect 12299 30756 13124 30784
rect 12299 30753 12311 30756
rect 12253 30747 12311 30753
rect 13096 30728 13124 30756
rect 16114 30744 16120 30796
rect 16172 30744 16178 30796
rect 16577 30787 16635 30793
rect 16577 30753 16589 30787
rect 16623 30784 16635 30787
rect 16684 30784 16712 30880
rect 16623 30756 16712 30784
rect 16623 30753 16635 30756
rect 16577 30747 16635 30753
rect 17034 30744 17040 30796
rect 17092 30784 17098 30796
rect 17681 30787 17739 30793
rect 17681 30784 17693 30787
rect 17092 30756 17693 30784
rect 17092 30744 17098 30756
rect 17681 30753 17693 30756
rect 17727 30753 17739 30787
rect 18892 30784 18920 30880
rect 19245 30787 19303 30793
rect 19245 30784 19257 30787
rect 18892 30756 19257 30784
rect 17681 30747 17739 30753
rect 19245 30753 19257 30756
rect 19291 30753 19303 30787
rect 20272 30784 20300 30880
rect 21729 30855 21787 30861
rect 21729 30821 21741 30855
rect 21775 30852 21787 30855
rect 21775 30824 22094 30852
rect 21775 30821 21787 30824
rect 21729 30815 21787 30821
rect 20349 30787 20407 30793
rect 20349 30784 20361 30787
rect 20272 30756 20361 30784
rect 19245 30747 19303 30753
rect 20349 30753 20361 30756
rect 20395 30753 20407 30787
rect 22066 30784 22094 30824
rect 22848 30793 22876 30892
rect 23658 30880 23664 30932
rect 23716 30880 23722 30932
rect 24946 30880 24952 30932
rect 25004 30920 25010 30932
rect 25869 30923 25927 30929
rect 25869 30920 25881 30923
rect 25004 30892 25881 30920
rect 25004 30880 25010 30892
rect 25869 30889 25881 30892
rect 25915 30889 25927 30923
rect 25869 30883 25927 30889
rect 26418 30880 26424 30932
rect 26476 30880 26482 30932
rect 33042 30920 33048 30932
rect 31404 30892 33048 30920
rect 23676 30793 23704 30880
rect 26053 30855 26111 30861
rect 26053 30821 26065 30855
rect 26099 30852 26111 30855
rect 26234 30852 26240 30864
rect 26099 30824 26240 30852
rect 26099 30821 26111 30824
rect 26053 30815 26111 30821
rect 26234 30812 26240 30824
rect 26292 30812 26298 30864
rect 22465 30787 22523 30793
rect 22465 30784 22477 30787
rect 22066 30756 22477 30784
rect 20349 30747 20407 30753
rect 22465 30753 22477 30756
rect 22511 30753 22523 30787
rect 22465 30747 22523 30753
rect 22833 30787 22891 30793
rect 22833 30753 22845 30787
rect 22879 30753 22891 30787
rect 22833 30747 22891 30753
rect 23661 30787 23719 30793
rect 23661 30753 23673 30787
rect 23707 30753 23719 30787
rect 26436 30784 26464 30880
rect 31404 30796 31432 30892
rect 33042 30880 33048 30892
rect 33100 30920 33106 30932
rect 33137 30923 33195 30929
rect 33137 30920 33149 30923
rect 33100 30892 33149 30920
rect 33100 30880 33106 30892
rect 33137 30889 33149 30892
rect 33183 30889 33195 30923
rect 33137 30883 33195 30889
rect 23661 30747 23719 30753
rect 24826 30756 26464 30784
rect 1820 30688 3188 30716
rect 5077 30719 5135 30725
rect 1820 30676 1826 30688
rect 5077 30685 5089 30719
rect 5123 30716 5135 30719
rect 5626 30716 5632 30728
rect 5123 30688 5632 30716
rect 5123 30685 5135 30688
rect 5077 30679 5135 30685
rect 5626 30676 5632 30688
rect 5684 30676 5690 30728
rect 5804 30719 5862 30725
rect 5804 30685 5816 30719
rect 5850 30685 5862 30719
rect 5804 30679 5862 30685
rect 2032 30651 2090 30657
rect 2032 30617 2044 30651
rect 2078 30648 2090 30651
rect 4154 30648 4160 30660
rect 2078 30620 4160 30648
rect 2078 30617 2090 30620
rect 2032 30611 2090 30617
rect 4154 30608 4160 30620
rect 4212 30608 4218 30660
rect 4709 30651 4767 30657
rect 4709 30617 4721 30651
rect 4755 30648 4767 30651
rect 5534 30648 5540 30660
rect 4755 30620 5540 30648
rect 4755 30617 4767 30620
rect 4709 30611 4767 30617
rect 5534 30608 5540 30620
rect 5592 30608 5598 30660
rect 5718 30608 5724 30660
rect 5776 30648 5782 30660
rect 5828 30648 5856 30679
rect 8018 30676 8024 30728
rect 8076 30676 8082 30728
rect 8386 30676 8392 30728
rect 8444 30716 8450 30728
rect 9401 30719 9459 30725
rect 9401 30716 9413 30719
rect 8444 30688 9413 30716
rect 8444 30676 8450 30688
rect 9401 30685 9413 30688
rect 9447 30685 9459 30719
rect 9401 30679 9459 30685
rect 11054 30676 11060 30728
rect 11112 30716 11118 30728
rect 11986 30719 12044 30725
rect 11986 30716 11998 30719
rect 11112 30688 11998 30716
rect 11112 30676 11118 30688
rect 11986 30685 11998 30688
rect 12032 30685 12044 30719
rect 11986 30679 12044 30685
rect 12894 30676 12900 30728
rect 12952 30676 12958 30728
rect 13078 30676 13084 30728
rect 13136 30676 13142 30728
rect 13357 30719 13415 30725
rect 13357 30685 13369 30719
rect 13403 30716 13415 30719
rect 13722 30716 13728 30728
rect 13403 30688 13728 30716
rect 13403 30685 13415 30688
rect 13357 30679 13415 30685
rect 13722 30676 13728 30688
rect 13780 30676 13786 30728
rect 13909 30719 13967 30725
rect 13909 30685 13921 30719
rect 13955 30716 13967 30719
rect 14185 30719 14243 30725
rect 14185 30716 14197 30719
rect 13955 30688 14197 30716
rect 13955 30685 13967 30688
rect 13909 30679 13967 30685
rect 14185 30685 14197 30688
rect 14231 30685 14243 30719
rect 14185 30679 14243 30685
rect 14274 30676 14280 30728
rect 14332 30716 14338 30728
rect 14553 30719 14611 30725
rect 14553 30716 14565 30719
rect 14332 30688 14565 30716
rect 14332 30676 14338 30688
rect 14553 30685 14565 30688
rect 14599 30685 14611 30719
rect 14553 30679 14611 30685
rect 17218 30676 17224 30728
rect 17276 30676 17282 30728
rect 19889 30719 19947 30725
rect 19889 30685 19901 30719
rect 19935 30716 19947 30719
rect 20898 30716 20904 30728
rect 19935 30688 20904 30716
rect 19935 30685 19947 30688
rect 19889 30679 19947 30685
rect 20898 30676 20904 30688
rect 20956 30676 20962 30728
rect 23477 30719 23535 30725
rect 23477 30685 23489 30719
rect 23523 30716 23535 30719
rect 24826 30716 24854 30756
rect 27430 30744 27436 30796
rect 27488 30744 27494 30796
rect 28353 30787 28411 30793
rect 28353 30784 28365 30787
rect 27908 30756 28365 30784
rect 23523 30688 24854 30716
rect 25777 30719 25835 30725
rect 23523 30685 23535 30688
rect 23477 30679 23535 30685
rect 25777 30685 25789 30719
rect 25823 30716 25835 30719
rect 26510 30716 26516 30728
rect 25823 30688 26516 30716
rect 25823 30685 25835 30688
rect 25777 30679 25835 30685
rect 26510 30676 26516 30688
rect 26568 30676 26574 30728
rect 27908 30725 27936 30756
rect 28353 30753 28365 30756
rect 28399 30753 28411 30787
rect 28353 30747 28411 30753
rect 30926 30744 30932 30796
rect 30984 30744 30990 30796
rect 31386 30744 31392 30796
rect 31444 30744 31450 30796
rect 27893 30719 27951 30725
rect 27893 30685 27905 30719
rect 27939 30685 27951 30719
rect 27893 30679 27951 30685
rect 28074 30676 28080 30728
rect 28132 30676 28138 30728
rect 30944 30716 30972 30744
rect 32401 30719 32459 30725
rect 32401 30716 32413 30719
rect 30944 30688 31754 30716
rect 5776 30620 5856 30648
rect 20616 30651 20674 30657
rect 5776 30608 5782 30620
rect 20616 30617 20628 30651
rect 20662 30648 20674 30651
rect 21174 30648 21180 30660
rect 20662 30620 21180 30648
rect 20662 30617 20674 30620
rect 20616 30611 20674 30617
rect 21174 30608 21180 30620
rect 21232 30608 21238 30660
rect 23290 30608 23296 30660
rect 23348 30648 23354 30660
rect 24581 30651 24639 30657
rect 24581 30648 24593 30651
rect 23348 30620 24593 30648
rect 23348 30608 23354 30620
rect 24581 30617 24593 30620
rect 24627 30617 24639 30651
rect 24581 30611 24639 30617
rect 25314 30608 25320 30660
rect 25372 30648 25378 30660
rect 26329 30651 26387 30657
rect 26329 30648 26341 30651
rect 25372 30620 26341 30648
rect 25372 30608 25378 30620
rect 26329 30617 26341 30620
rect 26375 30648 26387 30651
rect 27154 30648 27160 30660
rect 26375 30620 27160 30648
rect 26375 30617 26387 30620
rect 26329 30611 26387 30617
rect 27154 30608 27160 30620
rect 27212 30648 27218 30660
rect 27430 30648 27436 30660
rect 27212 30620 27436 30648
rect 27212 30608 27218 30620
rect 27430 30608 27436 30620
rect 27488 30608 27494 30660
rect 28902 30608 28908 30660
rect 28960 30648 28966 30660
rect 30662 30651 30720 30657
rect 30662 30648 30674 30651
rect 28960 30620 30674 30648
rect 28960 30608 28966 30620
rect 30662 30617 30674 30620
rect 30708 30617 30720 30651
rect 31726 30648 31754 30688
rect 32048 30688 32413 30716
rect 32048 30660 32076 30688
rect 32401 30685 32413 30688
rect 32447 30685 32459 30719
rect 32401 30679 32459 30685
rect 32493 30719 32551 30725
rect 32493 30685 32505 30719
rect 32539 30685 32551 30719
rect 32493 30679 32551 30685
rect 32030 30648 32036 30660
rect 31726 30620 32036 30648
rect 30662 30611 30720 30617
rect 32030 30608 32036 30620
rect 32088 30608 32094 30660
rect 32122 30608 32128 30660
rect 32180 30657 32186 30660
rect 32180 30611 32192 30657
rect 32180 30608 32186 30611
rect 3145 30583 3203 30589
rect 3145 30549 3157 30583
rect 3191 30580 3203 30583
rect 4614 30580 4620 30592
rect 3191 30552 4620 30580
rect 3191 30549 3203 30552
rect 3145 30543 3203 30549
rect 4614 30540 4620 30552
rect 4672 30540 4678 30592
rect 6914 30540 6920 30592
rect 6972 30540 6978 30592
rect 8938 30540 8944 30592
rect 8996 30580 9002 30592
rect 9125 30583 9183 30589
rect 9125 30580 9137 30583
rect 8996 30552 9137 30580
rect 8996 30540 9002 30552
rect 9125 30549 9137 30552
rect 9171 30549 9183 30583
rect 9125 30543 9183 30549
rect 10870 30540 10876 30592
rect 10928 30540 10934 30592
rect 24213 30583 24271 30589
rect 24213 30549 24225 30583
rect 24259 30580 24271 30583
rect 25406 30580 25412 30592
rect 24259 30552 25412 30580
rect 24259 30549 24271 30552
rect 24213 30543 24271 30549
rect 25406 30540 25412 30552
rect 25464 30540 25470 30592
rect 26694 30540 26700 30592
rect 26752 30580 26758 30592
rect 29549 30583 29607 30589
rect 29549 30580 29561 30583
rect 26752 30552 29561 30580
rect 26752 30540 26758 30552
rect 29549 30549 29561 30552
rect 29595 30549 29607 30583
rect 29549 30543 29607 30549
rect 30466 30540 30472 30592
rect 30524 30580 30530 30592
rect 31021 30583 31079 30589
rect 31021 30580 31033 30583
rect 30524 30552 31033 30580
rect 30524 30540 30530 30552
rect 31021 30549 31033 30552
rect 31067 30549 31079 30583
rect 31021 30543 31079 30549
rect 31110 30540 31116 30592
rect 31168 30580 31174 30592
rect 32508 30580 32536 30679
rect 31168 30552 32536 30580
rect 31168 30540 31174 30552
rect 1104 30490 34016 30512
rect 1104 30438 9138 30490
rect 9190 30438 9202 30490
rect 9254 30438 9266 30490
rect 9318 30438 9330 30490
rect 9382 30438 9394 30490
rect 9446 30438 17326 30490
rect 17378 30438 17390 30490
rect 17442 30438 17454 30490
rect 17506 30438 17518 30490
rect 17570 30438 17582 30490
rect 17634 30438 25514 30490
rect 25566 30438 25578 30490
rect 25630 30438 25642 30490
rect 25694 30438 25706 30490
rect 25758 30438 25770 30490
rect 25822 30438 33702 30490
rect 33754 30438 33766 30490
rect 33818 30438 33830 30490
rect 33882 30438 33894 30490
rect 33946 30438 33958 30490
rect 34010 30438 34016 30490
rect 1104 30416 34016 30438
rect 2498 30336 2504 30388
rect 2556 30376 2562 30388
rect 2556 30348 3096 30376
rect 2556 30336 2562 30348
rect 2317 30311 2375 30317
rect 2317 30277 2329 30311
rect 2363 30308 2375 30311
rect 2590 30308 2596 30320
rect 2363 30280 2596 30308
rect 2363 30277 2375 30280
rect 2317 30271 2375 30277
rect 2590 30268 2596 30280
rect 2648 30268 2654 30320
rect 3068 30317 3096 30348
rect 6822 30336 6828 30388
rect 6880 30336 6886 30388
rect 8294 30336 8300 30388
rect 8352 30336 8358 30388
rect 11330 30336 11336 30388
rect 11388 30336 11394 30388
rect 12986 30336 12992 30388
rect 13044 30376 13050 30388
rect 13081 30379 13139 30385
rect 13081 30376 13093 30379
rect 13044 30348 13093 30376
rect 13044 30336 13050 30348
rect 13081 30345 13093 30348
rect 13127 30345 13139 30379
rect 13081 30339 13139 30345
rect 13722 30336 13728 30388
rect 13780 30336 13786 30388
rect 14458 30336 14464 30388
rect 14516 30336 14522 30388
rect 16298 30336 16304 30388
rect 16356 30336 16362 30388
rect 17954 30336 17960 30388
rect 18012 30376 18018 30388
rect 18141 30379 18199 30385
rect 18141 30376 18153 30379
rect 18012 30348 18153 30376
rect 18012 30336 18018 30348
rect 18141 30345 18153 30348
rect 18187 30345 18199 30379
rect 18141 30339 18199 30345
rect 21174 30336 21180 30388
rect 21232 30336 21238 30388
rect 22462 30336 22468 30388
rect 22520 30376 22526 30388
rect 23382 30376 23388 30388
rect 22520 30348 23388 30376
rect 22520 30336 22526 30348
rect 23382 30336 23388 30348
rect 23440 30336 23446 30388
rect 26513 30379 26571 30385
rect 26513 30345 26525 30379
rect 26559 30376 26571 30379
rect 27614 30376 27620 30388
rect 26559 30348 27620 30376
rect 26559 30345 26571 30348
rect 26513 30339 26571 30345
rect 27614 30336 27620 30348
rect 27672 30336 27678 30388
rect 28166 30336 28172 30388
rect 28224 30376 28230 30388
rect 28224 30348 31432 30376
rect 28224 30336 28230 30348
rect 3053 30311 3111 30317
rect 3053 30277 3065 30311
rect 3099 30277 3111 30311
rect 4525 30311 4583 30317
rect 4525 30308 4537 30311
rect 3053 30271 3111 30277
rect 3160 30280 4537 30308
rect 2685 30243 2743 30249
rect 2685 30209 2697 30243
rect 2731 30240 2743 30243
rect 2958 30240 2964 30252
rect 2731 30212 2964 30240
rect 2731 30209 2743 30212
rect 2685 30203 2743 30209
rect 2958 30200 2964 30212
rect 3016 30200 3022 30252
rect 1026 30132 1032 30184
rect 1084 30172 1090 30184
rect 3160 30172 3188 30280
rect 4525 30277 4537 30280
rect 4571 30277 4583 30311
rect 4525 30271 4583 30277
rect 6178 30268 6184 30320
rect 6236 30308 6242 30320
rect 6362 30308 6368 30320
rect 6236 30280 6368 30308
rect 6236 30268 6242 30280
rect 6362 30268 6368 30280
rect 6420 30268 6426 30320
rect 4249 30243 4307 30249
rect 4249 30209 4261 30243
rect 4295 30240 4307 30243
rect 4295 30212 4568 30240
rect 4295 30209 4307 30212
rect 4249 30203 4307 30209
rect 1084 30144 3188 30172
rect 1084 30132 1090 30144
rect 4540 30048 4568 30212
rect 5534 30200 5540 30252
rect 5592 30200 5598 30252
rect 6914 30200 6920 30252
rect 6972 30240 6978 30252
rect 7009 30243 7067 30249
rect 7009 30240 7021 30243
rect 6972 30212 7021 30240
rect 6972 30200 6978 30212
rect 7009 30209 7021 30212
rect 7055 30209 7067 30243
rect 8312 30240 8340 30336
rect 8662 30268 8668 30320
rect 8720 30308 8726 30320
rect 9125 30311 9183 30317
rect 9125 30308 9137 30311
rect 8720 30280 9137 30308
rect 8720 30268 8726 30280
rect 9125 30277 9137 30280
rect 9171 30277 9183 30311
rect 9125 30271 9183 30277
rect 9858 30268 9864 30320
rect 9916 30308 9922 30320
rect 11885 30311 11943 30317
rect 11885 30308 11897 30311
rect 9916 30280 11897 30308
rect 9916 30268 9922 30280
rect 11885 30277 11897 30280
rect 11931 30277 11943 30311
rect 11885 30271 11943 30277
rect 24670 30268 24676 30320
rect 24728 30308 24734 30320
rect 24765 30311 24823 30317
rect 24765 30308 24777 30311
rect 24728 30280 24777 30308
rect 24728 30268 24734 30280
rect 24765 30277 24777 30280
rect 24811 30277 24823 30311
rect 31294 30308 31300 30320
rect 24765 30271 24823 30277
rect 28552 30280 31300 30308
rect 9677 30243 9735 30249
rect 9677 30240 9689 30243
rect 8312 30212 9689 30240
rect 7009 30203 7067 30209
rect 9677 30209 9689 30212
rect 9723 30209 9735 30243
rect 9677 30203 9735 30209
rect 10410 30200 10416 30252
rect 10468 30200 10474 30252
rect 10781 30243 10839 30249
rect 10781 30209 10793 30243
rect 10827 30240 10839 30243
rect 10870 30240 10876 30252
rect 10827 30212 10876 30240
rect 10827 30209 10839 30212
rect 10781 30203 10839 30209
rect 10870 30200 10876 30212
rect 10928 30200 10934 30252
rect 12434 30200 12440 30252
rect 12492 30200 12498 30252
rect 12621 30243 12679 30249
rect 12621 30209 12633 30243
rect 12667 30240 12679 30243
rect 13449 30243 13507 30249
rect 13449 30240 13461 30243
rect 12667 30212 13461 30240
rect 12667 30209 12679 30212
rect 12621 30203 12679 30209
rect 13449 30209 13461 30212
rect 13495 30240 13507 30243
rect 18601 30243 18659 30249
rect 13495 30212 14964 30240
rect 13495 30209 13507 30212
rect 13449 30203 13507 30209
rect 7653 30175 7711 30181
rect 7653 30141 7665 30175
rect 7699 30172 7711 30175
rect 8297 30175 8355 30181
rect 8297 30172 8309 30175
rect 7699 30144 8309 30172
rect 7699 30141 7711 30144
rect 7653 30135 7711 30141
rect 8297 30141 8309 30144
rect 8343 30141 8355 30175
rect 8297 30135 8355 30141
rect 11146 30132 11152 30184
rect 11204 30172 11210 30184
rect 12636 30172 12664 30203
rect 14936 30181 14964 30212
rect 18601 30209 18613 30243
rect 18647 30240 18659 30243
rect 18969 30243 19027 30249
rect 18969 30240 18981 30243
rect 18647 30212 18981 30240
rect 18647 30209 18659 30212
rect 18601 30203 18659 30209
rect 18969 30209 18981 30212
rect 19015 30240 19027 30243
rect 21266 30240 21272 30252
rect 19015 30212 21272 30240
rect 19015 30209 19027 30212
rect 18969 30203 19027 30209
rect 21266 30200 21272 30212
rect 21324 30240 21330 30252
rect 21637 30243 21695 30249
rect 21637 30240 21649 30243
rect 21324 30212 21649 30240
rect 21324 30200 21330 30212
rect 21637 30209 21649 30212
rect 21683 30240 21695 30243
rect 21683 30212 22140 30240
rect 21683 30209 21695 30212
rect 21637 30203 21695 30209
rect 11204 30144 12664 30172
rect 14277 30175 14335 30181
rect 11204 30132 11210 30144
rect 14277 30141 14289 30175
rect 14323 30141 14335 30175
rect 14277 30135 14335 30141
rect 14921 30175 14979 30181
rect 14921 30141 14933 30175
rect 14967 30172 14979 30175
rect 15841 30175 15899 30181
rect 15841 30172 15853 30175
rect 14967 30144 15332 30172
rect 14967 30141 14979 30144
rect 14921 30135 14979 30141
rect 6733 30107 6791 30113
rect 6733 30104 6745 30107
rect 6656 30076 6745 30104
rect 6656 30048 6684 30076
rect 6733 30073 6745 30076
rect 6779 30104 6791 30107
rect 7745 30107 7803 30113
rect 7745 30104 7757 30107
rect 6779 30076 7757 30104
rect 6779 30073 6791 30076
rect 6733 30067 6791 30073
rect 7745 30073 7757 30076
rect 7791 30073 7803 30107
rect 7745 30067 7803 30073
rect 9674 30064 9680 30116
rect 9732 30104 9738 30116
rect 9861 30107 9919 30113
rect 9861 30104 9873 30107
rect 9732 30076 9873 30104
rect 9732 30064 9738 30076
rect 9861 30073 9873 30076
rect 9907 30073 9919 30107
rect 9861 30067 9919 30073
rect 12989 30107 13047 30113
rect 12989 30073 13001 30107
rect 13035 30104 13047 30107
rect 13722 30104 13728 30116
rect 13035 30076 13728 30104
rect 13035 30073 13047 30076
rect 12989 30067 13047 30073
rect 13722 30064 13728 30076
rect 13780 30064 13786 30116
rect 4522 29996 4528 30048
rect 4580 29996 4586 30048
rect 6638 29996 6644 30048
rect 6696 29996 6702 30048
rect 13630 29996 13636 30048
rect 13688 30036 13694 30048
rect 14292 30036 14320 30135
rect 14550 30064 14556 30116
rect 14608 30064 14614 30116
rect 15304 30045 15332 30144
rect 15764 30144 15853 30172
rect 15764 30048 15792 30144
rect 15841 30141 15853 30144
rect 15887 30141 15899 30175
rect 15841 30135 15899 30141
rect 22002 30132 22008 30184
rect 22060 30132 22066 30184
rect 22112 30181 22140 30212
rect 25406 30200 25412 30252
rect 25464 30200 25470 30252
rect 22097 30175 22155 30181
rect 22097 30141 22109 30175
rect 22143 30172 22155 30175
rect 23385 30175 23443 30181
rect 23385 30172 23397 30175
rect 22143 30144 23397 30172
rect 22143 30141 22155 30144
rect 22097 30135 22155 30141
rect 23385 30141 23397 30144
rect 23431 30172 23443 30175
rect 23566 30172 23572 30184
rect 23431 30144 23572 30172
rect 23431 30141 23443 30144
rect 23385 30135 23443 30141
rect 23566 30132 23572 30144
rect 23624 30132 23630 30184
rect 24213 30175 24271 30181
rect 24213 30172 24225 30175
rect 23768 30144 24225 30172
rect 16209 30107 16267 30113
rect 16209 30073 16221 30107
rect 16255 30104 16267 30107
rect 17678 30104 17684 30116
rect 16255 30076 17684 30104
rect 16255 30073 16267 30076
rect 16209 30067 16267 30073
rect 17678 30064 17684 30076
rect 17736 30064 17742 30116
rect 18325 30107 18383 30113
rect 18325 30073 18337 30107
rect 18371 30104 18383 30107
rect 18506 30104 18512 30116
rect 18371 30076 18512 30104
rect 18371 30073 18383 30076
rect 18325 30067 18383 30073
rect 18506 30064 18512 30076
rect 18564 30064 18570 30116
rect 21361 30107 21419 30113
rect 21361 30073 21373 30107
rect 21407 30104 21419 30107
rect 22020 30104 22048 30132
rect 21407 30076 22048 30104
rect 21407 30073 21419 30076
rect 21361 30067 21419 30073
rect 22922 30064 22928 30116
rect 22980 30064 22986 30116
rect 23109 30107 23167 30113
rect 23109 30073 23121 30107
rect 23155 30104 23167 30107
rect 23768 30104 23796 30144
rect 24213 30141 24225 30144
rect 24259 30172 24271 30175
rect 24857 30175 24915 30181
rect 24857 30172 24869 30175
rect 24259 30144 24869 30172
rect 24259 30141 24271 30144
rect 24213 30135 24271 30141
rect 24857 30141 24869 30144
rect 24903 30141 24915 30175
rect 24857 30135 24915 30141
rect 25961 30175 26019 30181
rect 25961 30141 25973 30175
rect 26007 30172 26019 30175
rect 26234 30172 26240 30184
rect 26007 30144 26240 30172
rect 26007 30141 26019 30144
rect 25961 30135 26019 30141
rect 26234 30132 26240 30144
rect 26292 30132 26298 30184
rect 26326 30132 26332 30184
rect 26384 30172 26390 30184
rect 26973 30175 27031 30181
rect 26973 30172 26985 30175
rect 26384 30144 26985 30172
rect 26384 30132 26390 30144
rect 26973 30141 26985 30144
rect 27019 30141 27031 30175
rect 26973 30135 27031 30141
rect 27430 30132 27436 30184
rect 27488 30172 27494 30184
rect 27982 30172 27988 30184
rect 27488 30144 27988 30172
rect 27488 30132 27494 30144
rect 27982 30132 27988 30144
rect 28040 30132 28046 30184
rect 28552 30181 28580 30280
rect 31294 30268 31300 30280
rect 31352 30268 31358 30320
rect 31404 30308 31432 30348
rect 32370 30311 32428 30317
rect 32370 30308 32382 30311
rect 31404 30280 32382 30308
rect 32370 30277 32382 30280
rect 32416 30277 32428 30311
rect 32370 30271 32428 30277
rect 28994 30200 29000 30252
rect 29052 30200 29058 30252
rect 29733 30243 29791 30249
rect 29733 30209 29745 30243
rect 29779 30240 29791 30243
rect 30006 30240 30012 30252
rect 29779 30212 30012 30240
rect 29779 30209 29791 30212
rect 29733 30203 29791 30209
rect 30006 30200 30012 30212
rect 30064 30200 30070 30252
rect 30098 30200 30104 30252
rect 30156 30240 30162 30252
rect 30653 30243 30711 30249
rect 30653 30240 30665 30243
rect 30156 30212 30665 30240
rect 30156 30200 30162 30212
rect 30653 30209 30665 30212
rect 30699 30209 30711 30243
rect 30653 30203 30711 30209
rect 28537 30175 28595 30181
rect 28537 30141 28549 30175
rect 28583 30141 28595 30175
rect 28537 30135 28595 30141
rect 29178 30132 29184 30184
rect 29236 30132 29242 30184
rect 30926 30132 30932 30184
rect 30984 30132 30990 30184
rect 32122 30132 32128 30184
rect 32180 30132 32186 30184
rect 23155 30076 23796 30104
rect 23937 30107 23995 30113
rect 23155 30073 23167 30076
rect 23109 30067 23167 30073
rect 23937 30073 23949 30107
rect 23983 30104 23995 30107
rect 24946 30104 24952 30116
rect 23983 30076 24952 30104
rect 23983 30073 23995 30076
rect 23937 30067 23995 30073
rect 24946 30064 24952 30076
rect 25004 30064 25010 30116
rect 27157 30107 27215 30113
rect 27157 30073 27169 30107
rect 27203 30104 27215 30107
rect 27338 30104 27344 30116
rect 27203 30076 27344 30104
rect 27203 30073 27215 30076
rect 27157 30067 27215 30073
rect 27338 30064 27344 30076
rect 27396 30104 27402 30116
rect 31018 30104 31024 30116
rect 27396 30076 31024 30104
rect 27396 30064 27402 30076
rect 31018 30064 31024 30076
rect 31076 30064 31082 30116
rect 13688 30008 14320 30036
rect 15289 30039 15347 30045
rect 13688 29996 13694 30008
rect 15289 30005 15301 30039
rect 15335 30036 15347 30039
rect 15746 30036 15752 30048
rect 15335 30008 15752 30036
rect 15335 30005 15347 30008
rect 15289 29999 15347 30005
rect 15746 29996 15752 30008
rect 15804 29996 15810 30048
rect 24029 30039 24087 30045
rect 24029 30005 24041 30039
rect 24075 30036 24087 30039
rect 29270 30036 29276 30048
rect 24075 30008 29276 30036
rect 24075 30005 24087 30008
rect 24029 29999 24087 30005
rect 29270 29996 29276 30008
rect 29328 29996 29334 30048
rect 29362 29996 29368 30048
rect 29420 30036 29426 30048
rect 30101 30039 30159 30045
rect 30101 30036 30113 30039
rect 29420 30008 30113 30036
rect 29420 29996 29426 30008
rect 30101 30005 30113 30008
rect 30147 30036 30159 30039
rect 30190 30036 30196 30048
rect 30147 30008 30196 30036
rect 30147 30005 30159 30008
rect 30101 29999 30159 30005
rect 30190 29996 30196 30008
rect 30248 29996 30254 30048
rect 33502 29996 33508 30048
rect 33560 29996 33566 30048
rect 1104 29946 33856 29968
rect 1104 29894 5044 29946
rect 5096 29894 5108 29946
rect 5160 29894 5172 29946
rect 5224 29894 5236 29946
rect 5288 29894 5300 29946
rect 5352 29894 13232 29946
rect 13284 29894 13296 29946
rect 13348 29894 13360 29946
rect 13412 29894 13424 29946
rect 13476 29894 13488 29946
rect 13540 29894 21420 29946
rect 21472 29894 21484 29946
rect 21536 29894 21548 29946
rect 21600 29894 21612 29946
rect 21664 29894 21676 29946
rect 21728 29894 29608 29946
rect 29660 29894 29672 29946
rect 29724 29894 29736 29946
rect 29788 29894 29800 29946
rect 29852 29894 29864 29946
rect 29916 29894 33856 29946
rect 1104 29872 33856 29894
rect 4154 29792 4160 29844
rect 4212 29832 4218 29844
rect 5997 29835 6055 29841
rect 5997 29832 6009 29835
rect 4212 29804 6009 29832
rect 4212 29792 4218 29804
rect 5997 29801 6009 29804
rect 6043 29801 6055 29835
rect 5997 29795 6055 29801
rect 7006 29792 7012 29844
rect 7064 29792 7070 29844
rect 7098 29792 7104 29844
rect 7156 29832 7162 29844
rect 7193 29835 7251 29841
rect 7193 29832 7205 29835
rect 7156 29804 7205 29832
rect 7156 29792 7162 29804
rect 7193 29801 7205 29804
rect 7239 29801 7251 29835
rect 7193 29795 7251 29801
rect 10134 29792 10140 29844
rect 10192 29832 10198 29844
rect 10321 29835 10379 29841
rect 10321 29832 10333 29835
rect 10192 29804 10333 29832
rect 10192 29792 10198 29804
rect 10321 29801 10333 29804
rect 10367 29801 10379 29835
rect 10321 29795 10379 29801
rect 10962 29792 10968 29844
rect 11020 29832 11026 29844
rect 11241 29835 11299 29841
rect 11241 29832 11253 29835
rect 11020 29804 11253 29832
rect 11020 29792 11026 29804
rect 11241 29801 11253 29804
rect 11287 29801 11299 29835
rect 11241 29795 11299 29801
rect 26234 29792 26240 29844
rect 26292 29792 26298 29844
rect 27893 29835 27951 29841
rect 27893 29801 27905 29835
rect 27939 29832 27951 29835
rect 28442 29832 28448 29844
rect 27939 29804 28448 29832
rect 27939 29801 27951 29804
rect 27893 29795 27951 29801
rect 28442 29792 28448 29804
rect 28500 29792 28506 29844
rect 6178 29724 6184 29776
rect 6236 29724 6242 29776
rect 7024 29764 7052 29792
rect 7285 29767 7343 29773
rect 7285 29764 7297 29767
rect 7024 29736 7297 29764
rect 7285 29733 7297 29736
rect 7331 29733 7343 29767
rect 7285 29727 7343 29733
rect 10505 29767 10563 29773
rect 10505 29733 10517 29767
rect 10551 29764 10563 29767
rect 10686 29764 10692 29776
rect 10551 29736 10692 29764
rect 10551 29733 10563 29736
rect 10505 29727 10563 29733
rect 10686 29724 10692 29736
rect 10744 29764 10750 29776
rect 10744 29736 11836 29764
rect 10744 29724 10750 29736
rect 3418 29696 3424 29708
rect 2700 29668 3424 29696
rect 2700 29637 2728 29668
rect 3418 29656 3424 29668
rect 3476 29656 3482 29708
rect 4522 29656 4528 29708
rect 4580 29656 4586 29708
rect 4614 29656 4620 29708
rect 4672 29696 4678 29708
rect 5261 29699 5319 29705
rect 5261 29696 5273 29699
rect 4672 29668 5273 29696
rect 4672 29656 4678 29668
rect 5261 29665 5273 29668
rect 5307 29665 5319 29699
rect 5261 29659 5319 29665
rect 6362 29656 6368 29708
rect 6420 29696 6426 29708
rect 6457 29699 6515 29705
rect 6457 29696 6469 29699
rect 6420 29668 6469 29696
rect 6420 29656 6426 29668
rect 6457 29665 6469 29668
rect 6503 29665 6515 29699
rect 6457 29659 6515 29665
rect 6638 29656 6644 29708
rect 6696 29656 6702 29708
rect 7834 29656 7840 29708
rect 7892 29656 7898 29708
rect 8938 29656 8944 29708
rect 8996 29696 9002 29708
rect 10781 29699 10839 29705
rect 10781 29696 10793 29699
rect 8996 29668 10793 29696
rect 8996 29656 9002 29668
rect 10781 29665 10793 29668
rect 10827 29696 10839 29699
rect 11146 29696 11152 29708
rect 10827 29668 11152 29696
rect 10827 29665 10839 29668
rect 10781 29659 10839 29665
rect 11146 29656 11152 29668
rect 11204 29656 11210 29708
rect 11808 29705 11836 29736
rect 28258 29724 28264 29776
rect 28316 29764 28322 29776
rect 29549 29767 29607 29773
rect 29549 29764 29561 29767
rect 28316 29736 29561 29764
rect 28316 29724 28322 29736
rect 29549 29733 29561 29736
rect 29595 29733 29607 29767
rect 29549 29727 29607 29733
rect 29733 29767 29791 29773
rect 29733 29733 29745 29767
rect 29779 29764 29791 29767
rect 31386 29764 31392 29776
rect 29779 29736 31392 29764
rect 29779 29733 29791 29736
rect 29733 29727 29791 29733
rect 31386 29724 31392 29736
rect 31444 29724 31450 29776
rect 11793 29699 11851 29705
rect 11793 29665 11805 29699
rect 11839 29665 11851 29699
rect 11793 29659 11851 29665
rect 24854 29656 24860 29708
rect 24912 29656 24918 29708
rect 25409 29699 25467 29705
rect 25409 29665 25421 29699
rect 25455 29696 25467 29699
rect 25455 29668 28120 29696
rect 25455 29665 25467 29668
rect 25409 29659 25467 29665
rect 2685 29631 2743 29637
rect 2685 29597 2697 29631
rect 2731 29597 2743 29631
rect 2685 29591 2743 29597
rect 2961 29631 3019 29637
rect 2961 29597 2973 29631
rect 3007 29628 3019 29631
rect 4246 29628 4252 29640
rect 3007 29600 4252 29628
rect 3007 29597 3019 29600
rect 2961 29591 3019 29597
rect 4246 29588 4252 29600
rect 4304 29588 4310 29640
rect 4890 29588 4896 29640
rect 4948 29628 4954 29640
rect 5077 29631 5135 29637
rect 5077 29628 5089 29631
rect 4948 29600 5089 29628
rect 4948 29588 4954 29600
rect 5077 29597 5089 29600
rect 5123 29597 5135 29631
rect 5077 29591 5135 29597
rect 23566 29588 23572 29640
rect 23624 29628 23630 29640
rect 24213 29631 24271 29637
rect 24213 29628 24225 29631
rect 23624 29600 24225 29628
rect 23624 29588 23630 29600
rect 24213 29597 24225 29600
rect 24259 29628 24271 29631
rect 25314 29628 25320 29640
rect 24259 29600 25320 29628
rect 24259 29597 24271 29600
rect 24213 29591 24271 29597
rect 25314 29588 25320 29600
rect 25372 29588 25378 29640
rect 25593 29631 25651 29637
rect 25593 29597 25605 29631
rect 25639 29628 25651 29631
rect 26694 29628 26700 29640
rect 25639 29600 26700 29628
rect 25639 29597 25651 29600
rect 25593 29591 25651 29597
rect 26694 29588 26700 29600
rect 26752 29588 26758 29640
rect 26878 29588 26884 29640
rect 26936 29588 26942 29640
rect 27338 29588 27344 29640
rect 27396 29588 27402 29640
rect 28092 29637 28120 29668
rect 28994 29656 29000 29708
rect 29052 29696 29058 29708
rect 30561 29699 30619 29705
rect 30561 29696 30573 29699
rect 29052 29668 30573 29696
rect 29052 29656 29058 29668
rect 30561 29665 30573 29668
rect 30607 29665 30619 29699
rect 30561 29659 30619 29665
rect 28077 29631 28135 29637
rect 28077 29597 28089 29631
rect 28123 29597 28135 29631
rect 28077 29591 28135 29597
rect 30282 29588 30288 29640
rect 30340 29588 30346 29640
rect 31665 29631 31723 29637
rect 30760 29600 31064 29628
rect 2317 29563 2375 29569
rect 2317 29529 2329 29563
rect 2363 29560 2375 29563
rect 2363 29532 2912 29560
rect 2363 29529 2375 29532
rect 2317 29523 2375 29529
rect 2884 29504 2912 29532
rect 28626 29520 28632 29572
rect 28684 29520 28690 29572
rect 28718 29520 28724 29572
rect 28776 29560 28782 29572
rect 29362 29560 29368 29572
rect 28776 29532 29368 29560
rect 28776 29520 28782 29532
rect 29362 29520 29368 29532
rect 29420 29560 29426 29572
rect 30009 29563 30067 29569
rect 30009 29560 30021 29563
rect 29420 29532 30021 29560
rect 29420 29520 29426 29532
rect 30009 29529 30021 29532
rect 30055 29529 30067 29563
rect 30009 29523 30067 29529
rect 30190 29520 30196 29572
rect 30248 29560 30254 29572
rect 30760 29560 30788 29600
rect 30248 29532 30788 29560
rect 31036 29560 31064 29600
rect 31665 29597 31677 29631
rect 31711 29628 31723 29631
rect 31711 29600 32168 29628
rect 31711 29597 31723 29600
rect 31665 29591 31723 29597
rect 32140 29572 32168 29600
rect 31910 29563 31968 29569
rect 31910 29560 31922 29563
rect 31036 29532 31922 29560
rect 30248 29520 30254 29532
rect 31910 29529 31922 29532
rect 31956 29529 31968 29563
rect 31910 29523 31968 29529
rect 32122 29520 32128 29572
rect 32180 29520 32186 29572
rect 2866 29452 2872 29504
rect 2924 29452 2930 29504
rect 3510 29452 3516 29504
rect 3568 29452 3574 29504
rect 5902 29452 5908 29504
rect 5960 29452 5966 29504
rect 26145 29495 26203 29501
rect 26145 29461 26157 29495
rect 26191 29492 26203 29495
rect 29270 29492 29276 29504
rect 26191 29464 29276 29492
rect 26191 29461 26203 29464
rect 26145 29455 26203 29461
rect 29270 29452 29276 29464
rect 29328 29452 29334 29504
rect 29454 29452 29460 29504
rect 29512 29492 29518 29504
rect 33045 29495 33103 29501
rect 33045 29492 33057 29495
rect 29512 29464 33057 29492
rect 29512 29452 29518 29464
rect 33045 29461 33057 29464
rect 33091 29461 33103 29495
rect 33045 29455 33103 29461
rect 1104 29402 34016 29424
rect 1104 29350 9138 29402
rect 9190 29350 9202 29402
rect 9254 29350 9266 29402
rect 9318 29350 9330 29402
rect 9382 29350 9394 29402
rect 9446 29350 17326 29402
rect 17378 29350 17390 29402
rect 17442 29350 17454 29402
rect 17506 29350 17518 29402
rect 17570 29350 17582 29402
rect 17634 29350 25514 29402
rect 25566 29350 25578 29402
rect 25630 29350 25642 29402
rect 25694 29350 25706 29402
rect 25758 29350 25770 29402
rect 25822 29350 33702 29402
rect 33754 29350 33766 29402
rect 33818 29350 33830 29402
rect 33882 29350 33894 29402
rect 33946 29350 33958 29402
rect 34010 29350 34016 29402
rect 1104 29328 34016 29350
rect 7653 29291 7711 29297
rect 7653 29257 7665 29291
rect 7699 29288 7711 29291
rect 8018 29288 8024 29300
rect 7699 29260 8024 29288
rect 7699 29257 7711 29260
rect 7653 29251 7711 29257
rect 8018 29248 8024 29260
rect 8076 29248 8082 29300
rect 26053 29291 26111 29297
rect 26053 29257 26065 29291
rect 26099 29288 26111 29291
rect 28074 29288 28080 29300
rect 26099 29260 28080 29288
rect 26099 29257 26111 29260
rect 26053 29251 26111 29257
rect 28074 29248 28080 29260
rect 28132 29248 28138 29300
rect 28997 29291 29055 29297
rect 28997 29257 29009 29291
rect 29043 29288 29055 29291
rect 31110 29288 31116 29300
rect 29043 29260 31116 29288
rect 29043 29257 29055 29260
rect 28997 29251 29055 29257
rect 31110 29248 31116 29260
rect 31168 29248 31174 29300
rect 30285 29223 30343 29229
rect 2700 29192 3648 29220
rect 2700 29161 2728 29192
rect 3620 29164 3648 29192
rect 30285 29189 30297 29223
rect 30331 29220 30343 29223
rect 32950 29220 32956 29232
rect 30331 29192 32956 29220
rect 30331 29189 30343 29192
rect 30285 29183 30343 29189
rect 32950 29180 32956 29192
rect 33008 29180 33014 29232
rect 2685 29155 2743 29161
rect 2685 29121 2697 29155
rect 2731 29121 2743 29155
rect 2685 29115 2743 29121
rect 2866 29112 2872 29164
rect 2924 29112 2930 29164
rect 3602 29112 3608 29164
rect 3660 29112 3666 29164
rect 4430 29112 4436 29164
rect 4488 29112 4494 29164
rect 6270 29112 6276 29164
rect 6328 29152 6334 29164
rect 7009 29155 7067 29161
rect 7009 29152 7021 29155
rect 6328 29124 7021 29152
rect 6328 29112 6334 29124
rect 7009 29121 7021 29124
rect 7055 29121 7067 29155
rect 7009 29115 7067 29121
rect 26970 29112 26976 29164
rect 27028 29152 27034 29164
rect 27249 29155 27307 29161
rect 27249 29152 27261 29155
rect 27028 29124 27261 29152
rect 27028 29112 27034 29124
rect 27249 29121 27261 29124
rect 27295 29121 27307 29155
rect 27249 29115 27307 29121
rect 28445 29155 28503 29161
rect 28445 29121 28457 29155
rect 28491 29152 28503 29155
rect 29086 29152 29092 29164
rect 28491 29124 29092 29152
rect 28491 29121 28503 29124
rect 28445 29115 28503 29121
rect 29086 29112 29092 29124
rect 29144 29112 29150 29164
rect 29178 29112 29184 29164
rect 29236 29112 29242 29164
rect 31938 29112 31944 29164
rect 31996 29112 32002 29164
rect 32381 29155 32439 29161
rect 32381 29152 32393 29155
rect 32048 29124 32393 29152
rect 2133 29087 2191 29093
rect 2133 29053 2145 29087
rect 2179 29084 2191 29087
rect 2774 29084 2780 29096
rect 2179 29056 2780 29084
rect 2179 29053 2191 29056
rect 2133 29047 2191 29053
rect 2774 29044 2780 29056
rect 2832 29044 2838 29096
rect 3326 29044 3332 29096
rect 3384 29044 3390 29096
rect 4338 29044 4344 29096
rect 4396 29084 4402 29096
rect 4801 29087 4859 29093
rect 4801 29084 4813 29087
rect 4396 29056 4813 29084
rect 4396 29044 4402 29056
rect 4801 29053 4813 29056
rect 4847 29053 4859 29087
rect 4801 29047 4859 29053
rect 25501 29087 25559 29093
rect 25501 29053 25513 29087
rect 25547 29084 25559 29087
rect 25547 29056 26188 29084
rect 25547 29053 25559 29056
rect 25501 29047 25559 29053
rect 26160 28957 26188 29056
rect 26786 29044 26792 29096
rect 26844 29044 26850 29096
rect 27893 29087 27951 29093
rect 27893 29053 27905 29087
rect 27939 29084 27951 29087
rect 30374 29084 30380 29096
rect 27939 29056 30380 29084
rect 27939 29053 27951 29056
rect 27893 29047 27951 29053
rect 30374 29044 30380 29056
rect 30432 29044 30438 29096
rect 31478 29044 31484 29096
rect 31536 29044 31542 29096
rect 29362 28976 29368 29028
rect 29420 29016 29426 29028
rect 32048 29016 32076 29124
rect 32381 29121 32393 29124
rect 32427 29121 32439 29155
rect 32381 29115 32439 29121
rect 32122 29044 32128 29096
rect 32180 29044 32186 29096
rect 29420 28988 32076 29016
rect 29420 28976 29426 28988
rect 26145 28951 26203 28957
rect 26145 28917 26157 28951
rect 26191 28948 26203 28951
rect 27154 28948 27160 28960
rect 26191 28920 27160 28948
rect 26191 28917 26203 28920
rect 26145 28911 26203 28917
rect 27154 28908 27160 28920
rect 27212 28908 27218 28960
rect 28074 28908 28080 28960
rect 28132 28948 28138 28960
rect 28169 28951 28227 28957
rect 28169 28948 28181 28951
rect 28132 28920 28181 28948
rect 28132 28908 28138 28920
rect 28169 28917 28181 28920
rect 28215 28948 28227 28951
rect 28718 28948 28724 28960
rect 28215 28920 28724 28948
rect 28215 28917 28227 28920
rect 28169 28911 28227 28917
rect 28718 28908 28724 28920
rect 28776 28908 28782 28960
rect 30742 28908 30748 28960
rect 30800 28948 30806 28960
rect 33505 28951 33563 28957
rect 33505 28948 33517 28951
rect 30800 28920 33517 28948
rect 30800 28908 30806 28920
rect 33505 28917 33517 28920
rect 33551 28917 33563 28951
rect 33505 28911 33563 28917
rect 1104 28858 33856 28880
rect 1104 28806 5044 28858
rect 5096 28806 5108 28858
rect 5160 28806 5172 28858
rect 5224 28806 5236 28858
rect 5288 28806 5300 28858
rect 5352 28806 13232 28858
rect 13284 28806 13296 28858
rect 13348 28806 13360 28858
rect 13412 28806 13424 28858
rect 13476 28806 13488 28858
rect 13540 28806 21420 28858
rect 21472 28806 21484 28858
rect 21536 28806 21548 28858
rect 21600 28806 21612 28858
rect 21664 28806 21676 28858
rect 21728 28806 29608 28858
rect 29660 28806 29672 28858
rect 29724 28806 29736 28858
rect 29788 28806 29800 28858
rect 29852 28806 29864 28858
rect 29916 28806 33856 28858
rect 1104 28784 33856 28806
rect 29365 28747 29423 28753
rect 29365 28713 29377 28747
rect 29411 28744 29423 28747
rect 31570 28744 31576 28756
rect 29411 28716 31576 28744
rect 29411 28713 29423 28716
rect 29365 28707 29423 28713
rect 31570 28704 31576 28716
rect 31628 28704 31634 28756
rect 33502 28676 33508 28688
rect 25884 28648 33508 28676
rect 4430 28568 4436 28620
rect 4488 28568 4494 28620
rect 5902 28568 5908 28620
rect 5960 28568 5966 28620
rect 5994 28568 6000 28620
rect 6052 28568 6058 28620
rect 25884 28617 25912 28648
rect 33502 28636 33508 28648
rect 33560 28636 33566 28688
rect 25869 28611 25927 28617
rect 25869 28577 25881 28611
rect 25915 28577 25927 28611
rect 25869 28571 25927 28577
rect 27341 28611 27399 28617
rect 27341 28577 27353 28611
rect 27387 28608 27399 28611
rect 30742 28608 30748 28620
rect 27387 28580 30748 28608
rect 27387 28577 27399 28580
rect 27341 28571 27399 28577
rect 30742 28568 30748 28580
rect 30800 28568 30806 28620
rect 30834 28568 30840 28620
rect 30892 28568 30898 28620
rect 31938 28568 31944 28620
rect 31996 28608 32002 28620
rect 32493 28611 32551 28617
rect 32493 28608 32505 28611
rect 31996 28580 32505 28608
rect 31996 28568 32002 28580
rect 32493 28577 32505 28580
rect 32539 28577 32551 28611
rect 32493 28571 32551 28577
rect 2685 28543 2743 28549
rect 2685 28509 2697 28543
rect 2731 28509 2743 28543
rect 2685 28503 2743 28509
rect 2317 28475 2375 28481
rect 2317 28441 2329 28475
rect 2363 28472 2375 28475
rect 2700 28472 2728 28503
rect 2958 28500 2964 28552
rect 3016 28500 3022 28552
rect 3878 28500 3884 28552
rect 3936 28500 3942 28552
rect 6641 28543 6699 28549
rect 6641 28509 6653 28543
rect 6687 28540 6699 28543
rect 7285 28543 7343 28549
rect 7285 28540 7297 28543
rect 6687 28512 7297 28540
rect 6687 28509 6699 28512
rect 6641 28503 6699 28509
rect 7285 28509 7297 28512
rect 7331 28509 7343 28543
rect 7285 28503 7343 28509
rect 9585 28543 9643 28549
rect 9585 28509 9597 28543
rect 9631 28540 9643 28543
rect 10410 28540 10416 28552
rect 9631 28512 10416 28540
rect 9631 28509 9643 28512
rect 9585 28503 9643 28509
rect 10410 28500 10416 28512
rect 10468 28500 10474 28552
rect 24946 28500 24952 28552
rect 25004 28500 25010 28552
rect 26421 28543 26479 28549
rect 26421 28509 26433 28543
rect 26467 28540 26479 28543
rect 26513 28543 26571 28549
rect 26513 28540 26525 28543
rect 26467 28512 26525 28540
rect 26467 28509 26479 28512
rect 26421 28503 26479 28509
rect 26513 28509 26525 28512
rect 26559 28509 26571 28543
rect 26513 28503 26571 28509
rect 27982 28500 27988 28552
rect 28040 28500 28046 28552
rect 28718 28540 28724 28552
rect 28092 28512 28724 28540
rect 3786 28472 3792 28484
rect 2363 28444 2636 28472
rect 2700 28444 3792 28472
rect 2363 28441 2375 28444
rect 2317 28435 2375 28441
rect 2608 28416 2636 28444
rect 3786 28432 3792 28444
rect 3844 28432 3850 28484
rect 24964 28472 24992 28500
rect 28092 28472 28120 28512
rect 28718 28500 28724 28512
rect 28776 28500 28782 28552
rect 30558 28500 30564 28552
rect 30616 28500 30622 28552
rect 31846 28500 31852 28552
rect 31904 28500 31910 28552
rect 32217 28543 32275 28549
rect 32217 28509 32229 28543
rect 32263 28509 32275 28543
rect 32217 28503 32275 28509
rect 24964 28444 28120 28472
rect 28629 28475 28687 28481
rect 28629 28441 28641 28475
rect 28675 28472 28687 28475
rect 32232 28472 32260 28503
rect 28675 28444 32260 28472
rect 28675 28441 28687 28444
rect 28629 28435 28687 28441
rect 2590 28364 2596 28416
rect 2648 28364 2654 28416
rect 3513 28407 3571 28413
rect 3513 28373 3525 28407
rect 3559 28404 3571 28407
rect 4338 28404 4344 28416
rect 3559 28376 4344 28404
rect 3559 28373 3571 28376
rect 3513 28367 3571 28373
rect 4338 28364 4344 28376
rect 4396 28364 4402 28416
rect 4430 28364 4436 28416
rect 4488 28404 4494 28416
rect 5261 28407 5319 28413
rect 5261 28404 5273 28407
rect 4488 28376 5273 28404
rect 4488 28364 4494 28376
rect 5261 28373 5273 28376
rect 5307 28373 5319 28407
rect 5261 28367 5319 28373
rect 5718 28364 5724 28416
rect 5776 28404 5782 28416
rect 6178 28404 6184 28416
rect 5776 28376 6184 28404
rect 5776 28364 5782 28376
rect 6178 28364 6184 28376
rect 6236 28404 6242 28416
rect 6733 28407 6791 28413
rect 6733 28404 6745 28407
rect 6236 28376 6745 28404
rect 6236 28364 6242 28376
rect 6733 28373 6745 28376
rect 6779 28373 6791 28407
rect 6733 28367 6791 28373
rect 7098 28364 7104 28416
rect 7156 28404 7162 28416
rect 8941 28407 8999 28413
rect 8941 28404 8953 28407
rect 7156 28376 8953 28404
rect 7156 28364 7162 28376
rect 8941 28373 8953 28376
rect 8987 28373 8999 28407
rect 8941 28367 8999 28373
rect 27157 28407 27215 28413
rect 27157 28373 27169 28407
rect 27203 28404 27215 28407
rect 27706 28404 27712 28416
rect 27203 28376 27712 28404
rect 27203 28373 27215 28376
rect 27157 28367 27215 28373
rect 27706 28364 27712 28376
rect 27764 28364 27770 28416
rect 27890 28364 27896 28416
rect 27948 28364 27954 28416
rect 29914 28364 29920 28416
rect 29972 28364 29978 28416
rect 1104 28314 34016 28336
rect 1104 28262 9138 28314
rect 9190 28262 9202 28314
rect 9254 28262 9266 28314
rect 9318 28262 9330 28314
rect 9382 28262 9394 28314
rect 9446 28262 17326 28314
rect 17378 28262 17390 28314
rect 17442 28262 17454 28314
rect 17506 28262 17518 28314
rect 17570 28262 17582 28314
rect 17634 28262 25514 28314
rect 25566 28262 25578 28314
rect 25630 28262 25642 28314
rect 25694 28262 25706 28314
rect 25758 28262 25770 28314
rect 25822 28262 33702 28314
rect 33754 28262 33766 28314
rect 33818 28262 33830 28314
rect 33882 28262 33894 28314
rect 33946 28262 33958 28314
rect 34010 28262 34016 28314
rect 1104 28240 34016 28262
rect 4890 28160 4896 28212
rect 4948 28200 4954 28212
rect 5077 28203 5135 28209
rect 5077 28200 5089 28203
rect 4948 28172 5089 28200
rect 4948 28160 4954 28172
rect 5077 28169 5089 28172
rect 5123 28169 5135 28203
rect 5077 28163 5135 28169
rect 26786 28160 26792 28212
rect 26844 28200 26850 28212
rect 27525 28203 27583 28209
rect 27525 28200 27537 28203
rect 26844 28172 27537 28200
rect 26844 28160 26850 28172
rect 27525 28169 27537 28172
rect 27571 28169 27583 28203
rect 27525 28163 27583 28169
rect 29641 28203 29699 28209
rect 29641 28169 29653 28203
rect 29687 28200 29699 28203
rect 30098 28200 30104 28212
rect 29687 28172 30104 28200
rect 29687 28169 29699 28172
rect 29641 28163 29699 28169
rect 30098 28160 30104 28172
rect 30156 28160 30162 28212
rect 30558 28160 30564 28212
rect 30616 28200 30622 28212
rect 33505 28203 33563 28209
rect 33505 28200 33517 28203
rect 30616 28172 33517 28200
rect 30616 28160 30622 28172
rect 33505 28169 33517 28172
rect 33551 28169 33563 28203
rect 33505 28163 33563 28169
rect 3602 28092 3608 28144
rect 3660 28092 3666 28144
rect 32370 28135 32428 28141
rect 32370 28132 32382 28135
rect 27448 28104 32382 28132
rect 2590 28024 2596 28076
rect 2648 28024 2654 28076
rect 4154 28024 4160 28076
rect 4212 28024 4218 28076
rect 5718 28024 5724 28076
rect 5776 28024 5782 28076
rect 1578 27956 1584 28008
rect 1636 27956 1642 28008
rect 4433 27999 4491 28005
rect 4433 27965 4445 27999
rect 4479 27996 4491 27999
rect 4798 27996 4804 28008
rect 4479 27968 4804 27996
rect 4479 27965 4491 27968
rect 4433 27959 4491 27965
rect 4798 27956 4804 27968
rect 4856 27956 4862 28008
rect 27448 28005 27476 28104
rect 32370 28101 32382 28104
rect 32416 28101 32428 28135
rect 32370 28095 32428 28101
rect 27890 28024 27896 28076
rect 27948 28064 27954 28076
rect 28813 28067 28871 28073
rect 28813 28064 28825 28067
rect 27948 28036 28825 28064
rect 27948 28024 27954 28036
rect 28813 28033 28825 28036
rect 28859 28033 28871 28067
rect 29454 28064 29460 28076
rect 28813 28027 28871 28033
rect 28920 28036 29460 28064
rect 26973 27999 27031 28005
rect 26973 27996 26985 27999
rect 26896 27968 26985 27996
rect 26896 27872 26924 27968
rect 26973 27965 26985 27968
rect 27019 27965 27031 27999
rect 26973 27959 27031 27965
rect 27433 27999 27491 28005
rect 27433 27965 27445 27999
rect 27479 27965 27491 27999
rect 27433 27959 27491 27965
rect 28169 27999 28227 28005
rect 28169 27965 28181 27999
rect 28215 27996 28227 27999
rect 28920 27996 28948 28036
rect 29454 28024 29460 28036
rect 29512 28024 29518 28076
rect 29914 28024 29920 28076
rect 29972 28064 29978 28076
rect 30377 28067 30435 28073
rect 30377 28064 30389 28067
rect 29972 28036 30389 28064
rect 29972 28024 29978 28036
rect 30377 28033 30389 28036
rect 30423 28033 30435 28067
rect 30377 28027 30435 28033
rect 31938 28024 31944 28076
rect 31996 28024 32002 28076
rect 28215 27968 28948 27996
rect 29089 27999 29147 28005
rect 28215 27965 28227 27968
rect 28169 27959 28227 27965
rect 29089 27965 29101 27999
rect 29135 27996 29147 27999
rect 29178 27996 29184 28008
rect 29135 27968 29184 27996
rect 29135 27965 29147 27968
rect 29089 27959 29147 27965
rect 29178 27956 29184 27968
rect 29236 27996 29242 28008
rect 31386 27996 31392 28008
rect 29236 27968 31392 27996
rect 29236 27956 29242 27968
rect 31386 27956 31392 27968
rect 31444 27956 31450 28008
rect 31478 27956 31484 28008
rect 31536 27956 31542 28008
rect 31662 27956 31668 28008
rect 31720 27996 31726 28008
rect 32122 27996 32128 28008
rect 31720 27968 32128 27996
rect 31720 27956 31726 27968
rect 32122 27956 32128 27968
rect 32180 27956 32186 28008
rect 27341 27931 27399 27937
rect 27341 27897 27353 27931
rect 27387 27928 27399 27931
rect 27982 27928 27988 27940
rect 27387 27900 27988 27928
rect 27387 27897 27399 27900
rect 27341 27891 27399 27897
rect 27982 27888 27988 27900
rect 28040 27928 28046 27940
rect 28261 27931 28319 27937
rect 28261 27928 28273 27931
rect 28040 27900 28273 27928
rect 28040 27888 28046 27900
rect 28261 27897 28273 27900
rect 28307 27897 28319 27931
rect 28261 27891 28319 27897
rect 4890 27820 4896 27872
rect 4948 27860 4954 27872
rect 4985 27863 5043 27869
rect 4985 27860 4997 27863
rect 4948 27832 4997 27860
rect 4948 27820 4954 27832
rect 4985 27829 4997 27832
rect 5031 27829 5043 27863
rect 4985 27823 5043 27829
rect 26789 27863 26847 27869
rect 26789 27829 26801 27863
rect 26835 27860 26847 27863
rect 26878 27860 26884 27872
rect 26835 27832 26884 27860
rect 26835 27829 26847 27832
rect 26789 27823 26847 27829
rect 26878 27820 26884 27832
rect 26936 27820 26942 27872
rect 29825 27863 29883 27869
rect 29825 27829 29837 27863
rect 29871 27860 29883 27863
rect 30098 27860 30104 27872
rect 29871 27832 30104 27860
rect 29871 27829 29883 27832
rect 29825 27823 29883 27829
rect 30098 27820 30104 27832
rect 30156 27820 30162 27872
rect 1104 27770 33856 27792
rect 1104 27718 5044 27770
rect 5096 27718 5108 27770
rect 5160 27718 5172 27770
rect 5224 27718 5236 27770
rect 5288 27718 5300 27770
rect 5352 27718 13232 27770
rect 13284 27718 13296 27770
rect 13348 27718 13360 27770
rect 13412 27718 13424 27770
rect 13476 27718 13488 27770
rect 13540 27718 21420 27770
rect 21472 27718 21484 27770
rect 21536 27718 21548 27770
rect 21600 27718 21612 27770
rect 21664 27718 21676 27770
rect 21728 27718 29608 27770
rect 29660 27718 29672 27770
rect 29724 27718 29736 27770
rect 29788 27718 29800 27770
rect 29852 27718 29864 27770
rect 29916 27718 33856 27770
rect 1104 27696 33856 27718
rect 2958 27616 2964 27668
rect 3016 27656 3022 27668
rect 3145 27659 3203 27665
rect 3145 27656 3157 27659
rect 3016 27628 3157 27656
rect 3016 27616 3022 27628
rect 3145 27625 3157 27628
rect 3191 27625 3203 27659
rect 3145 27619 3203 27625
rect 3789 27659 3847 27665
rect 3789 27625 3801 27659
rect 3835 27656 3847 27659
rect 3878 27656 3884 27668
rect 3835 27628 3884 27656
rect 3835 27625 3847 27628
rect 3789 27619 3847 27625
rect 3878 27616 3884 27628
rect 3936 27616 3942 27668
rect 4154 27616 4160 27668
rect 4212 27656 4218 27668
rect 4525 27659 4583 27665
rect 4525 27656 4537 27659
rect 4212 27628 4537 27656
rect 4212 27616 4218 27628
rect 4525 27625 4537 27628
rect 4571 27625 4583 27659
rect 4525 27619 4583 27625
rect 4798 27616 4804 27668
rect 4856 27656 4862 27668
rect 5261 27659 5319 27665
rect 5261 27656 5273 27659
rect 4856 27628 5273 27656
rect 4856 27616 4862 27628
rect 5261 27625 5273 27628
rect 5307 27625 5319 27659
rect 27893 27659 27951 27665
rect 5261 27619 5319 27625
rect 24872 27628 27752 27656
rect 24872 27600 24900 27628
rect 24854 27548 24860 27600
rect 24912 27548 24918 27600
rect 27154 27548 27160 27600
rect 27212 27548 27218 27600
rect 27724 27597 27752 27628
rect 27893 27625 27905 27659
rect 27939 27656 27951 27659
rect 28902 27656 28908 27668
rect 27939 27628 28908 27656
rect 27939 27625 27951 27628
rect 27893 27619 27951 27625
rect 28902 27616 28908 27628
rect 28960 27616 28966 27668
rect 30193 27659 30251 27665
rect 30193 27625 30205 27659
rect 30239 27656 30251 27659
rect 30282 27656 30288 27668
rect 30239 27628 30288 27656
rect 30239 27625 30251 27628
rect 30193 27619 30251 27625
rect 30282 27616 30288 27628
rect 30340 27616 30346 27668
rect 27709 27591 27767 27597
rect 27709 27557 27721 27591
rect 27755 27588 27767 27591
rect 28350 27588 28356 27600
rect 27755 27560 28356 27588
rect 27755 27557 27767 27560
rect 27709 27551 27767 27557
rect 28350 27548 28356 27560
rect 28408 27548 28414 27600
rect 30466 27588 30472 27600
rect 28552 27560 30472 27588
rect 4430 27480 4436 27532
rect 4488 27480 4494 27532
rect 4890 27480 4896 27532
rect 4948 27520 4954 27532
rect 5077 27523 5135 27529
rect 5077 27520 5089 27523
rect 4948 27492 5089 27520
rect 4948 27480 4954 27492
rect 5077 27489 5089 27492
rect 5123 27489 5135 27523
rect 5077 27483 5135 27489
rect 27341 27523 27399 27529
rect 27341 27489 27353 27523
rect 27387 27520 27399 27523
rect 28166 27520 28172 27532
rect 27387 27492 28172 27520
rect 27387 27489 27399 27492
rect 27341 27483 27399 27489
rect 28166 27480 28172 27492
rect 28224 27480 28230 27532
rect 28552 27529 28580 27560
rect 30466 27548 30472 27560
rect 30524 27548 30530 27600
rect 32214 27588 32220 27600
rect 31864 27560 32220 27588
rect 31864 27529 31892 27560
rect 32214 27548 32220 27560
rect 32272 27548 32278 27600
rect 28537 27523 28595 27529
rect 28537 27489 28549 27523
rect 28583 27489 28595 27523
rect 31849 27523 31907 27529
rect 28537 27483 28595 27489
rect 28644 27492 30374 27520
rect 28644 27464 28672 27492
rect 1762 27412 1768 27464
rect 1820 27412 1826 27464
rect 5810 27412 5816 27464
rect 5868 27412 5874 27464
rect 28626 27412 28632 27464
rect 28684 27412 28690 27464
rect 28718 27412 28724 27464
rect 28776 27412 28782 27464
rect 29270 27412 29276 27464
rect 29328 27412 29334 27464
rect 29546 27412 29552 27464
rect 29604 27412 29610 27464
rect 30346 27452 30374 27492
rect 31849 27489 31861 27523
rect 31895 27489 31907 27523
rect 31849 27483 31907 27489
rect 31938 27480 31944 27532
rect 31996 27520 32002 27532
rect 32493 27523 32551 27529
rect 32493 27520 32505 27523
rect 31996 27492 32505 27520
rect 31996 27480 32002 27492
rect 32493 27489 32505 27492
rect 32539 27489 32551 27523
rect 32493 27483 32551 27489
rect 30653 27455 30711 27461
rect 30653 27452 30665 27455
rect 30346 27424 30665 27452
rect 30653 27421 30665 27424
rect 30699 27421 30711 27455
rect 30653 27415 30711 27421
rect 32214 27412 32220 27464
rect 32272 27412 32278 27464
rect 2032 27387 2090 27393
rect 2032 27353 2044 27387
rect 2078 27384 2090 27387
rect 3602 27384 3608 27396
rect 2078 27356 3608 27384
rect 2078 27353 2090 27356
rect 2032 27347 2090 27353
rect 3602 27344 3608 27356
rect 3660 27344 3666 27396
rect 26878 27344 26884 27396
rect 26936 27344 26942 27396
rect 27433 27387 27491 27393
rect 27433 27353 27445 27387
rect 27479 27384 27491 27387
rect 28074 27384 28080 27396
rect 27479 27356 28080 27384
rect 27479 27353 27491 27356
rect 27433 27347 27491 27353
rect 28074 27344 28080 27356
rect 28132 27344 28138 27396
rect 27982 27276 27988 27328
rect 28040 27276 28046 27328
rect 1104 27226 34016 27248
rect 1104 27174 9138 27226
rect 9190 27174 9202 27226
rect 9254 27174 9266 27226
rect 9318 27174 9330 27226
rect 9382 27174 9394 27226
rect 9446 27174 17326 27226
rect 17378 27174 17390 27226
rect 17442 27174 17454 27226
rect 17506 27174 17518 27226
rect 17570 27174 17582 27226
rect 17634 27174 25514 27226
rect 25566 27174 25578 27226
rect 25630 27174 25642 27226
rect 25694 27174 25706 27226
rect 25758 27174 25770 27226
rect 25822 27174 33702 27226
rect 33754 27174 33766 27226
rect 33818 27174 33830 27226
rect 33882 27174 33894 27226
rect 33946 27174 33958 27226
rect 34010 27174 34016 27226
rect 1104 27152 34016 27174
rect 3602 27072 3608 27124
rect 3660 27072 3666 27124
rect 4249 27115 4307 27121
rect 4249 27081 4261 27115
rect 4295 27112 4307 27115
rect 5810 27112 5816 27124
rect 4295 27084 5816 27112
rect 4295 27081 4307 27084
rect 4249 27075 4307 27081
rect 5810 27072 5816 27084
rect 5868 27072 5874 27124
rect 10410 27072 10416 27124
rect 10468 27072 10474 27124
rect 28261 27115 28319 27121
rect 28261 27081 28273 27115
rect 28307 27081 28319 27115
rect 28261 27075 28319 27081
rect 3620 27044 3648 27072
rect 5537 27047 5595 27053
rect 3620 27016 5120 27044
rect 1762 26936 1768 26988
rect 1820 26976 1826 26988
rect 2685 26979 2743 26985
rect 1820 26948 2636 26976
rect 1820 26936 1826 26948
rect 2409 26911 2467 26917
rect 2409 26877 2421 26911
rect 2455 26877 2467 26911
rect 2608 26908 2636 26948
rect 2685 26945 2697 26979
rect 2731 26976 2743 26979
rect 2774 26976 2780 26988
rect 2731 26948 2780 26976
rect 2731 26945 2743 26948
rect 2685 26939 2743 26945
rect 2774 26936 2780 26948
rect 2832 26936 2838 26988
rect 3136 26979 3194 26985
rect 3136 26945 3148 26979
rect 3182 26976 3194 26979
rect 4154 26976 4160 26988
rect 3182 26948 4160 26976
rect 3182 26945 3194 26948
rect 3136 26939 3194 26945
rect 4154 26936 4160 26948
rect 4212 26936 4218 26988
rect 4338 26936 4344 26988
rect 4396 26936 4402 26988
rect 5092 26917 5120 27016
rect 5537 27013 5549 27047
rect 5583 27044 5595 27047
rect 5718 27044 5724 27056
rect 5583 27016 5724 27044
rect 5583 27013 5595 27016
rect 5537 27007 5595 27013
rect 5718 27004 5724 27016
rect 5776 27044 5782 27056
rect 6362 27044 6368 27056
rect 5776 27016 6368 27044
rect 5776 27004 5782 27016
rect 6362 27004 6368 27016
rect 6420 27004 6426 27056
rect 28276 27044 28304 27075
rect 28350 27072 28356 27124
rect 28408 27072 28414 27124
rect 29733 27115 29791 27121
rect 29733 27081 29745 27115
rect 29779 27112 29791 27115
rect 30006 27112 30012 27124
rect 29779 27084 30012 27112
rect 29779 27081 29791 27084
rect 29733 27075 29791 27081
rect 30006 27072 30012 27084
rect 30064 27072 30070 27124
rect 30190 27072 30196 27124
rect 30248 27072 30254 27124
rect 30469 27115 30527 27121
rect 30469 27081 30481 27115
rect 30515 27112 30527 27115
rect 32214 27112 32220 27124
rect 30515 27084 32220 27112
rect 30515 27081 30527 27084
rect 30469 27075 30527 27081
rect 32214 27072 32220 27084
rect 32272 27072 32278 27124
rect 30208 27044 30236 27072
rect 28276 27016 30236 27044
rect 31757 27047 31815 27053
rect 31757 27013 31769 27047
rect 31803 27044 31815 27047
rect 33410 27044 33416 27056
rect 31803 27016 33416 27044
rect 31803 27013 31815 27016
rect 31757 27007 31815 27013
rect 33410 27004 33416 27016
rect 33468 27004 33474 27056
rect 5626 26936 5632 26988
rect 5684 26976 5690 26988
rect 6457 26979 6515 26985
rect 6457 26976 6469 26979
rect 5684 26948 6469 26976
rect 5684 26936 5690 26948
rect 6457 26945 6469 26948
rect 6503 26945 6515 26979
rect 6457 26939 6515 26945
rect 7098 26936 7104 26988
rect 7156 26936 7162 26988
rect 27706 26936 27712 26988
rect 27764 26976 27770 26988
rect 27764 26948 27936 26976
rect 27764 26936 27770 26948
rect 2869 26911 2927 26917
rect 2869 26908 2881 26911
rect 2608 26880 2881 26908
rect 2409 26871 2467 26877
rect 2869 26877 2881 26880
rect 2915 26877 2927 26911
rect 2869 26871 2927 26877
rect 5077 26911 5135 26917
rect 5077 26877 5089 26911
rect 5123 26877 5135 26911
rect 5077 26871 5135 26877
rect 11057 26911 11115 26917
rect 11057 26877 11069 26911
rect 11103 26908 11115 26911
rect 12066 26908 12072 26920
rect 11103 26880 12072 26908
rect 11103 26877 11115 26880
rect 11057 26871 11115 26877
rect 2424 26772 2452 26871
rect 12066 26868 12072 26880
rect 12124 26868 12130 26920
rect 26878 26868 26884 26920
rect 26936 26908 26942 26920
rect 27525 26911 27583 26917
rect 27525 26908 27537 26911
rect 26936 26880 27537 26908
rect 26936 26868 26942 26880
rect 27525 26877 27537 26880
rect 27571 26908 27583 26911
rect 27798 26908 27804 26920
rect 27571 26880 27804 26908
rect 27571 26877 27583 26880
rect 27525 26871 27583 26877
rect 27798 26868 27804 26880
rect 27856 26868 27862 26920
rect 27908 26908 27936 26948
rect 27982 26936 27988 26988
rect 28040 26976 28046 26988
rect 28905 26979 28963 26985
rect 28905 26976 28917 26979
rect 28040 26948 28917 26976
rect 28040 26936 28046 26948
rect 28905 26945 28917 26948
rect 28951 26945 28963 26979
rect 28905 26939 28963 26945
rect 29917 26979 29975 26985
rect 29917 26945 29929 26979
rect 29963 26976 29975 26979
rect 30098 26976 30104 26988
rect 29963 26948 30104 26976
rect 29963 26945 29975 26948
rect 29917 26939 29975 26945
rect 30098 26936 30104 26948
rect 30156 26936 30162 26988
rect 30745 26979 30803 26985
rect 30745 26945 30757 26979
rect 30791 26976 30803 26979
rect 30926 26976 30932 26988
rect 30791 26948 30932 26976
rect 30791 26945 30803 26948
rect 30745 26939 30803 26945
rect 30926 26936 30932 26948
rect 30984 26936 30990 26988
rect 32306 26936 32312 26988
rect 32364 26936 32370 26988
rect 29086 26908 29092 26920
rect 27908 26880 29092 26908
rect 29086 26868 29092 26880
rect 29144 26868 29150 26920
rect 33318 26868 33324 26920
rect 33376 26868 33382 26920
rect 4890 26800 4896 26852
rect 4948 26840 4954 26852
rect 5169 26843 5227 26849
rect 5169 26840 5181 26843
rect 4948 26812 5181 26840
rect 4948 26800 4954 26812
rect 5169 26809 5181 26812
rect 5215 26809 5227 26843
rect 5169 26803 5227 26809
rect 27614 26800 27620 26852
rect 27672 26840 27678 26852
rect 28077 26843 28135 26849
rect 28077 26840 28089 26843
rect 27672 26812 28089 26840
rect 27672 26800 27678 26812
rect 28077 26809 28089 26812
rect 28123 26840 28135 26843
rect 29546 26840 29552 26852
rect 28123 26812 29552 26840
rect 28123 26809 28135 26812
rect 28077 26803 28135 26809
rect 29546 26800 29552 26812
rect 29604 26800 29610 26852
rect 2590 26772 2596 26784
rect 2424 26744 2596 26772
rect 2590 26732 2596 26744
rect 2648 26732 2654 26784
rect 4430 26732 4436 26784
rect 4488 26772 4494 26784
rect 4985 26775 5043 26781
rect 4985 26772 4997 26775
rect 4488 26744 4997 26772
rect 4488 26732 4494 26744
rect 4985 26741 4997 26744
rect 5031 26741 5043 26775
rect 4985 26735 5043 26741
rect 1104 26682 33856 26704
rect 1104 26630 5044 26682
rect 5096 26630 5108 26682
rect 5160 26630 5172 26682
rect 5224 26630 5236 26682
rect 5288 26630 5300 26682
rect 5352 26630 13232 26682
rect 13284 26630 13296 26682
rect 13348 26630 13360 26682
rect 13412 26630 13424 26682
rect 13476 26630 13488 26682
rect 13540 26630 21420 26682
rect 21472 26630 21484 26682
rect 21536 26630 21548 26682
rect 21600 26630 21612 26682
rect 21664 26630 21676 26682
rect 21728 26630 29608 26682
rect 29660 26630 29672 26682
rect 29724 26630 29736 26682
rect 29788 26630 29800 26682
rect 29852 26630 29864 26682
rect 29916 26630 33856 26682
rect 1104 26608 33856 26630
rect 3786 26528 3792 26580
rect 3844 26528 3850 26580
rect 4154 26528 4160 26580
rect 4212 26568 4218 26580
rect 5261 26571 5319 26577
rect 5261 26568 5273 26571
rect 4212 26540 5273 26568
rect 4212 26528 4218 26540
rect 5261 26537 5273 26540
rect 5307 26537 5319 26571
rect 5261 26531 5319 26537
rect 29362 26528 29368 26580
rect 29420 26528 29426 26580
rect 4246 26460 4252 26512
rect 4304 26500 4310 26512
rect 4525 26503 4583 26509
rect 4525 26500 4537 26503
rect 4304 26472 4537 26500
rect 4304 26460 4310 26472
rect 4525 26469 4537 26472
rect 4571 26469 4583 26503
rect 4525 26463 4583 26469
rect 5442 26460 5448 26512
rect 5500 26460 5506 26512
rect 29086 26460 29092 26512
rect 29144 26500 29150 26512
rect 29181 26503 29239 26509
rect 29181 26500 29193 26503
rect 29144 26472 29193 26500
rect 29144 26460 29150 26472
rect 29181 26469 29193 26472
rect 29227 26469 29239 26503
rect 29181 26463 29239 26469
rect 30009 26503 30067 26509
rect 30009 26469 30021 26503
rect 30055 26500 30067 26503
rect 30098 26500 30104 26512
rect 30055 26472 30104 26500
rect 30055 26469 30067 26472
rect 30009 26463 30067 26469
rect 30098 26460 30104 26472
rect 30156 26460 30162 26512
rect 2317 26435 2375 26441
rect 2317 26401 2329 26435
rect 2363 26432 2375 26435
rect 2774 26432 2780 26444
rect 2363 26404 2780 26432
rect 2363 26401 2375 26404
rect 2317 26395 2375 26401
rect 2774 26392 2780 26404
rect 2832 26392 2838 26444
rect 4430 26392 4436 26444
rect 4488 26392 4494 26444
rect 5718 26392 5724 26444
rect 5776 26392 5782 26444
rect 28074 26392 28080 26444
rect 28132 26432 28138 26444
rect 30742 26432 30748 26444
rect 28132 26404 30748 26432
rect 28132 26392 28138 26404
rect 30742 26392 30748 26404
rect 30800 26392 30806 26444
rect 2590 26324 2596 26376
rect 2648 26324 2654 26376
rect 2961 26367 3019 26373
rect 2961 26333 2973 26367
rect 3007 26364 3019 26367
rect 3970 26364 3976 26376
rect 3007 26336 3976 26364
rect 3007 26333 3019 26336
rect 2961 26327 3019 26333
rect 3970 26324 3976 26336
rect 4028 26324 4034 26376
rect 4154 26324 4160 26376
rect 4212 26364 4218 26376
rect 5077 26367 5135 26373
rect 5077 26364 5089 26367
rect 4212 26336 5089 26364
rect 4212 26324 4218 26336
rect 5077 26333 5089 26336
rect 5123 26333 5135 26367
rect 5077 26327 5135 26333
rect 18138 26324 18144 26376
rect 18196 26324 18202 26376
rect 30190 26324 30196 26376
rect 30248 26324 30254 26376
rect 30926 26324 30932 26376
rect 30984 26324 30990 26376
rect 31662 26324 31668 26376
rect 31720 26324 31726 26376
rect 27798 26256 27804 26308
rect 27856 26296 27862 26308
rect 28445 26299 28503 26305
rect 28445 26296 28457 26299
rect 27856 26268 28457 26296
rect 27856 26256 27862 26268
rect 28445 26265 28457 26268
rect 28491 26296 28503 26299
rect 28905 26299 28963 26305
rect 28905 26296 28917 26299
rect 28491 26268 28917 26296
rect 28491 26265 28503 26268
rect 28445 26259 28503 26265
rect 28828 26240 28856 26268
rect 28905 26265 28917 26268
rect 28951 26296 28963 26299
rect 29641 26299 29699 26305
rect 29641 26296 29653 26299
rect 28951 26268 29653 26296
rect 28951 26265 28963 26268
rect 28905 26259 28963 26265
rect 29641 26265 29653 26268
rect 29687 26265 29699 26299
rect 31910 26299 31968 26305
rect 31910 26296 31922 26299
rect 29641 26259 29699 26265
rect 30116 26268 31922 26296
rect 3513 26231 3571 26237
rect 3513 26197 3525 26231
rect 3559 26228 3571 26231
rect 3786 26228 3792 26240
rect 3559 26200 3792 26228
rect 3559 26197 3571 26200
rect 3513 26191 3571 26197
rect 3786 26188 3792 26200
rect 3844 26188 3850 26240
rect 16758 26188 16764 26240
rect 16816 26228 16822 26240
rect 17589 26231 17647 26237
rect 17589 26228 17601 26231
rect 16816 26200 17601 26228
rect 16816 26188 16822 26200
rect 17589 26197 17601 26200
rect 17635 26197 17647 26231
rect 17589 26191 17647 26197
rect 28810 26188 28816 26240
rect 28868 26188 28874 26240
rect 30116 26237 30144 26268
rect 31910 26265 31922 26268
rect 31956 26265 31968 26299
rect 31910 26259 31968 26265
rect 30101 26231 30159 26237
rect 30101 26197 30113 26231
rect 30147 26197 30159 26231
rect 30101 26191 30159 26197
rect 30834 26188 30840 26240
rect 30892 26188 30898 26240
rect 31573 26231 31631 26237
rect 31573 26197 31585 26231
rect 31619 26228 31631 26231
rect 32214 26228 32220 26240
rect 31619 26200 32220 26228
rect 31619 26197 31631 26200
rect 31573 26191 31631 26197
rect 32214 26188 32220 26200
rect 32272 26188 32278 26240
rect 33042 26188 33048 26240
rect 33100 26188 33106 26240
rect 1104 26138 34016 26160
rect 1104 26086 9138 26138
rect 9190 26086 9202 26138
rect 9254 26086 9266 26138
rect 9318 26086 9330 26138
rect 9382 26086 9394 26138
rect 9446 26086 17326 26138
rect 17378 26086 17390 26138
rect 17442 26086 17454 26138
rect 17506 26086 17518 26138
rect 17570 26086 17582 26138
rect 17634 26086 25514 26138
rect 25566 26086 25578 26138
rect 25630 26086 25642 26138
rect 25694 26086 25706 26138
rect 25758 26086 25770 26138
rect 25822 26086 33702 26138
rect 33754 26086 33766 26138
rect 33818 26086 33830 26138
rect 33882 26086 33894 26138
rect 33946 26086 33958 26138
rect 34010 26086 34016 26138
rect 1104 26064 34016 26086
rect 2866 25984 2872 26036
rect 2924 26024 2930 26036
rect 3237 26027 3295 26033
rect 3237 26024 3249 26027
rect 2924 25996 3249 26024
rect 2924 25984 2930 25996
rect 3237 25993 3249 25996
rect 3283 25993 3295 26027
rect 3237 25987 3295 25993
rect 3970 25984 3976 26036
rect 4028 25984 4034 26036
rect 17126 25984 17132 26036
rect 17184 26024 17190 26036
rect 17405 26027 17463 26033
rect 17405 26024 17417 26027
rect 17184 25996 17417 26024
rect 17184 25984 17190 25996
rect 17405 25993 17417 25996
rect 17451 25993 17463 26027
rect 17405 25987 17463 25993
rect 29825 26027 29883 26033
rect 29825 25993 29837 26027
rect 29871 26024 29883 26027
rect 30190 26024 30196 26036
rect 29871 25996 30196 26024
rect 29871 25993 29883 25996
rect 29825 25987 29883 25993
rect 30190 25984 30196 25996
rect 30248 25984 30254 26036
rect 33042 26024 33048 26036
rect 30484 25996 33048 26024
rect 30374 25956 30380 25968
rect 30346 25916 30380 25956
rect 30432 25916 30438 25968
rect 1762 25848 1768 25900
rect 1820 25848 1826 25900
rect 2032 25891 2090 25897
rect 2032 25857 2044 25891
rect 2078 25888 2090 25891
rect 2078 25860 4752 25888
rect 2078 25857 2090 25860
rect 2032 25851 2090 25857
rect 3786 25780 3792 25832
rect 3844 25780 3850 25832
rect 4724 25829 4752 25860
rect 4525 25823 4583 25829
rect 4525 25820 4537 25823
rect 3896 25792 4537 25820
rect 3145 25755 3203 25761
rect 3145 25721 3157 25755
rect 3191 25752 3203 25755
rect 3896 25752 3924 25792
rect 4525 25789 4537 25792
rect 4571 25789 4583 25823
rect 4525 25783 4583 25789
rect 4709 25823 4767 25829
rect 4709 25789 4721 25823
rect 4755 25789 4767 25823
rect 4709 25783 4767 25789
rect 4890 25780 4896 25832
rect 4948 25820 4954 25832
rect 5169 25823 5227 25829
rect 5169 25820 5181 25823
rect 4948 25792 5181 25820
rect 4948 25780 4954 25792
rect 5169 25789 5181 25792
rect 5215 25820 5227 25823
rect 5902 25820 5908 25832
rect 5215 25792 5908 25820
rect 5215 25789 5227 25792
rect 5169 25783 5227 25789
rect 5902 25780 5908 25792
rect 5960 25780 5966 25832
rect 16758 25780 16764 25832
rect 16816 25780 16822 25832
rect 28810 25780 28816 25832
rect 28868 25820 28874 25832
rect 29181 25823 29239 25829
rect 29181 25820 29193 25823
rect 28868 25792 29193 25820
rect 28868 25780 28874 25792
rect 29181 25789 29193 25792
rect 29227 25820 29239 25823
rect 29273 25823 29331 25829
rect 29273 25820 29285 25823
rect 29227 25792 29285 25820
rect 29227 25789 29239 25792
rect 29181 25783 29239 25789
rect 29273 25789 29285 25792
rect 29319 25820 29331 25823
rect 30346 25820 30374 25916
rect 30484 25897 30512 25996
rect 33042 25984 33048 25996
rect 33100 25984 33106 26036
rect 32306 25916 32312 25968
rect 32364 25956 32370 25968
rect 32585 25959 32643 25965
rect 32585 25956 32597 25959
rect 32364 25928 32597 25956
rect 32364 25916 32370 25928
rect 32585 25925 32597 25928
rect 32631 25925 32643 25959
rect 32585 25919 32643 25925
rect 30469 25891 30527 25897
rect 30469 25857 30481 25891
rect 30515 25857 30527 25891
rect 30469 25851 30527 25857
rect 32214 25848 32220 25900
rect 32272 25848 32278 25900
rect 29319 25792 30374 25820
rect 29319 25789 29331 25792
rect 29273 25783 29331 25789
rect 30558 25780 30564 25832
rect 30616 25780 30622 25832
rect 31202 25780 31208 25832
rect 31260 25780 31266 25832
rect 31294 25780 31300 25832
rect 31352 25780 31358 25832
rect 3191 25724 3924 25752
rect 3191 25721 3203 25724
rect 3145 25715 3203 25721
rect 4430 25712 4436 25764
rect 4488 25752 4494 25764
rect 4801 25755 4859 25761
rect 4801 25752 4813 25755
rect 4488 25724 4813 25752
rect 4488 25712 4494 25724
rect 4801 25721 4813 25724
rect 4847 25721 4859 25755
rect 4801 25715 4859 25721
rect 29641 25755 29699 25761
rect 29641 25721 29653 25755
rect 29687 25752 29699 25755
rect 30834 25752 30840 25764
rect 29687 25724 30840 25752
rect 29687 25721 29699 25724
rect 29641 25715 29699 25721
rect 30834 25712 30840 25724
rect 30892 25712 30898 25764
rect 29733 25687 29791 25693
rect 29733 25653 29745 25687
rect 29779 25684 29791 25687
rect 31754 25684 31760 25696
rect 29779 25656 31760 25684
rect 29779 25653 29791 25656
rect 29733 25647 29791 25653
rect 31754 25644 31760 25656
rect 31812 25644 31818 25696
rect 31938 25644 31944 25696
rect 31996 25644 32002 25696
rect 1104 25594 33856 25616
rect 1104 25542 5044 25594
rect 5096 25542 5108 25594
rect 5160 25542 5172 25594
rect 5224 25542 5236 25594
rect 5288 25542 5300 25594
rect 5352 25542 13232 25594
rect 13284 25542 13296 25594
rect 13348 25542 13360 25594
rect 13412 25542 13424 25594
rect 13476 25542 13488 25594
rect 13540 25542 21420 25594
rect 21472 25542 21484 25594
rect 21536 25542 21548 25594
rect 21600 25542 21612 25594
rect 21664 25542 21676 25594
rect 21728 25542 29608 25594
rect 29660 25542 29672 25594
rect 29724 25542 29736 25594
rect 29788 25542 29800 25594
rect 29852 25542 29864 25594
rect 29916 25542 33856 25594
rect 1104 25520 33856 25542
rect 1765 25483 1823 25489
rect 1765 25449 1777 25483
rect 1811 25480 1823 25483
rect 1811 25452 3188 25480
rect 1811 25449 1823 25452
rect 1765 25443 1823 25449
rect 3160 25412 3188 25452
rect 3418 25440 3424 25492
rect 3476 25480 3482 25492
rect 3789 25483 3847 25489
rect 3789 25480 3801 25483
rect 3476 25452 3801 25480
rect 3476 25440 3482 25452
rect 3789 25449 3801 25452
rect 3835 25449 3847 25483
rect 3789 25443 3847 25449
rect 4154 25440 4160 25492
rect 4212 25440 4218 25492
rect 29178 25440 29184 25492
rect 29236 25480 29242 25492
rect 29365 25483 29423 25489
rect 29365 25480 29377 25483
rect 29236 25452 29377 25480
rect 29236 25440 29242 25452
rect 29365 25449 29377 25452
rect 29411 25449 29423 25483
rect 29365 25443 29423 25449
rect 31202 25440 31208 25492
rect 31260 25480 31266 25492
rect 33045 25483 33103 25489
rect 33045 25480 33057 25483
rect 31260 25452 33057 25480
rect 31260 25440 31266 25452
rect 33045 25449 33057 25452
rect 33091 25449 33103 25483
rect 33045 25443 33103 25449
rect 4172 25412 4200 25440
rect 3160 25384 4200 25412
rect 7006 25344 7012 25356
rect 3620 25316 7012 25344
rect 3142 25236 3148 25288
rect 3200 25236 3206 25288
rect 3620 25285 3648 25316
rect 7006 25304 7012 25316
rect 7064 25304 7070 25356
rect 26970 25304 26976 25356
rect 27028 25344 27034 25356
rect 28534 25344 28540 25356
rect 27028 25316 28540 25344
rect 27028 25304 27034 25316
rect 28534 25304 28540 25316
rect 28592 25344 28598 25356
rect 30101 25347 30159 25353
rect 30101 25344 30113 25347
rect 28592 25316 30113 25344
rect 28592 25304 28598 25316
rect 30101 25313 30113 25316
rect 30147 25344 30159 25347
rect 31665 25347 31723 25353
rect 31665 25344 31677 25347
rect 30147 25316 31677 25344
rect 30147 25313 30159 25316
rect 30101 25307 30159 25313
rect 31665 25313 31677 25316
rect 31711 25313 31723 25347
rect 31665 25307 31723 25313
rect 3605 25279 3663 25285
rect 3605 25245 3617 25279
rect 3651 25245 3663 25279
rect 3605 25239 3663 25245
rect 4430 25236 4436 25288
rect 4488 25276 4494 25288
rect 5442 25276 5448 25288
rect 4488 25248 5448 25276
rect 4488 25236 4494 25248
rect 5442 25236 5448 25248
rect 5500 25236 5506 25288
rect 28718 25236 28724 25288
rect 28776 25236 28782 25288
rect 31570 25236 31576 25288
rect 31628 25236 31634 25288
rect 31754 25236 31760 25288
rect 31812 25276 31818 25288
rect 31921 25279 31979 25285
rect 31921 25276 31933 25279
rect 31812 25248 31933 25276
rect 31812 25236 31818 25248
rect 31921 25245 31933 25248
rect 31967 25245 31979 25279
rect 31921 25239 31979 25245
rect 2900 25211 2958 25217
rect 2900 25177 2912 25211
rect 2946 25208 2958 25211
rect 3237 25211 3295 25217
rect 3237 25208 3249 25211
rect 2946 25180 3249 25208
rect 2946 25177 2958 25180
rect 2900 25171 2958 25177
rect 3237 25177 3249 25180
rect 3283 25177 3295 25211
rect 3237 25171 3295 25177
rect 3421 25211 3479 25217
rect 3421 25177 3433 25211
rect 3467 25208 3479 25211
rect 4062 25208 4068 25220
rect 3467 25180 4068 25208
rect 3467 25177 3479 25180
rect 3421 25171 3479 25177
rect 4062 25168 4068 25180
rect 4120 25168 4126 25220
rect 30653 25211 30711 25217
rect 30653 25177 30665 25211
rect 30699 25208 30711 25211
rect 31110 25208 31116 25220
rect 30699 25180 31116 25208
rect 30699 25177 30711 25180
rect 30653 25171 30711 25177
rect 31110 25168 31116 25180
rect 31168 25168 31174 25220
rect 1104 25050 34016 25072
rect 1104 24998 9138 25050
rect 9190 24998 9202 25050
rect 9254 24998 9266 25050
rect 9318 24998 9330 25050
rect 9382 24998 9394 25050
rect 9446 24998 17326 25050
rect 17378 24998 17390 25050
rect 17442 24998 17454 25050
rect 17506 24998 17518 25050
rect 17570 24998 17582 25050
rect 17634 24998 25514 25050
rect 25566 24998 25578 25050
rect 25630 24998 25642 25050
rect 25694 24998 25706 25050
rect 25758 24998 25770 25050
rect 25822 24998 33702 25050
rect 33754 24998 33766 25050
rect 33818 24998 33830 25050
rect 33882 24998 33894 25050
rect 33946 24998 33958 25050
rect 34010 24998 34016 25050
rect 1104 24976 34016 24998
rect 31205 24939 31263 24945
rect 31205 24905 31217 24939
rect 31251 24936 31263 24939
rect 31294 24936 31300 24948
rect 31251 24908 31300 24936
rect 31251 24905 31263 24908
rect 31205 24899 31263 24905
rect 31294 24896 31300 24908
rect 31352 24896 31358 24948
rect 4062 24828 4068 24880
rect 4120 24868 4126 24880
rect 4890 24868 4896 24880
rect 4120 24840 4896 24868
rect 4120 24828 4126 24840
rect 4890 24828 4896 24840
rect 4948 24828 4954 24880
rect 31570 24828 31576 24880
rect 31628 24868 31634 24880
rect 32585 24871 32643 24877
rect 32585 24868 32597 24871
rect 31628 24840 32597 24868
rect 31628 24828 31634 24840
rect 32585 24837 32597 24840
rect 32631 24837 32643 24871
rect 32585 24831 32643 24837
rect 2590 24760 2596 24812
rect 2648 24760 2654 24812
rect 13193 24803 13251 24809
rect 13193 24769 13205 24803
rect 13239 24800 13251 24803
rect 15565 24803 15623 24809
rect 13239 24772 15148 24800
rect 13239 24769 13251 24772
rect 13193 24763 13251 24769
rect 934 24692 940 24744
rect 992 24732 998 24744
rect 1581 24735 1639 24741
rect 1581 24732 1593 24735
rect 992 24704 1593 24732
rect 992 24692 998 24704
rect 1581 24701 1593 24704
rect 1627 24701 1639 24735
rect 1581 24695 1639 24701
rect 2961 24735 3019 24741
rect 2961 24701 2973 24735
rect 3007 24732 3019 24735
rect 3326 24732 3332 24744
rect 3007 24704 3332 24732
rect 3007 24701 3019 24704
rect 2961 24695 3019 24701
rect 3326 24692 3332 24704
rect 3384 24692 3390 24744
rect 15120 24741 15148 24772
rect 15565 24769 15577 24803
rect 15611 24800 15623 24803
rect 15746 24800 15752 24812
rect 15611 24772 15752 24800
rect 15611 24769 15623 24772
rect 15565 24763 15623 24769
rect 15746 24760 15752 24772
rect 15804 24760 15810 24812
rect 15930 24760 15936 24812
rect 15988 24800 15994 24812
rect 16209 24803 16267 24809
rect 16209 24800 16221 24803
rect 15988 24772 16221 24800
rect 15988 24760 15994 24772
rect 16209 24769 16221 24772
rect 16255 24769 16267 24803
rect 16209 24763 16267 24769
rect 30558 24760 30564 24812
rect 30616 24760 30622 24812
rect 31938 24760 31944 24812
rect 31996 24800 32002 24812
rect 32217 24803 32275 24809
rect 32217 24800 32229 24803
rect 31996 24772 32229 24800
rect 31996 24760 32002 24772
rect 32217 24769 32229 24772
rect 32263 24769 32275 24803
rect 32217 24763 32275 24769
rect 13449 24735 13507 24741
rect 13449 24701 13461 24735
rect 13495 24701 13507 24735
rect 13449 24695 13507 24701
rect 15105 24735 15163 24741
rect 15105 24701 15117 24735
rect 15151 24701 15163 24735
rect 16758 24732 16764 24744
rect 15105 24695 15163 24701
rect 16546 24704 16764 24732
rect 3786 24624 3792 24676
rect 3844 24624 3850 24676
rect 3510 24556 3516 24608
rect 3568 24556 3574 24608
rect 3602 24556 3608 24608
rect 3660 24556 3666 24608
rect 12066 24556 12072 24608
rect 12124 24556 12130 24608
rect 13078 24556 13084 24608
rect 13136 24596 13142 24608
rect 13464 24596 13492 24695
rect 15289 24667 15347 24673
rect 15289 24633 15301 24667
rect 15335 24664 15347 24667
rect 16546 24664 16574 24704
rect 16758 24692 16764 24704
rect 16816 24692 16822 24744
rect 31846 24692 31852 24744
rect 31904 24692 31910 24744
rect 15335 24636 16574 24664
rect 15335 24633 15347 24636
rect 15289 24627 15347 24633
rect 13136 24568 13492 24596
rect 13136 24556 13142 24568
rect 15746 24556 15752 24608
rect 15804 24556 15810 24608
rect 30650 24556 30656 24608
rect 30708 24596 30714 24608
rect 31297 24599 31355 24605
rect 31297 24596 31309 24599
rect 30708 24568 31309 24596
rect 30708 24556 30714 24568
rect 31297 24565 31309 24568
rect 31343 24565 31355 24599
rect 31297 24559 31355 24565
rect 1104 24506 33856 24528
rect 1104 24454 5044 24506
rect 5096 24454 5108 24506
rect 5160 24454 5172 24506
rect 5224 24454 5236 24506
rect 5288 24454 5300 24506
rect 5352 24454 13232 24506
rect 13284 24454 13296 24506
rect 13348 24454 13360 24506
rect 13412 24454 13424 24506
rect 13476 24454 13488 24506
rect 13540 24454 21420 24506
rect 21472 24454 21484 24506
rect 21536 24454 21548 24506
rect 21600 24454 21612 24506
rect 21664 24454 21676 24506
rect 21728 24454 29608 24506
rect 29660 24454 29672 24506
rect 29724 24454 29736 24506
rect 29788 24454 29800 24506
rect 29852 24454 29864 24506
rect 29916 24454 33856 24506
rect 1104 24432 33856 24454
rect 2590 24392 2596 24404
rect 2424 24364 2596 24392
rect 2424 24265 2452 24364
rect 2590 24352 2596 24364
rect 2648 24352 2654 24404
rect 2958 24352 2964 24404
rect 3016 24352 3022 24404
rect 3326 24352 3332 24404
rect 3384 24392 3390 24404
rect 3789 24395 3847 24401
rect 3789 24392 3801 24395
rect 3384 24364 3801 24392
rect 3384 24352 3390 24364
rect 3789 24361 3801 24364
rect 3835 24361 3847 24395
rect 3789 24355 3847 24361
rect 15746 24352 15752 24404
rect 15804 24352 15810 24404
rect 30742 24352 30748 24404
rect 30800 24352 30806 24404
rect 2409 24259 2467 24265
rect 2409 24225 2421 24259
rect 2455 24225 2467 24259
rect 2409 24219 2467 24225
rect 3605 24259 3663 24265
rect 3605 24225 3617 24259
rect 3651 24256 3663 24259
rect 3694 24256 3700 24268
rect 3651 24228 3700 24256
rect 3651 24225 3663 24228
rect 3605 24219 3663 24225
rect 3694 24216 3700 24228
rect 3752 24256 3758 24268
rect 30760 24256 30788 24352
rect 31205 24327 31263 24333
rect 31205 24293 31217 24327
rect 31251 24324 31263 24327
rect 31294 24324 31300 24336
rect 31251 24296 31300 24324
rect 31251 24293 31263 24296
rect 31205 24287 31263 24293
rect 31294 24284 31300 24296
rect 31352 24284 31358 24336
rect 30837 24259 30895 24265
rect 30837 24256 30849 24259
rect 3752 24228 4752 24256
rect 30760 24228 30849 24256
rect 3752 24216 3758 24228
rect 4724 24200 4752 24228
rect 30837 24225 30849 24228
rect 30883 24225 30895 24259
rect 30837 24219 30895 24225
rect 2685 24191 2743 24197
rect 2685 24157 2697 24191
rect 2731 24188 2743 24191
rect 2958 24188 2964 24200
rect 2731 24160 2964 24188
rect 2731 24157 2743 24160
rect 2685 24151 2743 24157
rect 2958 24148 2964 24160
rect 3016 24148 3022 24200
rect 4338 24148 4344 24200
rect 4396 24148 4402 24200
rect 4706 24148 4712 24200
rect 4764 24148 4770 24200
rect 31386 24148 31392 24200
rect 31444 24148 31450 24200
rect 32306 24148 32312 24200
rect 32364 24148 32370 24200
rect 33318 24080 33324 24132
rect 33376 24080 33382 24132
rect 31294 24012 31300 24064
rect 31352 24012 31358 24064
rect 32030 24012 32036 24064
rect 32088 24012 32094 24064
rect 1104 23962 34016 23984
rect 1104 23910 9138 23962
rect 9190 23910 9202 23962
rect 9254 23910 9266 23962
rect 9318 23910 9330 23962
rect 9382 23910 9394 23962
rect 9446 23910 17326 23962
rect 17378 23910 17390 23962
rect 17442 23910 17454 23962
rect 17506 23910 17518 23962
rect 17570 23910 17582 23962
rect 17634 23910 25514 23962
rect 25566 23910 25578 23962
rect 25630 23910 25642 23962
rect 25694 23910 25706 23962
rect 25758 23910 25770 23962
rect 25822 23910 33702 23962
rect 33754 23910 33766 23962
rect 33818 23910 33830 23962
rect 33882 23910 33894 23962
rect 33946 23910 33958 23962
rect 34010 23910 34016 23962
rect 1104 23888 34016 23910
rect 3602 23808 3608 23860
rect 3660 23808 3666 23860
rect 4249 23851 4307 23857
rect 4249 23817 4261 23851
rect 4295 23848 4307 23851
rect 4338 23848 4344 23860
rect 4295 23820 4344 23848
rect 4295 23817 4307 23820
rect 4249 23811 4307 23817
rect 4338 23808 4344 23820
rect 4396 23808 4402 23860
rect 8297 23851 8355 23857
rect 8297 23848 8309 23851
rect 6886 23820 8309 23848
rect 3136 23783 3194 23789
rect 3136 23749 3148 23783
rect 3182 23780 3194 23783
rect 3620 23780 3648 23808
rect 3182 23752 3648 23780
rect 3182 23749 3194 23752
rect 3136 23743 3194 23749
rect 2590 23672 2596 23724
rect 2648 23672 2654 23724
rect 1578 23604 1584 23656
rect 1636 23604 1642 23656
rect 2869 23647 2927 23653
rect 2869 23613 2881 23647
rect 2915 23613 2927 23647
rect 2869 23607 2927 23613
rect 2884 23508 2912 23607
rect 6886 23576 6914 23820
rect 8297 23817 8309 23820
rect 8343 23848 8355 23851
rect 13078 23848 13084 23860
rect 8343 23820 13084 23848
rect 8343 23817 8355 23820
rect 8297 23811 8355 23817
rect 13078 23808 13084 23820
rect 13136 23808 13142 23860
rect 27614 23808 27620 23860
rect 27672 23808 27678 23860
rect 31205 23851 31263 23857
rect 31205 23817 31217 23851
rect 31251 23848 31263 23851
rect 31386 23848 31392 23860
rect 31251 23820 31392 23848
rect 31251 23817 31263 23820
rect 31205 23811 31263 23817
rect 31386 23808 31392 23820
rect 31444 23808 31450 23860
rect 31846 23808 31852 23860
rect 31904 23848 31910 23860
rect 33505 23851 33563 23857
rect 33505 23848 33517 23851
rect 31904 23820 33517 23848
rect 31904 23808 31910 23820
rect 33505 23817 33517 23820
rect 33551 23817 33563 23851
rect 33505 23811 33563 23817
rect 31294 23740 31300 23792
rect 31352 23780 31358 23792
rect 32370 23783 32428 23789
rect 32370 23780 32382 23783
rect 31352 23752 32382 23780
rect 31352 23740 31358 23752
rect 32370 23749 32382 23752
rect 32416 23749 32428 23783
rect 32370 23743 32428 23749
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23681 9643 23715
rect 28629 23715 28687 23721
rect 28629 23712 28641 23715
rect 9585 23675 9643 23681
rect 28460 23684 28641 23712
rect 4172 23548 6914 23576
rect 3142 23508 3148 23520
rect 2884 23480 3148 23508
rect 3142 23468 3148 23480
rect 3200 23508 3206 23520
rect 4172 23508 4200 23548
rect 9600 23520 9628 23675
rect 25406 23604 25412 23656
rect 25464 23644 25470 23656
rect 26973 23647 27031 23653
rect 26973 23644 26985 23647
rect 25464 23616 26985 23644
rect 25464 23604 25470 23616
rect 26973 23613 26985 23616
rect 27019 23613 27031 23647
rect 26973 23607 27031 23613
rect 28460 23585 28488 23684
rect 28629 23681 28641 23684
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 30377 23715 30435 23721
rect 30377 23681 30389 23715
rect 30423 23712 30435 23715
rect 31662 23712 31668 23724
rect 30423 23684 31668 23712
rect 30423 23681 30435 23684
rect 30377 23675 30435 23681
rect 31662 23672 31668 23684
rect 31720 23712 31726 23724
rect 32125 23715 32183 23721
rect 32125 23712 32137 23715
rect 31720 23684 32137 23712
rect 31720 23672 31726 23684
rect 32125 23681 32137 23684
rect 32171 23681 32183 23715
rect 32125 23675 32183 23681
rect 30650 23604 30656 23656
rect 30708 23604 30714 23656
rect 31941 23647 31999 23653
rect 31941 23613 31953 23647
rect 31987 23613 31999 23647
rect 31941 23607 31999 23613
rect 28445 23579 28503 23585
rect 28445 23576 28457 23579
rect 25884 23548 28457 23576
rect 25884 23520 25912 23548
rect 28445 23545 28457 23548
rect 28491 23545 28503 23579
rect 28445 23539 28503 23545
rect 3200 23480 4200 23508
rect 3200 23468 3206 23480
rect 9582 23468 9588 23520
rect 9640 23508 9646 23520
rect 9861 23511 9919 23517
rect 9861 23508 9873 23511
rect 9640 23480 9873 23508
rect 9640 23468 9646 23480
rect 9861 23477 9873 23480
rect 9907 23477 9919 23511
rect 9861 23471 9919 23477
rect 25866 23468 25872 23520
rect 25924 23468 25930 23520
rect 31294 23468 31300 23520
rect 31352 23468 31358 23520
rect 31956 23508 31984 23607
rect 33042 23508 33048 23520
rect 31956 23480 33048 23508
rect 33042 23468 33048 23480
rect 33100 23468 33106 23520
rect 1104 23418 33856 23440
rect 1104 23366 5044 23418
rect 5096 23366 5108 23418
rect 5160 23366 5172 23418
rect 5224 23366 5236 23418
rect 5288 23366 5300 23418
rect 5352 23366 13232 23418
rect 13284 23366 13296 23418
rect 13348 23366 13360 23418
rect 13412 23366 13424 23418
rect 13476 23366 13488 23418
rect 13540 23366 21420 23418
rect 21472 23366 21484 23418
rect 21536 23366 21548 23418
rect 21600 23366 21612 23418
rect 21664 23366 21676 23418
rect 21728 23366 29608 23418
rect 29660 23366 29672 23418
rect 29724 23366 29736 23418
rect 29788 23366 29800 23418
rect 29852 23366 29864 23418
rect 29916 23366 33856 23418
rect 1104 23344 33856 23366
rect 2958 23264 2964 23316
rect 3016 23264 3022 23316
rect 4430 23264 4436 23316
rect 4488 23264 4494 23316
rect 18138 23264 18144 23316
rect 18196 23264 18202 23316
rect 26970 23264 26976 23316
rect 27028 23304 27034 23316
rect 27341 23307 27399 23313
rect 27341 23304 27353 23307
rect 27028 23276 27353 23304
rect 27028 23264 27034 23276
rect 27341 23273 27353 23276
rect 27387 23273 27399 23307
rect 27341 23267 27399 23273
rect 30742 23264 30748 23316
rect 30800 23304 30806 23316
rect 30800 23276 30880 23304
rect 30800 23264 30806 23276
rect 4614 23196 4620 23248
rect 4672 23196 4678 23248
rect 2409 23171 2467 23177
rect 2409 23137 2421 23171
rect 2455 23168 2467 23171
rect 2590 23168 2596 23180
rect 2455 23140 2596 23168
rect 2455 23137 2467 23140
rect 2409 23131 2467 23137
rect 2590 23128 2596 23140
rect 2648 23128 2654 23180
rect 3510 23128 3516 23180
rect 3568 23128 3574 23180
rect 30852 23177 30880 23276
rect 31205 23239 31263 23245
rect 31205 23205 31217 23239
rect 31251 23236 31263 23239
rect 31386 23236 31392 23248
rect 31251 23208 31392 23236
rect 31251 23205 31263 23208
rect 31205 23199 31263 23205
rect 31386 23196 31392 23208
rect 31444 23196 31450 23248
rect 30837 23171 30895 23177
rect 30837 23137 30849 23171
rect 30883 23137 30895 23171
rect 30837 23131 30895 23137
rect 31294 23128 31300 23180
rect 31352 23168 31358 23180
rect 31941 23171 31999 23177
rect 31941 23168 31953 23171
rect 31352 23140 31953 23168
rect 31352 23128 31358 23140
rect 31941 23137 31953 23140
rect 31987 23137 31999 23171
rect 31941 23131 31999 23137
rect 32306 23128 32312 23180
rect 32364 23168 32370 23180
rect 32493 23171 32551 23177
rect 32493 23168 32505 23171
rect 32364 23140 32505 23168
rect 32364 23128 32370 23140
rect 32493 23137 32505 23140
rect 32539 23137 32551 23171
rect 32493 23131 32551 23137
rect 2685 23103 2743 23109
rect 2685 23069 2697 23103
rect 2731 23100 2743 23103
rect 3234 23100 3240 23112
rect 2731 23072 3240 23100
rect 2731 23069 2743 23072
rect 2685 23063 2743 23069
rect 3234 23060 3240 23072
rect 3292 23060 3298 23112
rect 3786 23060 3792 23112
rect 3844 23060 3850 23112
rect 17218 23060 17224 23112
rect 17276 23100 17282 23112
rect 17497 23103 17555 23109
rect 17497 23100 17509 23103
rect 17276 23072 17509 23100
rect 17276 23060 17282 23072
rect 17497 23069 17509 23072
rect 17543 23069 17555 23103
rect 17497 23063 17555 23069
rect 32214 23060 32220 23112
rect 32272 23060 32278 23112
rect 4890 22992 4896 23044
rect 4948 23032 4954 23044
rect 4985 23035 5043 23041
rect 4985 23032 4997 23035
rect 4948 23004 4997 23032
rect 4948 22992 4954 23004
rect 4985 23001 4997 23004
rect 5031 23001 5043 23035
rect 26053 23035 26111 23041
rect 26053 23032 26065 23035
rect 4985 22995 5043 23001
rect 25884 23004 26065 23032
rect 25884 22976 25912 23004
rect 26053 23001 26065 23004
rect 26099 23001 26111 23035
rect 26053 22995 26111 23001
rect 4522 22924 4528 22976
rect 4580 22924 4586 22976
rect 25866 22924 25872 22976
rect 25924 22924 25930 22976
rect 31294 22924 31300 22976
rect 31352 22924 31358 22976
rect 31386 22924 31392 22976
rect 31444 22924 31450 22976
rect 1104 22874 34016 22896
rect 1104 22822 9138 22874
rect 9190 22822 9202 22874
rect 9254 22822 9266 22874
rect 9318 22822 9330 22874
rect 9382 22822 9394 22874
rect 9446 22822 17326 22874
rect 17378 22822 17390 22874
rect 17442 22822 17454 22874
rect 17506 22822 17518 22874
rect 17570 22822 17582 22874
rect 17634 22822 25514 22874
rect 25566 22822 25578 22874
rect 25630 22822 25642 22874
rect 25694 22822 25706 22874
rect 25758 22822 25770 22874
rect 25822 22822 33702 22874
rect 33754 22822 33766 22874
rect 33818 22822 33830 22874
rect 33882 22822 33894 22874
rect 33946 22822 33958 22874
rect 34010 22822 34016 22874
rect 1104 22800 34016 22822
rect 3510 22720 3516 22772
rect 3568 22720 3574 22772
rect 28537 22763 28595 22769
rect 28537 22729 28549 22763
rect 28583 22760 28595 22763
rect 28718 22760 28724 22772
rect 28583 22732 28724 22760
rect 28583 22729 28595 22732
rect 28537 22723 28595 22729
rect 28718 22720 28724 22732
rect 28776 22720 28782 22772
rect 3528 22692 3556 22720
rect 3528 22664 4844 22692
rect 1762 22584 1768 22636
rect 1820 22584 1826 22636
rect 2032 22627 2090 22633
rect 2032 22593 2044 22627
rect 2078 22624 2090 22627
rect 2078 22596 4752 22624
rect 2078 22593 2090 22596
rect 2032 22587 2090 22593
rect 4724 22565 4752 22596
rect 3329 22559 3387 22565
rect 3329 22525 3341 22559
rect 3375 22556 3387 22559
rect 3973 22559 4031 22565
rect 3973 22556 3985 22559
rect 3375 22528 3985 22556
rect 3375 22525 3387 22528
rect 3329 22519 3387 22525
rect 3973 22525 3985 22528
rect 4019 22525 4031 22559
rect 3973 22519 4031 22525
rect 4525 22559 4583 22565
rect 4525 22525 4537 22559
rect 4571 22525 4583 22559
rect 4525 22519 4583 22525
rect 4709 22559 4767 22565
rect 4709 22525 4721 22559
rect 4755 22525 4767 22559
rect 4709 22519 4767 22525
rect 3145 22491 3203 22497
rect 3145 22457 3157 22491
rect 3191 22488 3203 22491
rect 4540 22488 4568 22519
rect 4816 22497 4844 22664
rect 31941 22627 31999 22633
rect 31941 22593 31953 22627
rect 31987 22593 31999 22627
rect 31941 22587 31999 22593
rect 4890 22516 4896 22568
rect 4948 22556 4954 22568
rect 5169 22559 5227 22565
rect 5169 22556 5181 22559
rect 4948 22528 5181 22556
rect 4948 22516 4954 22528
rect 5169 22525 5181 22528
rect 5215 22525 5227 22559
rect 5169 22519 5227 22525
rect 26786 22516 26792 22568
rect 26844 22556 26850 22568
rect 27893 22559 27951 22565
rect 27893 22556 27905 22559
rect 26844 22528 27905 22556
rect 26844 22516 26850 22528
rect 27893 22525 27905 22528
rect 27939 22525 27951 22559
rect 27893 22519 27951 22525
rect 31478 22516 31484 22568
rect 31536 22516 31542 22568
rect 31956 22556 31984 22587
rect 32030 22584 32036 22636
rect 32088 22624 32094 22636
rect 32217 22627 32275 22633
rect 32217 22624 32229 22627
rect 32088 22596 32229 22624
rect 32088 22584 32094 22596
rect 32217 22593 32229 22596
rect 32263 22593 32275 22627
rect 32217 22587 32275 22593
rect 32493 22559 32551 22565
rect 32493 22556 32505 22559
rect 31956 22528 32505 22556
rect 32493 22525 32505 22528
rect 32539 22525 32551 22559
rect 32493 22519 32551 22525
rect 3191 22460 4568 22488
rect 4801 22491 4859 22497
rect 3191 22457 3203 22460
rect 3145 22451 3203 22457
rect 4801 22457 4813 22491
rect 4847 22457 4859 22491
rect 4801 22451 4859 22457
rect 3881 22423 3939 22429
rect 3881 22389 3893 22423
rect 3927 22420 3939 22423
rect 4338 22420 4344 22432
rect 3927 22392 4344 22420
rect 3927 22389 3939 22392
rect 3881 22383 3939 22389
rect 4338 22380 4344 22392
rect 4396 22380 4402 22432
rect 1104 22330 33856 22352
rect 1104 22278 5044 22330
rect 5096 22278 5108 22330
rect 5160 22278 5172 22330
rect 5224 22278 5236 22330
rect 5288 22278 5300 22330
rect 5352 22278 13232 22330
rect 13284 22278 13296 22330
rect 13348 22278 13360 22330
rect 13412 22278 13424 22330
rect 13476 22278 13488 22330
rect 13540 22278 21420 22330
rect 21472 22278 21484 22330
rect 21536 22278 21548 22330
rect 21600 22278 21612 22330
rect 21664 22278 21676 22330
rect 21728 22278 29608 22330
rect 29660 22278 29672 22330
rect 29724 22278 29736 22330
rect 29788 22278 29800 22330
rect 29852 22278 29864 22330
rect 29916 22278 33856 22330
rect 1104 22256 33856 22278
rect 3234 22176 3240 22228
rect 3292 22216 3298 22228
rect 3789 22219 3847 22225
rect 3789 22216 3801 22219
rect 3292 22188 3801 22216
rect 3292 22176 3298 22188
rect 3789 22185 3801 22188
rect 3835 22185 3847 22219
rect 3789 22179 3847 22185
rect 31573 22219 31631 22225
rect 31573 22185 31585 22219
rect 31619 22216 31631 22219
rect 32030 22216 32036 22228
rect 31619 22188 32036 22216
rect 31619 22185 31631 22188
rect 31573 22179 31631 22185
rect 32030 22176 32036 22188
rect 32088 22176 32094 22228
rect 33042 22176 33048 22228
rect 33100 22176 33106 22228
rect 1762 22040 1768 22092
rect 1820 22040 1826 22092
rect 4338 22040 4344 22092
rect 4396 22040 4402 22092
rect 31021 22083 31079 22089
rect 31021 22049 31033 22083
rect 31067 22080 31079 22083
rect 31386 22080 31392 22092
rect 31067 22052 31392 22080
rect 31067 22049 31079 22052
rect 31021 22043 31079 22049
rect 31386 22040 31392 22052
rect 31444 22040 31450 22092
rect 2032 22015 2090 22021
rect 2032 21981 2044 22015
rect 2078 22012 2090 22015
rect 4522 22012 4528 22024
rect 2078 21984 4528 22012
rect 2078 21981 2090 21984
rect 2032 21975 2090 21981
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 31662 21972 31668 22024
rect 31720 21972 31726 22024
rect 31294 21904 31300 21956
rect 31352 21944 31358 21956
rect 31910 21947 31968 21953
rect 31910 21944 31922 21947
rect 31352 21916 31922 21944
rect 31352 21904 31358 21916
rect 31910 21913 31922 21916
rect 31956 21913 31968 21947
rect 31910 21907 31968 21913
rect 3145 21879 3203 21885
rect 3145 21845 3157 21879
rect 3191 21876 3203 21879
rect 4614 21876 4620 21888
rect 3191 21848 4620 21876
rect 3191 21845 3203 21848
rect 3145 21839 3203 21845
rect 4614 21836 4620 21848
rect 4672 21836 4678 21888
rect 1104 21786 34016 21808
rect 1104 21734 9138 21786
rect 9190 21734 9202 21786
rect 9254 21734 9266 21786
rect 9318 21734 9330 21786
rect 9382 21734 9394 21786
rect 9446 21734 17326 21786
rect 17378 21734 17390 21786
rect 17442 21734 17454 21786
rect 17506 21734 17518 21786
rect 17570 21734 17582 21786
rect 17634 21734 25514 21786
rect 25566 21734 25578 21786
rect 25630 21734 25642 21786
rect 25694 21734 25706 21786
rect 25758 21734 25770 21786
rect 25822 21734 33702 21786
rect 33754 21734 33766 21786
rect 33818 21734 33830 21786
rect 33882 21734 33894 21786
rect 33946 21734 33958 21786
rect 34010 21734 34016 21786
rect 1104 21712 34016 21734
rect 30653 21607 30711 21613
rect 30653 21573 30665 21607
rect 30699 21604 30711 21607
rect 30742 21604 30748 21616
rect 30699 21576 30748 21604
rect 30699 21573 30711 21576
rect 30653 21567 30711 21573
rect 30742 21564 30748 21576
rect 30800 21564 30806 21616
rect 2590 21496 2596 21548
rect 2648 21496 2654 21548
rect 32306 21496 32312 21548
rect 32364 21496 32370 21548
rect 934 21428 940 21480
rect 992 21468 998 21480
rect 1581 21471 1639 21477
rect 1581 21468 1593 21471
rect 992 21440 1593 21468
rect 992 21428 998 21440
rect 1581 21437 1593 21440
rect 1627 21437 1639 21471
rect 1581 21431 1639 21437
rect 2961 21471 3019 21477
rect 2961 21437 2973 21471
rect 3007 21468 3019 21471
rect 3605 21471 3663 21477
rect 3605 21468 3617 21471
rect 3007 21440 3617 21468
rect 3007 21437 3019 21440
rect 2961 21431 3019 21437
rect 3605 21437 3617 21440
rect 3651 21437 3663 21471
rect 3605 21431 3663 21437
rect 3694 21428 3700 21480
rect 3752 21468 3758 21480
rect 4157 21471 4215 21477
rect 4157 21468 4169 21471
rect 3752 21440 4169 21468
rect 3752 21428 3758 21440
rect 4157 21437 4169 21440
rect 4203 21437 4215 21471
rect 4157 21431 4215 21437
rect 4338 21428 4344 21480
rect 4396 21428 4402 21480
rect 4798 21428 4804 21480
rect 4856 21428 4862 21480
rect 31938 21428 31944 21480
rect 31996 21428 32002 21480
rect 33318 21428 33324 21480
rect 33376 21428 33382 21480
rect 4356 21400 4384 21428
rect 4433 21403 4491 21409
rect 4433 21400 4445 21403
rect 4356 21372 4445 21400
rect 4433 21369 4445 21372
rect 4479 21369 4491 21403
rect 4433 21363 4491 21369
rect 31113 21403 31171 21409
rect 31113 21369 31125 21403
rect 31159 21400 31171 21403
rect 31386 21400 31392 21412
rect 31159 21372 31392 21400
rect 31159 21369 31171 21372
rect 31113 21363 31171 21369
rect 31386 21360 31392 21372
rect 31444 21360 31450 21412
rect 3510 21292 3516 21344
rect 3568 21292 3574 21344
rect 3602 21292 3608 21344
rect 3660 21332 3666 21344
rect 4341 21335 4399 21341
rect 4341 21332 4353 21335
rect 3660 21304 4353 21332
rect 3660 21292 3666 21304
rect 4341 21301 4353 21304
rect 4387 21301 4399 21335
rect 4341 21295 4399 21301
rect 31202 21292 31208 21344
rect 31260 21292 31266 21344
rect 31294 21292 31300 21344
rect 31352 21292 31358 21344
rect 1104 21242 33856 21264
rect 1104 21190 5044 21242
rect 5096 21190 5108 21242
rect 5160 21190 5172 21242
rect 5224 21190 5236 21242
rect 5288 21190 5300 21242
rect 5352 21190 13232 21242
rect 13284 21190 13296 21242
rect 13348 21190 13360 21242
rect 13412 21190 13424 21242
rect 13476 21190 13488 21242
rect 13540 21190 21420 21242
rect 21472 21190 21484 21242
rect 21536 21190 21548 21242
rect 21600 21190 21612 21242
rect 21664 21190 21676 21242
rect 21728 21190 29608 21242
rect 29660 21190 29672 21242
rect 29724 21190 29736 21242
rect 29788 21190 29800 21242
rect 29852 21190 29864 21242
rect 29916 21190 33856 21242
rect 1104 21168 33856 21190
rect 3145 21131 3203 21137
rect 3145 21097 3157 21131
rect 3191 21128 3203 21131
rect 3694 21128 3700 21140
rect 3191 21100 3700 21128
rect 3191 21097 3203 21100
rect 3145 21091 3203 21097
rect 3694 21088 3700 21100
rect 3752 21088 3758 21140
rect 3786 21088 3792 21140
rect 3844 21088 3850 21140
rect 25406 21088 25412 21140
rect 25464 21088 25470 21140
rect 31938 21088 31944 21140
rect 31996 21128 32002 21140
rect 33045 21131 33103 21137
rect 33045 21128 33057 21131
rect 31996 21100 33057 21128
rect 31996 21088 32002 21100
rect 33045 21097 33057 21100
rect 33091 21097 33103 21131
rect 33045 21091 33103 21097
rect 1762 20952 1768 21004
rect 1820 20952 1826 21004
rect 5261 20995 5319 21001
rect 5261 20992 5273 20995
rect 2792 20964 5273 20992
rect 1780 20924 1808 20952
rect 2792 20924 2820 20964
rect 5261 20961 5273 20964
rect 5307 20961 5319 20995
rect 5261 20955 5319 20961
rect 31021 20995 31079 21001
rect 31021 20961 31033 20995
rect 31067 20992 31079 20995
rect 31294 20992 31300 21004
rect 31067 20964 31300 20992
rect 31067 20961 31079 20964
rect 31021 20955 31079 20961
rect 31294 20952 31300 20964
rect 31352 20952 31358 21004
rect 1780 20896 2820 20924
rect 3602 20884 3608 20936
rect 3660 20884 3666 20936
rect 4433 20927 4491 20933
rect 4433 20893 4445 20927
rect 4479 20924 4491 20927
rect 4522 20924 4528 20936
rect 4479 20896 4528 20924
rect 4479 20893 4491 20896
rect 4433 20887 4491 20893
rect 4522 20884 4528 20896
rect 4580 20884 4586 20936
rect 24762 20884 24768 20936
rect 24820 20884 24826 20936
rect 31202 20884 31208 20936
rect 31260 20884 31266 20936
rect 31662 20884 31668 20936
rect 31720 20884 31726 20936
rect 2032 20859 2090 20865
rect 2032 20825 2044 20859
rect 2078 20856 2090 20859
rect 3620 20856 3648 20884
rect 2078 20828 3648 20856
rect 7009 20859 7067 20865
rect 2078 20825 2090 20828
rect 2032 20819 2090 20825
rect 7009 20825 7021 20859
rect 7055 20825 7067 20859
rect 31220 20856 31248 20884
rect 31910 20859 31968 20865
rect 31910 20856 31922 20859
rect 31220 20828 31922 20856
rect 7009 20819 7067 20825
rect 31910 20825 31922 20828
rect 31956 20825 31968 20859
rect 31910 20819 31968 20825
rect 7024 20788 7052 20819
rect 7377 20791 7435 20797
rect 7377 20788 7389 20791
rect 7024 20760 7389 20788
rect 7377 20757 7389 20760
rect 7423 20788 7435 20791
rect 9582 20788 9588 20800
rect 7423 20760 9588 20788
rect 7423 20757 7435 20760
rect 7377 20751 7435 20757
rect 9582 20748 9588 20760
rect 9640 20788 9646 20800
rect 10318 20788 10324 20800
rect 9640 20760 10324 20788
rect 9640 20748 9646 20760
rect 10318 20748 10324 20760
rect 10376 20748 10382 20800
rect 31570 20748 31576 20800
rect 31628 20748 31634 20800
rect 1104 20698 34016 20720
rect 1104 20646 9138 20698
rect 9190 20646 9202 20698
rect 9254 20646 9266 20698
rect 9318 20646 9330 20698
rect 9382 20646 9394 20698
rect 9446 20646 17326 20698
rect 17378 20646 17390 20698
rect 17442 20646 17454 20698
rect 17506 20646 17518 20698
rect 17570 20646 17582 20698
rect 17634 20646 25514 20698
rect 25566 20646 25578 20698
rect 25630 20646 25642 20698
rect 25694 20646 25706 20698
rect 25758 20646 25770 20698
rect 25822 20646 33702 20698
rect 33754 20646 33766 20698
rect 33818 20646 33830 20698
rect 33882 20646 33894 20698
rect 33946 20646 33958 20698
rect 34010 20646 34016 20698
rect 1104 20624 34016 20646
rect 2317 20519 2375 20525
rect 2317 20485 2329 20519
rect 2363 20516 2375 20519
rect 2590 20516 2596 20528
rect 2363 20488 2596 20516
rect 2363 20485 2375 20488
rect 2317 20479 2375 20485
rect 2590 20476 2596 20488
rect 2648 20476 2654 20528
rect 32306 20476 32312 20528
rect 32364 20516 32370 20528
rect 32585 20519 32643 20525
rect 32585 20516 32597 20519
rect 32364 20488 32597 20516
rect 32364 20476 32370 20488
rect 32585 20485 32597 20488
rect 32631 20485 32643 20519
rect 32585 20479 32643 20485
rect 2685 20451 2743 20457
rect 2685 20417 2697 20451
rect 2731 20448 2743 20451
rect 2961 20451 3019 20457
rect 2961 20448 2973 20451
rect 2731 20420 2973 20448
rect 2731 20417 2743 20420
rect 2685 20411 2743 20417
rect 2961 20417 2973 20420
rect 3007 20417 3019 20451
rect 2961 20411 3019 20417
rect 31941 20451 31999 20457
rect 31941 20417 31953 20451
rect 31987 20448 31999 20451
rect 32217 20451 32275 20457
rect 32217 20448 32229 20451
rect 31987 20420 32229 20448
rect 31987 20417 31999 20420
rect 31941 20411 31999 20417
rect 32217 20417 32229 20420
rect 32263 20417 32275 20451
rect 32217 20411 32275 20417
rect 3602 20340 3608 20392
rect 3660 20340 3666 20392
rect 31389 20383 31447 20389
rect 31389 20349 31401 20383
rect 31435 20380 31447 20383
rect 31570 20380 31576 20392
rect 31435 20352 31576 20380
rect 31435 20349 31447 20352
rect 31389 20343 31447 20349
rect 31570 20340 31576 20352
rect 31628 20380 31634 20392
rect 31846 20380 31852 20392
rect 31628 20352 31852 20380
rect 31628 20340 31634 20352
rect 31846 20340 31852 20352
rect 31904 20340 31910 20392
rect 1104 20154 33856 20176
rect 1104 20102 5044 20154
rect 5096 20102 5108 20154
rect 5160 20102 5172 20154
rect 5224 20102 5236 20154
rect 5288 20102 5300 20154
rect 5352 20102 13232 20154
rect 13284 20102 13296 20154
rect 13348 20102 13360 20154
rect 13412 20102 13424 20154
rect 13476 20102 13488 20154
rect 13540 20102 21420 20154
rect 21472 20102 21484 20154
rect 21536 20102 21548 20154
rect 21600 20102 21612 20154
rect 21664 20102 21676 20154
rect 21728 20102 29608 20154
rect 29660 20102 29672 20154
rect 29724 20102 29736 20154
rect 29788 20102 29800 20154
rect 29852 20102 29864 20154
rect 29916 20102 33856 20154
rect 1104 20080 33856 20102
rect 17218 20000 17224 20052
rect 17276 20000 17282 20052
rect 30742 20000 30748 20052
rect 30800 20040 30806 20052
rect 31389 20043 31447 20049
rect 31389 20040 31401 20043
rect 30800 20012 31401 20040
rect 30800 20000 30806 20012
rect 31389 20009 31401 20012
rect 31435 20009 31447 20043
rect 31389 20003 31447 20009
rect 1762 19864 1768 19916
rect 1820 19864 1826 19916
rect 31404 19904 31432 20003
rect 31846 19932 31852 19984
rect 31904 19932 31910 19984
rect 31573 19907 31631 19913
rect 31573 19904 31585 19907
rect 31404 19876 31585 19904
rect 31573 19873 31585 19876
rect 31619 19873 31631 19907
rect 31573 19867 31631 19873
rect 4430 19796 4436 19848
rect 4488 19796 4494 19848
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19836 18659 19839
rect 18647 19808 19012 19836
rect 18647 19805 18659 19808
rect 18601 19799 18659 19805
rect 2032 19771 2090 19777
rect 2032 19737 2044 19771
rect 2078 19768 2090 19771
rect 3234 19768 3240 19780
rect 2078 19740 3240 19768
rect 2078 19737 2090 19740
rect 2032 19731 2090 19737
rect 3234 19728 3240 19740
rect 3292 19728 3298 19780
rect 18046 19728 18052 19780
rect 18104 19768 18110 19780
rect 18334 19771 18392 19777
rect 18334 19768 18346 19771
rect 18104 19740 18346 19768
rect 18104 19728 18110 19740
rect 18334 19737 18346 19740
rect 18380 19737 18392 19771
rect 18334 19731 18392 19737
rect 3142 19660 3148 19712
rect 3200 19660 3206 19712
rect 3786 19660 3792 19712
rect 3844 19660 3850 19712
rect 18984 19709 19012 19808
rect 28534 19796 28540 19848
rect 28592 19836 28598 19848
rect 32217 19839 32275 19845
rect 32217 19836 32229 19839
rect 28592 19808 32229 19836
rect 28592 19796 28598 19808
rect 32217 19805 32229 19808
rect 32263 19805 32275 19839
rect 32217 19799 32275 19805
rect 32582 19728 32588 19780
rect 32640 19728 32646 19780
rect 18969 19703 19027 19709
rect 18969 19669 18981 19703
rect 19015 19700 19027 19703
rect 25406 19700 25412 19712
rect 19015 19672 25412 19700
rect 19015 19669 19027 19672
rect 18969 19663 19027 19669
rect 25406 19660 25412 19672
rect 25464 19700 25470 19712
rect 26970 19700 26976 19712
rect 25464 19672 26976 19700
rect 25464 19660 25470 19672
rect 26970 19660 26976 19672
rect 27028 19660 27034 19712
rect 32030 19660 32036 19712
rect 32088 19660 32094 19712
rect 1104 19610 34016 19632
rect 1104 19558 9138 19610
rect 9190 19558 9202 19610
rect 9254 19558 9266 19610
rect 9318 19558 9330 19610
rect 9382 19558 9394 19610
rect 9446 19558 17326 19610
rect 17378 19558 17390 19610
rect 17442 19558 17454 19610
rect 17506 19558 17518 19610
rect 17570 19558 17582 19610
rect 17634 19558 25514 19610
rect 25566 19558 25578 19610
rect 25630 19558 25642 19610
rect 25694 19558 25706 19610
rect 25758 19558 25770 19610
rect 25822 19558 33702 19610
rect 33754 19558 33766 19610
rect 33818 19558 33830 19610
rect 33882 19558 33894 19610
rect 33946 19558 33958 19610
rect 34010 19558 34016 19610
rect 1104 19536 34016 19558
rect 3234 19456 3240 19508
rect 3292 19496 3298 19508
rect 4341 19499 4399 19505
rect 4341 19496 4353 19499
rect 3292 19468 4353 19496
rect 3292 19456 3298 19468
rect 4341 19465 4353 19468
rect 4387 19465 4399 19499
rect 4341 19459 4399 19465
rect 26786 19456 26792 19508
rect 26844 19456 26850 19508
rect 26970 19456 26976 19508
rect 27028 19496 27034 19508
rect 27157 19499 27215 19505
rect 27157 19496 27169 19499
rect 27028 19468 27169 19496
rect 27028 19456 27034 19468
rect 27157 19465 27169 19468
rect 27203 19465 27215 19499
rect 27157 19459 27215 19465
rect 25498 19388 25504 19440
rect 25556 19428 25562 19440
rect 25556 19400 25728 19428
rect 25556 19388 25562 19400
rect 934 19320 940 19372
rect 992 19360 998 19372
rect 1581 19363 1639 19369
rect 1581 19360 1593 19363
rect 992 19332 1593 19360
rect 992 19320 998 19332
rect 1581 19329 1593 19332
rect 1627 19329 1639 19363
rect 1581 19323 1639 19329
rect 2590 19320 2596 19372
rect 2648 19320 2654 19372
rect 3513 19363 3571 19369
rect 3513 19329 3525 19363
rect 3559 19360 3571 19363
rect 4430 19360 4436 19372
rect 3559 19332 4436 19360
rect 3559 19329 3571 19332
rect 3513 19323 3571 19329
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 25406 19320 25412 19372
rect 25464 19369 25470 19372
rect 25700 19369 25728 19400
rect 25464 19360 25474 19369
rect 25665 19363 25728 19369
rect 25464 19332 25509 19360
rect 25464 19323 25474 19332
rect 25665 19329 25677 19363
rect 25711 19332 25728 19363
rect 32309 19363 32367 19369
rect 25711 19329 25723 19332
rect 25665 19323 25723 19329
rect 32309 19329 32321 19363
rect 32355 19360 32367 19363
rect 32582 19360 32588 19372
rect 32355 19332 32588 19360
rect 32355 19329 32367 19332
rect 32309 19323 32367 19329
rect 25464 19320 25470 19323
rect 32582 19320 32588 19332
rect 32640 19320 32646 19372
rect 33318 19320 33324 19372
rect 33376 19320 33382 19372
rect 2866 19252 2872 19304
rect 2924 19252 2930 19304
rect 3694 19252 3700 19304
rect 3752 19252 3758 19304
rect 4798 19252 4804 19304
rect 4856 19252 4862 19304
rect 31294 19252 31300 19304
rect 31352 19252 31358 19304
rect 3602 19184 3608 19236
rect 3660 19224 3666 19236
rect 4433 19227 4491 19233
rect 4433 19224 4445 19227
rect 3660 19196 4445 19224
rect 3660 19184 3666 19196
rect 4433 19193 4445 19196
rect 4479 19193 4491 19227
rect 4433 19187 4491 19193
rect 4246 19116 4252 19168
rect 4304 19116 4310 19168
rect 31938 19116 31944 19168
rect 31996 19116 32002 19168
rect 1104 19066 33856 19088
rect 1104 19014 5044 19066
rect 5096 19014 5108 19066
rect 5160 19014 5172 19066
rect 5224 19014 5236 19066
rect 5288 19014 5300 19066
rect 5352 19014 13232 19066
rect 13284 19014 13296 19066
rect 13348 19014 13360 19066
rect 13412 19014 13424 19066
rect 13476 19014 13488 19066
rect 13540 19014 21420 19066
rect 21472 19014 21484 19066
rect 21536 19014 21548 19066
rect 21600 19014 21612 19066
rect 21664 19014 21676 19066
rect 21728 19014 29608 19066
rect 29660 19014 29672 19066
rect 29724 19014 29736 19066
rect 29788 19014 29800 19066
rect 29852 19014 29864 19066
rect 29916 19014 33856 19066
rect 1104 18992 33856 19014
rect 2866 18912 2872 18964
rect 2924 18912 2930 18964
rect 3694 18912 3700 18964
rect 3752 18952 3758 18964
rect 4525 18955 4583 18961
rect 4525 18952 4537 18955
rect 3752 18924 4537 18952
rect 3752 18912 3758 18924
rect 4525 18921 4537 18924
rect 4571 18921 4583 18955
rect 8938 18952 8944 18964
rect 4525 18915 4583 18921
rect 4632 18924 8944 18952
rect 1946 18844 1952 18896
rect 2004 18884 2010 18896
rect 4632 18884 4660 18924
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 18046 18912 18052 18964
rect 18104 18912 18110 18964
rect 2004 18856 4660 18884
rect 2004 18844 2010 18856
rect 4706 18844 4712 18896
rect 4764 18884 4770 18896
rect 5353 18887 5411 18893
rect 5353 18884 5365 18887
rect 4764 18856 5365 18884
rect 4764 18844 4770 18856
rect 5353 18853 5365 18856
rect 5399 18853 5411 18887
rect 5353 18847 5411 18853
rect 18233 18887 18291 18893
rect 18233 18853 18245 18887
rect 18279 18884 18291 18887
rect 19426 18884 19432 18896
rect 18279 18856 19432 18884
rect 18279 18853 18291 18856
rect 18233 18847 18291 18853
rect 19426 18844 19432 18856
rect 19484 18844 19490 18896
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18816 2467 18819
rect 2590 18816 2596 18828
rect 2455 18788 2596 18816
rect 2455 18785 2467 18788
rect 2409 18779 2467 18785
rect 2590 18776 2596 18788
rect 2648 18776 2654 18828
rect 3142 18776 3148 18828
rect 3200 18816 3206 18828
rect 3421 18819 3479 18825
rect 3421 18816 3433 18819
rect 3200 18788 3433 18816
rect 3200 18776 3206 18788
rect 3421 18785 3433 18788
rect 3467 18785 3479 18819
rect 3421 18779 3479 18785
rect 4246 18776 4252 18828
rect 4304 18816 4310 18828
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 4304 18788 4353 18816
rect 4304 18776 4310 18788
rect 4341 18785 4353 18788
rect 4387 18785 4399 18819
rect 4341 18779 4399 18785
rect 4798 18776 4804 18828
rect 4856 18816 4862 18828
rect 5721 18819 5779 18825
rect 5721 18816 5733 18819
rect 4856 18788 5733 18816
rect 4856 18776 4862 18788
rect 5721 18785 5733 18788
rect 5767 18785 5779 18819
rect 5721 18779 5779 18785
rect 31662 18776 31668 18828
rect 31720 18776 31726 18828
rect 2685 18751 2743 18757
rect 2685 18717 2697 18751
rect 2731 18748 2743 18751
rect 3786 18748 3792 18760
rect 2731 18720 3792 18748
rect 2731 18717 2743 18720
rect 2685 18711 2743 18717
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 4154 18708 4160 18760
rect 4212 18748 4218 18760
rect 5077 18751 5135 18757
rect 5077 18748 5089 18751
rect 4212 18720 5089 18748
rect 4212 18708 4218 18720
rect 5077 18717 5089 18720
rect 5123 18717 5135 18751
rect 5077 18711 5135 18717
rect 31021 18751 31079 18757
rect 31021 18717 31033 18751
rect 31067 18748 31079 18751
rect 31932 18751 31990 18757
rect 31067 18720 31754 18748
rect 31067 18717 31079 18720
rect 31021 18711 31079 18717
rect 18509 18683 18567 18689
rect 18509 18649 18521 18683
rect 18555 18680 18567 18683
rect 18877 18683 18935 18689
rect 18877 18680 18889 18683
rect 18555 18652 18889 18680
rect 18555 18649 18567 18652
rect 18509 18643 18567 18649
rect 18877 18649 18889 18652
rect 18923 18680 18935 18683
rect 30282 18680 30288 18692
rect 18923 18652 30288 18680
rect 18923 18649 18935 18652
rect 18877 18643 18935 18649
rect 30282 18640 30288 18652
rect 30340 18640 30346 18692
rect 3786 18572 3792 18624
rect 3844 18572 3850 18624
rect 3878 18572 3884 18624
rect 3936 18612 3942 18624
rect 5261 18615 5319 18621
rect 5261 18612 5273 18615
rect 3936 18584 5273 18612
rect 3936 18572 3942 18584
rect 5261 18581 5273 18584
rect 5307 18581 5319 18615
rect 5261 18575 5319 18581
rect 31570 18572 31576 18624
rect 31628 18572 31634 18624
rect 31726 18612 31754 18720
rect 31932 18717 31944 18751
rect 31978 18748 31990 18751
rect 31978 18720 32076 18748
rect 31978 18717 31990 18720
rect 31932 18711 31990 18717
rect 32048 18692 32076 18720
rect 32030 18640 32036 18692
rect 32088 18640 32094 18692
rect 33045 18615 33103 18621
rect 33045 18612 33057 18615
rect 31726 18584 33057 18612
rect 33045 18581 33057 18584
rect 33091 18581 33103 18615
rect 33045 18575 33103 18581
rect 1104 18522 34016 18544
rect 1104 18470 9138 18522
rect 9190 18470 9202 18522
rect 9254 18470 9266 18522
rect 9318 18470 9330 18522
rect 9382 18470 9394 18522
rect 9446 18470 17326 18522
rect 17378 18470 17390 18522
rect 17442 18470 17454 18522
rect 17506 18470 17518 18522
rect 17570 18470 17582 18522
rect 17634 18470 25514 18522
rect 25566 18470 25578 18522
rect 25630 18470 25642 18522
rect 25694 18470 25706 18522
rect 25758 18470 25770 18522
rect 25822 18470 33702 18522
rect 33754 18470 33766 18522
rect 33818 18470 33830 18522
rect 33882 18470 33894 18522
rect 33946 18470 33958 18522
rect 34010 18470 34016 18522
rect 1104 18448 34016 18470
rect 1946 18368 1952 18420
rect 2004 18368 2010 18420
rect 3786 18368 3792 18420
rect 3844 18368 3850 18420
rect 30374 18368 30380 18420
rect 30432 18408 30438 18420
rect 30653 18411 30711 18417
rect 30653 18408 30665 18411
rect 30432 18380 30665 18408
rect 30432 18368 30438 18380
rect 30653 18377 30665 18380
rect 30699 18377 30711 18411
rect 30653 18371 30711 18377
rect 30742 18368 30748 18420
rect 30800 18408 30806 18420
rect 31018 18408 31024 18420
rect 30800 18380 31024 18408
rect 30800 18368 30806 18380
rect 31018 18368 31024 18380
rect 31076 18368 31082 18420
rect 31294 18368 31300 18420
rect 31352 18368 31358 18420
rect 1765 18343 1823 18349
rect 1765 18309 1777 18343
rect 1811 18340 1823 18343
rect 1964 18340 1992 18368
rect 3804 18340 3832 18368
rect 1811 18312 1992 18340
rect 2700 18312 3832 18340
rect 1811 18309 1823 18312
rect 1765 18303 1823 18309
rect 2700 18281 2728 18312
rect 2685 18275 2743 18281
rect 2685 18241 2697 18275
rect 2731 18241 2743 18275
rect 2685 18235 2743 18241
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18241 2927 18275
rect 2869 18235 2927 18241
rect 2409 18207 2467 18213
rect 2409 18173 2421 18207
rect 2455 18204 2467 18207
rect 2884 18204 2912 18235
rect 31570 18232 31576 18284
rect 31628 18272 31634 18284
rect 31849 18275 31907 18281
rect 31849 18272 31861 18275
rect 31628 18244 31861 18272
rect 31628 18232 31634 18244
rect 31849 18241 31861 18244
rect 31895 18241 31907 18275
rect 31849 18235 31907 18241
rect 31938 18232 31944 18284
rect 31996 18272 32002 18284
rect 32217 18275 32275 18281
rect 32217 18272 32229 18275
rect 31996 18244 32229 18272
rect 31996 18232 32002 18244
rect 32217 18241 32229 18244
rect 32263 18241 32275 18275
rect 32217 18235 32275 18241
rect 2455 18176 2912 18204
rect 3329 18207 3387 18213
rect 2455 18173 2467 18176
rect 2409 18167 2467 18173
rect 3329 18173 3341 18207
rect 3375 18173 3387 18207
rect 4798 18204 4804 18216
rect 3329 18167 3387 18173
rect 4172 18176 4804 18204
rect 1302 18096 1308 18148
rect 1360 18136 1366 18148
rect 3344 18136 3372 18167
rect 1360 18108 3372 18136
rect 1360 18096 1366 18108
rect 1673 18071 1731 18077
rect 1673 18037 1685 18071
rect 1719 18068 1731 18071
rect 4172 18068 4200 18176
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 32490 18164 32496 18216
rect 32548 18164 32554 18216
rect 4430 18096 4436 18148
rect 4488 18096 4494 18148
rect 1719 18040 4200 18068
rect 1719 18037 1731 18040
rect 1673 18031 1731 18037
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 4341 18071 4399 18077
rect 4341 18068 4353 18071
rect 4304 18040 4353 18068
rect 4304 18028 4310 18040
rect 4341 18037 4353 18040
rect 4387 18037 4399 18071
rect 4341 18031 4399 18037
rect 1104 17978 33856 18000
rect 1104 17926 5044 17978
rect 5096 17926 5108 17978
rect 5160 17926 5172 17978
rect 5224 17926 5236 17978
rect 5288 17926 5300 17978
rect 5352 17926 13232 17978
rect 13284 17926 13296 17978
rect 13348 17926 13360 17978
rect 13412 17926 13424 17978
rect 13476 17926 13488 17978
rect 13540 17926 21420 17978
rect 21472 17926 21484 17978
rect 21536 17926 21548 17978
rect 21600 17926 21612 17978
rect 21664 17926 21676 17978
rect 21728 17926 29608 17978
rect 29660 17926 29672 17978
rect 29724 17926 29736 17978
rect 29788 17926 29800 17978
rect 29852 17926 29864 17978
rect 29916 17926 33856 17978
rect 1104 17904 33856 17926
rect 3145 17867 3203 17873
rect 3145 17833 3157 17867
rect 3191 17864 3203 17867
rect 4154 17864 4160 17876
rect 3191 17836 4160 17864
rect 3191 17833 3203 17836
rect 3145 17827 3203 17833
rect 4154 17824 4160 17836
rect 4212 17824 4218 17876
rect 21818 17824 21824 17876
rect 21876 17864 21882 17876
rect 22833 17867 22891 17873
rect 21876 17836 22416 17864
rect 21876 17824 21882 17836
rect 4338 17756 4344 17808
rect 4396 17796 4402 17808
rect 4617 17799 4675 17805
rect 4617 17796 4629 17799
rect 4396 17768 4629 17796
rect 4396 17756 4402 17768
rect 4617 17765 4629 17768
rect 4663 17765 4675 17799
rect 22388 17796 22416 17836
rect 22833 17833 22845 17867
rect 22879 17864 22891 17867
rect 24762 17864 24768 17876
rect 22879 17836 24768 17864
rect 22879 17833 22891 17836
rect 22833 17827 22891 17833
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 24397 17799 24455 17805
rect 24397 17796 24409 17799
rect 22388 17768 24409 17796
rect 4617 17759 4675 17765
rect 24397 17765 24409 17768
rect 24443 17765 24455 17799
rect 24397 17759 24455 17765
rect 30653 17799 30711 17805
rect 30653 17765 30665 17799
rect 30699 17796 30711 17799
rect 31294 17796 31300 17808
rect 30699 17768 31300 17796
rect 30699 17765 30711 17768
rect 30653 17759 30711 17765
rect 31294 17756 31300 17768
rect 31352 17756 31358 17808
rect 1762 17688 1768 17740
rect 1820 17688 1826 17740
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 4985 17731 5043 17737
rect 4985 17728 4997 17731
rect 4856 17700 4997 17728
rect 4856 17688 4862 17700
rect 4985 17697 4997 17700
rect 5031 17697 5043 17731
rect 4985 17691 5043 17697
rect 30282 17688 30288 17740
rect 30340 17728 30346 17740
rect 31018 17728 31024 17740
rect 30340 17700 31024 17728
rect 30340 17688 30346 17700
rect 31018 17688 31024 17700
rect 31076 17688 31082 17740
rect 33318 17688 33324 17740
rect 33376 17688 33382 17740
rect 4246 17620 4252 17672
rect 4304 17620 4310 17672
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17660 4491 17663
rect 4614 17660 4620 17672
rect 4479 17632 4620 17660
rect 4479 17629 4491 17632
rect 4433 17623 4491 17629
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 10376 17632 17325 17660
rect 10376 17620 10382 17632
rect 17313 17629 17325 17632
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 21453 17663 21511 17669
rect 21453 17629 21465 17663
rect 21499 17660 21511 17663
rect 22002 17660 22008 17672
rect 21499 17632 22008 17660
rect 21499 17629 21511 17632
rect 21453 17623 21511 17629
rect 2032 17595 2090 17601
rect 2032 17561 2044 17595
rect 2078 17592 2090 17595
rect 4264 17592 4292 17620
rect 2078 17564 4292 17592
rect 2078 17561 2090 17564
rect 2032 17555 2090 17561
rect 3510 17484 3516 17536
rect 3568 17524 3574 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 3568 17496 3801 17524
rect 3568 17484 3574 17496
rect 3789 17493 3801 17496
rect 3835 17493 3847 17527
rect 3789 17487 3847 17493
rect 4246 17484 4252 17536
rect 4304 17524 4310 17536
rect 4525 17527 4583 17533
rect 4525 17524 4537 17527
rect 4304 17496 4537 17524
rect 4304 17484 4310 17496
rect 4525 17493 4537 17496
rect 4571 17493 4583 17527
rect 17328 17524 17356 17623
rect 22002 17620 22008 17632
rect 22060 17660 22066 17672
rect 23109 17663 23167 17669
rect 23109 17660 23121 17663
rect 22060 17632 23121 17660
rect 22060 17620 22066 17632
rect 23109 17629 23121 17632
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 24946 17620 24952 17672
rect 25004 17620 25010 17672
rect 30374 17620 30380 17672
rect 30432 17660 30438 17672
rect 30837 17663 30895 17669
rect 30837 17660 30849 17663
rect 30432 17632 30849 17660
rect 30432 17620 30438 17632
rect 30837 17629 30849 17632
rect 30883 17629 30895 17663
rect 30837 17623 30895 17629
rect 32030 17620 32036 17672
rect 32088 17620 32094 17672
rect 32309 17663 32367 17669
rect 32309 17629 32321 17663
rect 32355 17660 32367 17663
rect 32490 17660 32496 17672
rect 32355 17632 32496 17660
rect 32355 17629 32367 17632
rect 32309 17623 32367 17629
rect 32490 17620 32496 17632
rect 32548 17620 32554 17672
rect 19058 17552 19064 17604
rect 19116 17552 19122 17604
rect 19150 17552 19156 17604
rect 19208 17592 19214 17604
rect 21698 17595 21756 17601
rect 21698 17592 21710 17595
rect 19208 17564 21710 17592
rect 19208 17552 19214 17564
rect 21698 17561 21710 17564
rect 21744 17561 21756 17595
rect 25866 17592 25872 17604
rect 21698 17555 21756 17561
rect 22756 17564 25872 17592
rect 22756 17524 22784 17564
rect 25866 17552 25872 17564
rect 25924 17552 25930 17604
rect 17328 17496 22784 17524
rect 4525 17487 4583 17493
rect 30742 17484 30748 17536
rect 30800 17484 30806 17536
rect 31386 17484 31392 17536
rect 31444 17484 31450 17536
rect 1104 17434 34016 17456
rect 1104 17382 9138 17434
rect 9190 17382 9202 17434
rect 9254 17382 9266 17434
rect 9318 17382 9330 17434
rect 9382 17382 9394 17434
rect 9446 17382 17326 17434
rect 17378 17382 17390 17434
rect 17442 17382 17454 17434
rect 17506 17382 17518 17434
rect 17570 17382 17582 17434
rect 17634 17382 25514 17434
rect 25566 17382 25578 17434
rect 25630 17382 25642 17434
rect 25694 17382 25706 17434
rect 25758 17382 25770 17434
rect 25822 17382 33702 17434
rect 33754 17382 33766 17434
rect 33818 17382 33830 17434
rect 33882 17382 33894 17434
rect 33946 17382 33958 17434
rect 34010 17382 34016 17434
rect 1104 17360 34016 17382
rect 3145 17323 3203 17329
rect 3145 17289 3157 17323
rect 3191 17320 3203 17323
rect 4522 17320 4528 17332
rect 3191 17292 4528 17320
rect 3191 17289 3203 17292
rect 3145 17283 3203 17289
rect 4522 17280 4528 17292
rect 4580 17280 4586 17332
rect 32030 17280 32036 17332
rect 32088 17320 32094 17332
rect 33505 17323 33563 17329
rect 33505 17320 33517 17323
rect 32088 17292 33517 17320
rect 32088 17280 32094 17292
rect 33505 17289 33517 17292
rect 33551 17289 33563 17323
rect 33505 17283 33563 17289
rect 30742 17212 30748 17264
rect 30800 17252 30806 17264
rect 32370 17255 32428 17261
rect 32370 17252 32382 17255
rect 30800 17224 32382 17252
rect 30800 17212 30806 17224
rect 32370 17221 32382 17224
rect 32416 17221 32428 17255
rect 32370 17215 32428 17221
rect 1762 17144 1768 17196
rect 1820 17144 1826 17196
rect 2032 17187 2090 17193
rect 2032 17153 2044 17187
rect 2078 17184 2090 17187
rect 4154 17184 4160 17196
rect 2078 17156 4160 17184
rect 2078 17153 2090 17156
rect 2032 17147 2090 17153
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 31938 17144 31944 17196
rect 31996 17144 32002 17196
rect 3326 17076 3332 17128
rect 3384 17076 3390 17128
rect 4522 17076 4528 17128
rect 4580 17076 4586 17128
rect 31478 17076 31484 17128
rect 31536 17076 31542 17128
rect 31662 17076 31668 17128
rect 31720 17116 31726 17128
rect 32125 17119 32183 17125
rect 32125 17116 32137 17119
rect 31720 17088 32137 17116
rect 31720 17076 31726 17088
rect 32125 17085 32137 17088
rect 32171 17085 32183 17119
rect 32125 17079 32183 17085
rect 3881 17051 3939 17057
rect 3881 17017 3893 17051
rect 3927 17048 3939 17051
rect 7466 17048 7472 17060
rect 3927 17020 7472 17048
rect 3927 17017 3939 17020
rect 3881 17011 3939 17017
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 3970 16940 3976 16992
rect 4028 16940 4034 16992
rect 1104 16890 33856 16912
rect 1104 16838 5044 16890
rect 5096 16838 5108 16890
rect 5160 16838 5172 16890
rect 5224 16838 5236 16890
rect 5288 16838 5300 16890
rect 5352 16838 13232 16890
rect 13284 16838 13296 16890
rect 13348 16838 13360 16890
rect 13412 16838 13424 16890
rect 13476 16838 13488 16890
rect 13540 16838 21420 16890
rect 21472 16838 21484 16890
rect 21536 16838 21548 16890
rect 21600 16838 21612 16890
rect 21664 16838 21676 16890
rect 21728 16838 29608 16890
rect 29660 16838 29672 16890
rect 29724 16838 29736 16890
rect 29788 16838 29800 16890
rect 29852 16838 29864 16890
rect 29916 16838 33856 16890
rect 1104 16816 33856 16838
rect 3326 16736 3332 16788
rect 3384 16776 3390 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3384 16748 3801 16776
rect 3384 16736 3390 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 4154 16736 4160 16788
rect 4212 16776 4218 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4212 16748 4537 16776
rect 4212 16736 4218 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 21818 16736 21824 16788
rect 21876 16736 21882 16788
rect 31938 16736 31944 16788
rect 31996 16776 32002 16788
rect 31996 16748 32536 16776
rect 31996 16736 32002 16748
rect 4614 16668 4620 16720
rect 4672 16668 4678 16720
rect 1762 16600 1768 16652
rect 1820 16600 1826 16652
rect 19518 16600 19524 16652
rect 19576 16600 19582 16652
rect 2032 16575 2090 16581
rect 2032 16541 2044 16575
rect 2078 16572 2090 16575
rect 3878 16572 3884 16584
rect 2078 16544 3884 16572
rect 2078 16541 2090 16544
rect 2032 16535 2090 16541
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4338 16532 4344 16584
rect 4396 16532 4402 16584
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 21453 16575 21511 16581
rect 21453 16572 21465 16575
rect 20772 16544 21465 16572
rect 20772 16532 20778 16544
rect 21453 16541 21465 16544
rect 21499 16572 21511 16575
rect 21836 16572 21864 16736
rect 31386 16600 31392 16652
rect 31444 16640 31450 16652
rect 32508 16649 32536 16748
rect 31941 16643 31999 16649
rect 31941 16640 31953 16643
rect 31444 16612 31953 16640
rect 31444 16600 31450 16612
rect 31941 16609 31953 16612
rect 31987 16609 31999 16643
rect 31941 16603 31999 16609
rect 32493 16643 32551 16649
rect 32493 16609 32505 16643
rect 32539 16609 32551 16643
rect 32493 16603 32551 16609
rect 21499 16544 21864 16572
rect 21499 16541 21511 16544
rect 21453 16535 21511 16541
rect 32214 16532 32220 16584
rect 32272 16532 32278 16584
rect 4985 16507 5043 16513
rect 4985 16473 4997 16507
rect 5031 16504 5043 16507
rect 20165 16507 20223 16513
rect 5031 16476 5065 16504
rect 5031 16473 5043 16476
rect 4985 16467 5043 16473
rect 20165 16473 20177 16507
rect 20211 16504 20223 16507
rect 24946 16504 24952 16516
rect 20211 16476 24952 16504
rect 20211 16473 20223 16476
rect 20165 16467 20223 16473
rect 3145 16439 3203 16445
rect 3145 16405 3157 16439
rect 3191 16436 3203 16439
rect 4522 16436 4528 16448
rect 3191 16408 4528 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 4798 16396 4804 16448
rect 4856 16436 4862 16448
rect 5000 16436 5028 16467
rect 24946 16464 24952 16476
rect 25004 16464 25010 16516
rect 5261 16439 5319 16445
rect 5261 16436 5273 16439
rect 4856 16408 5273 16436
rect 4856 16396 4862 16408
rect 5261 16405 5273 16408
rect 5307 16405 5319 16439
rect 5261 16399 5319 16405
rect 21637 16439 21695 16445
rect 21637 16405 21649 16439
rect 21683 16436 21695 16439
rect 28534 16436 28540 16448
rect 21683 16408 28540 16436
rect 21683 16405 21695 16408
rect 21637 16399 21695 16405
rect 28534 16396 28540 16408
rect 28592 16396 28598 16448
rect 31386 16396 31392 16448
rect 31444 16396 31450 16448
rect 1104 16346 34016 16368
rect 1104 16294 9138 16346
rect 9190 16294 9202 16346
rect 9254 16294 9266 16346
rect 9318 16294 9330 16346
rect 9382 16294 9394 16346
rect 9446 16294 17326 16346
rect 17378 16294 17390 16346
rect 17442 16294 17454 16346
rect 17506 16294 17518 16346
rect 17570 16294 17582 16346
rect 17634 16294 25514 16346
rect 25566 16294 25578 16346
rect 25630 16294 25642 16346
rect 25694 16294 25706 16346
rect 25758 16294 25770 16346
rect 25822 16294 33702 16346
rect 33754 16294 33766 16346
rect 33818 16294 33830 16346
rect 33882 16294 33894 16346
rect 33946 16294 33958 16346
rect 34010 16294 34016 16346
rect 1104 16272 34016 16294
rect 3513 16235 3571 16241
rect 3513 16201 3525 16235
rect 3559 16232 3571 16235
rect 4338 16232 4344 16244
rect 3559 16204 4344 16232
rect 3559 16201 3571 16204
rect 3513 16195 3571 16201
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 30374 16192 30380 16244
rect 30432 16232 30438 16244
rect 30561 16235 30619 16241
rect 30561 16232 30573 16235
rect 30432 16204 30573 16232
rect 30432 16192 30438 16204
rect 30561 16201 30573 16204
rect 30607 16201 30619 16235
rect 30561 16195 30619 16201
rect 31941 16235 31999 16241
rect 31941 16201 31953 16235
rect 31987 16232 31999 16235
rect 32214 16232 32220 16244
rect 31987 16204 32220 16232
rect 31987 16201 31999 16204
rect 31941 16195 31999 16201
rect 2400 16167 2458 16173
rect 2400 16133 2412 16167
rect 2446 16164 2458 16167
rect 4246 16164 4252 16176
rect 2446 16136 4252 16164
rect 2446 16133 2458 16136
rect 2400 16127 2458 16133
rect 4246 16124 4252 16136
rect 4304 16124 4310 16176
rect 30576 16164 30604 16195
rect 32214 16192 32220 16204
rect 32272 16192 32278 16244
rect 30745 16167 30803 16173
rect 30745 16164 30757 16167
rect 30576 16136 30757 16164
rect 30745 16133 30757 16136
rect 30791 16133 30803 16167
rect 30745 16127 30803 16133
rect 1489 16099 1547 16105
rect 1489 16065 1501 16099
rect 1535 16096 1547 16099
rect 3970 16096 3976 16108
rect 1535 16068 3976 16096
rect 1535 16065 1547 16068
rect 1489 16059 1547 16065
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4890 16056 4896 16108
rect 4948 16056 4954 16108
rect 31386 16056 31392 16108
rect 31444 16056 31450 16108
rect 32306 16056 32312 16108
rect 32364 16056 32370 16108
rect 1762 15988 1768 16040
rect 1820 16028 1826 16040
rect 2133 16031 2191 16037
rect 2133 16028 2145 16031
rect 1820 16000 2145 16028
rect 1820 15988 1826 16000
rect 2133 15997 2145 16000
rect 2179 15997 2191 16031
rect 2133 15991 2191 15997
rect 4338 15988 4344 16040
rect 4396 15988 4402 16040
rect 31113 15963 31171 15969
rect 31113 15929 31125 15963
rect 31159 15960 31171 15963
rect 31404 15960 31432 16056
rect 33318 15988 33324 16040
rect 33376 15988 33382 16040
rect 31159 15932 31432 15960
rect 31159 15929 31171 15932
rect 31113 15923 31171 15929
rect 2041 15895 2099 15901
rect 2041 15861 2053 15895
rect 2087 15892 2099 15895
rect 3418 15892 3424 15904
rect 2087 15864 3424 15892
rect 2087 15861 2099 15864
rect 2041 15855 2099 15861
rect 3418 15852 3424 15864
rect 3476 15852 3482 15904
rect 31205 15895 31263 15901
rect 31205 15861 31217 15895
rect 31251 15892 31263 15895
rect 31754 15892 31760 15904
rect 31251 15864 31760 15892
rect 31251 15861 31263 15864
rect 31205 15855 31263 15861
rect 31754 15852 31760 15864
rect 31812 15852 31818 15904
rect 1104 15802 33856 15824
rect 1104 15750 5044 15802
rect 5096 15750 5108 15802
rect 5160 15750 5172 15802
rect 5224 15750 5236 15802
rect 5288 15750 5300 15802
rect 5352 15750 13232 15802
rect 13284 15750 13296 15802
rect 13348 15750 13360 15802
rect 13412 15750 13424 15802
rect 13476 15750 13488 15802
rect 13540 15750 21420 15802
rect 21472 15750 21484 15802
rect 21536 15750 21548 15802
rect 21600 15750 21612 15802
rect 21664 15750 21676 15802
rect 21728 15750 29608 15802
rect 29660 15750 29672 15802
rect 29724 15750 29736 15802
rect 29788 15750 29800 15802
rect 29852 15750 29864 15802
rect 29916 15750 33856 15802
rect 1104 15728 33856 15750
rect 4338 15648 4344 15700
rect 4396 15648 4402 15700
rect 4890 15648 4896 15700
rect 4948 15688 4954 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 4948 15660 6929 15688
rect 4948 15648 4954 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 25041 15691 25099 15697
rect 25041 15657 25053 15691
rect 25087 15688 25099 15691
rect 25406 15688 25412 15700
rect 25087 15660 25412 15688
rect 25087 15657 25099 15660
rect 25041 15651 25099 15657
rect 25406 15648 25412 15660
rect 25464 15648 25470 15700
rect 1578 15512 1584 15564
rect 1636 15512 1642 15564
rect 4356 15552 4384 15648
rect 24946 15580 24952 15632
rect 25004 15580 25010 15632
rect 2700 15524 4384 15552
rect 30193 15555 30251 15561
rect 2700 15493 2728 15524
rect 30193 15521 30205 15555
rect 30239 15552 30251 15555
rect 30282 15552 30288 15564
rect 30239 15524 30288 15552
rect 30239 15521 30251 15524
rect 30193 15515 30251 15521
rect 30282 15512 30288 15524
rect 30340 15552 30346 15564
rect 30929 15555 30987 15561
rect 30929 15552 30941 15555
rect 30340 15524 30941 15552
rect 30340 15512 30346 15524
rect 30929 15521 30941 15524
rect 30975 15521 30987 15555
rect 30929 15515 30987 15521
rect 2685 15487 2743 15493
rect 2685 15453 2697 15487
rect 2731 15453 2743 15487
rect 2685 15447 2743 15453
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 3620 15416 3648 15447
rect 3786 15444 3792 15496
rect 3844 15444 3850 15496
rect 4433 15487 4491 15493
rect 4433 15453 4445 15487
rect 4479 15484 4491 15487
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 4479 15456 5089 15484
rect 4479 15453 4491 15456
rect 4433 15447 4491 15453
rect 5077 15453 5089 15456
rect 5123 15453 5135 15487
rect 5077 15447 5135 15453
rect 7558 15444 7564 15496
rect 7616 15484 7622 15496
rect 10594 15484 10600 15496
rect 7616 15456 10600 15484
rect 7616 15444 7622 15456
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 30834 15444 30840 15496
rect 30892 15444 30898 15496
rect 31662 15444 31668 15496
rect 31720 15444 31726 15496
rect 31754 15444 31760 15496
rect 31812 15484 31818 15496
rect 31921 15487 31979 15493
rect 31921 15484 31933 15487
rect 31812 15456 31933 15484
rect 31812 15444 31818 15456
rect 31921 15453 31933 15456
rect 31967 15453 31979 15487
rect 31921 15447 31979 15453
rect 3970 15416 3976 15428
rect 3620 15388 3976 15416
rect 3970 15376 3976 15388
rect 4028 15416 4034 15428
rect 4525 15419 4583 15425
rect 4525 15416 4537 15419
rect 4028 15388 4537 15416
rect 4028 15376 4034 15388
rect 4525 15385 4537 15388
rect 4571 15385 4583 15419
rect 4525 15379 4583 15385
rect 24578 15376 24584 15428
rect 24636 15416 24642 15428
rect 25222 15416 25228 15428
rect 24636 15388 25228 15416
rect 24636 15376 24642 15388
rect 25222 15376 25228 15388
rect 25280 15416 25286 15428
rect 25317 15419 25375 15425
rect 25317 15416 25329 15419
rect 25280 15388 25329 15416
rect 25280 15376 25286 15388
rect 25317 15385 25329 15388
rect 25363 15385 25375 15419
rect 25317 15379 25375 15385
rect 2958 15308 2964 15360
rect 3016 15308 3022 15360
rect 31570 15308 31576 15360
rect 31628 15308 31634 15360
rect 33042 15308 33048 15360
rect 33100 15308 33106 15360
rect 1104 15258 34016 15280
rect 1104 15206 9138 15258
rect 9190 15206 9202 15258
rect 9254 15206 9266 15258
rect 9318 15206 9330 15258
rect 9382 15206 9394 15258
rect 9446 15206 17326 15258
rect 17378 15206 17390 15258
rect 17442 15206 17454 15258
rect 17506 15206 17518 15258
rect 17570 15206 17582 15258
rect 17634 15206 25514 15258
rect 25566 15206 25578 15258
rect 25630 15206 25642 15258
rect 25694 15206 25706 15258
rect 25758 15206 25770 15258
rect 25822 15206 33702 15258
rect 33754 15206 33766 15258
rect 33818 15206 33830 15258
rect 33882 15206 33894 15258
rect 33946 15206 33958 15258
rect 34010 15206 34016 15258
rect 1104 15184 34016 15206
rect 3329 15147 3387 15153
rect 3329 15113 3341 15147
rect 3375 15144 3387 15147
rect 3786 15144 3792 15156
rect 3375 15116 3792 15144
rect 3375 15113 3387 15116
rect 3329 15107 3387 15113
rect 3786 15104 3792 15116
rect 3844 15104 3850 15156
rect 20165 15147 20223 15153
rect 20165 15113 20177 15147
rect 20211 15144 20223 15147
rect 24578 15144 24584 15156
rect 20211 15116 24584 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 18141 15079 18199 15085
rect 1964 15048 3648 15076
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 1964 14949 1992 15048
rect 3620 15017 3648 15048
rect 18141 15045 18153 15079
rect 18187 15076 18199 15079
rect 18506 15076 18512 15088
rect 18187 15048 18512 15076
rect 18187 15045 18199 15048
rect 18141 15039 18199 15045
rect 18506 15036 18512 15048
rect 18564 15076 18570 15088
rect 18969 15079 19027 15085
rect 18969 15076 18981 15079
rect 18564 15048 18981 15076
rect 18564 15036 18570 15048
rect 18969 15045 18981 15048
rect 19015 15076 19027 15079
rect 19337 15079 19395 15085
rect 19337 15076 19349 15079
rect 19015 15048 19349 15076
rect 19015 15045 19027 15048
rect 18969 15039 19027 15045
rect 19337 15045 19349 15048
rect 19383 15076 19395 15079
rect 20180 15076 20208 15107
rect 24578 15104 24584 15116
rect 24636 15104 24642 15156
rect 30834 15104 30840 15156
rect 30892 15144 30898 15156
rect 31297 15147 31355 15153
rect 31297 15144 31309 15147
rect 30892 15116 31309 15144
rect 30892 15104 30898 15116
rect 31297 15113 31309 15116
rect 31343 15113 31355 15147
rect 31297 15107 31355 15113
rect 19383 15048 20208 15076
rect 19383 15045 19395 15048
rect 19337 15039 19395 15045
rect 32306 15036 32312 15088
rect 32364 15076 32370 15088
rect 32585 15079 32643 15085
rect 32585 15076 32597 15079
rect 32364 15048 32597 15076
rect 32364 15036 32370 15048
rect 32585 15045 32597 15048
rect 32631 15045 32643 15079
rect 32585 15039 32643 15045
rect 2216 15011 2274 15017
rect 2216 14977 2228 15011
rect 2262 15008 2274 15011
rect 3605 15011 3663 15017
rect 2262 14980 3464 15008
rect 2262 14977 2274 14980
rect 2216 14971 2274 14977
rect 1949 14943 2007 14949
rect 1949 14940 1961 14943
rect 1820 14912 1961 14940
rect 1820 14900 1826 14912
rect 1949 14909 1961 14912
rect 1995 14909 2007 14943
rect 1949 14903 2007 14909
rect 3436 14804 3464 14980
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 3694 14968 3700 15020
rect 3752 15008 3758 15020
rect 3861 15011 3919 15017
rect 3861 15008 3873 15011
rect 3752 14980 3873 15008
rect 3752 14968 3758 14980
rect 3861 14977 3873 14980
rect 3907 14977 3919 15011
rect 3861 14971 3919 14977
rect 11606 14968 11612 15020
rect 11664 15008 11670 15020
rect 13981 15011 14039 15017
rect 13981 15008 13993 15011
rect 11664 14980 13993 15008
rect 11664 14968 11670 14980
rect 13981 14977 13993 14980
rect 14027 14977 14039 15011
rect 20714 15008 20720 15020
rect 13981 14971 14039 14977
rect 18432 14980 20720 15008
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 12768 14912 13737 14940
rect 12768 14900 12774 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 18432 14881 18460 14980
rect 20714 14968 20720 14980
rect 20772 14968 20778 15020
rect 31570 14968 31576 15020
rect 31628 15008 31634 15020
rect 32217 15011 32275 15017
rect 32217 15008 32229 15011
rect 31628 14980 32229 15008
rect 31628 14968 31634 14980
rect 32217 14977 32229 14980
rect 32263 14977 32275 15011
rect 32217 14971 32275 14977
rect 33042 14968 33048 15020
rect 33100 14968 33106 15020
rect 30009 14943 30067 14949
rect 30009 14909 30021 14943
rect 30055 14940 30067 14943
rect 30374 14940 30380 14952
rect 30055 14912 30380 14940
rect 30055 14909 30067 14912
rect 30009 14903 30067 14909
rect 18417 14875 18475 14881
rect 18417 14841 18429 14875
rect 18463 14841 18475 14875
rect 19705 14875 19763 14881
rect 18417 14835 18475 14841
rect 18524 14844 19564 14872
rect 4338 14804 4344 14816
rect 3436 14776 4344 14804
rect 4338 14764 4344 14776
rect 4396 14764 4402 14816
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5442 14804 5448 14816
rect 5031 14776 5448 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 15105 14807 15163 14813
rect 15105 14773 15117 14807
rect 15151 14804 15163 14807
rect 18524 14804 18552 14844
rect 19536 14816 19564 14844
rect 19705 14841 19717 14875
rect 19751 14872 19763 14875
rect 23474 14872 23480 14884
rect 19751 14844 23480 14872
rect 19751 14841 19763 14844
rect 19705 14835 19763 14841
rect 23474 14832 23480 14844
rect 23532 14832 23538 14884
rect 30024 14816 30052 14903
rect 30374 14900 30380 14912
rect 30432 14900 30438 14952
rect 30558 14900 30564 14952
rect 30616 14900 30622 14952
rect 31941 14943 31999 14949
rect 31941 14909 31953 14943
rect 31987 14940 31999 14943
rect 33060 14940 33088 14968
rect 31987 14912 33088 14940
rect 31987 14909 31999 14912
rect 31941 14903 31999 14909
rect 30282 14832 30288 14884
rect 30340 14832 30346 14884
rect 30469 14875 30527 14881
rect 30469 14841 30481 14875
rect 30515 14872 30527 14875
rect 31754 14872 31760 14884
rect 30515 14844 31760 14872
rect 30515 14841 30527 14844
rect 30469 14835 30527 14841
rect 31754 14832 31760 14844
rect 31812 14832 31818 14884
rect 15151 14776 18552 14804
rect 15151 14773 15163 14776
rect 15105 14767 15163 14773
rect 18598 14764 18604 14816
rect 18656 14764 18662 14816
rect 19518 14764 19524 14816
rect 19576 14764 19582 14816
rect 19794 14764 19800 14816
rect 19852 14764 19858 14816
rect 29917 14807 29975 14813
rect 29917 14773 29929 14807
rect 29963 14804 29975 14807
rect 30006 14804 30012 14816
rect 29963 14776 30012 14804
rect 29963 14773 29975 14776
rect 29917 14767 29975 14773
rect 30006 14764 30012 14776
rect 30064 14764 30070 14816
rect 31205 14807 31263 14813
rect 31205 14773 31217 14807
rect 31251 14804 31263 14807
rect 31294 14804 31300 14816
rect 31251 14776 31300 14804
rect 31251 14773 31263 14776
rect 31205 14767 31263 14773
rect 31294 14764 31300 14776
rect 31352 14764 31358 14816
rect 1104 14714 33856 14736
rect 1104 14662 5044 14714
rect 5096 14662 5108 14714
rect 5160 14662 5172 14714
rect 5224 14662 5236 14714
rect 5288 14662 5300 14714
rect 5352 14662 13232 14714
rect 13284 14662 13296 14714
rect 13348 14662 13360 14714
rect 13412 14662 13424 14714
rect 13476 14662 13488 14714
rect 13540 14662 21420 14714
rect 21472 14662 21484 14714
rect 21536 14662 21548 14714
rect 21600 14662 21612 14714
rect 21664 14662 21676 14714
rect 21728 14662 29608 14714
rect 29660 14662 29672 14714
rect 29724 14662 29736 14714
rect 29788 14662 29800 14714
rect 29852 14662 29864 14714
rect 29916 14662 33856 14714
rect 1104 14640 33856 14662
rect 3694 14560 3700 14612
rect 3752 14600 3758 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3752 14572 3801 14600
rect 3752 14560 3758 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 3789 14563 3847 14569
rect 4338 14560 4344 14612
rect 4396 14560 4402 14612
rect 11606 14560 11612 14612
rect 11664 14560 11670 14612
rect 18506 14560 18512 14612
rect 18564 14560 18570 14612
rect 18598 14560 18604 14612
rect 18656 14560 18662 14612
rect 19061 14603 19119 14609
rect 19061 14569 19073 14603
rect 19107 14600 19119 14603
rect 19150 14600 19156 14612
rect 19107 14572 19156 14600
rect 19107 14569 19119 14572
rect 19061 14563 19119 14569
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 3970 14492 3976 14544
rect 4028 14492 4034 14544
rect 4430 14492 4436 14544
rect 4488 14492 4494 14544
rect 11422 14492 11428 14544
rect 11480 14492 11486 14544
rect 1578 14424 1584 14476
rect 1636 14424 1642 14476
rect 3418 14424 3424 14476
rect 3476 14424 3482 14476
rect 2590 14356 2596 14408
rect 2648 14356 2654 14408
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14328 4307 14331
rect 4798 14328 4804 14340
rect 4295 14300 4804 14328
rect 4295 14297 4307 14300
rect 4249 14291 4307 14297
rect 4798 14288 4804 14300
rect 4856 14328 4862 14340
rect 5169 14331 5227 14337
rect 5169 14328 5181 14331
rect 4856 14300 5181 14328
rect 4856 14288 4862 14300
rect 5169 14297 5181 14300
rect 5215 14328 5227 14331
rect 5537 14331 5595 14337
rect 5537 14328 5549 14331
rect 5215 14300 5549 14328
rect 5215 14297 5227 14300
rect 5169 14291 5227 14297
rect 5537 14297 5549 14300
rect 5583 14297 5595 14331
rect 5537 14291 5595 14297
rect 11149 14331 11207 14337
rect 11149 14297 11161 14331
rect 11195 14328 11207 14331
rect 18524 14328 18552 14560
rect 18616 14396 18644 14560
rect 18874 14492 18880 14544
rect 18932 14492 18938 14544
rect 20625 14535 20683 14541
rect 20625 14501 20637 14535
rect 20671 14532 20683 14535
rect 24394 14532 24400 14544
rect 20671 14504 24400 14532
rect 20671 14501 20683 14504
rect 20625 14495 20683 14501
rect 24394 14492 24400 14504
rect 24452 14492 24458 14544
rect 31113 14467 31171 14473
rect 31113 14433 31125 14467
rect 31159 14433 31171 14467
rect 31113 14427 31171 14433
rect 19245 14399 19303 14405
rect 18616 14368 19104 14396
rect 18601 14331 18659 14337
rect 18601 14328 18613 14331
rect 11195 14300 12020 14328
rect 18524 14300 18613 14328
rect 11195 14297 11207 14300
rect 11149 14291 11207 14297
rect 11992 14272 12020 14300
rect 18601 14297 18613 14300
rect 18647 14297 18659 14331
rect 19076 14328 19104 14368
rect 19245 14365 19257 14399
rect 19291 14396 19303 14399
rect 19291 14368 21036 14396
rect 19291 14365 19303 14368
rect 19245 14359 19303 14365
rect 19490 14331 19548 14337
rect 19490 14328 19502 14331
rect 19076 14300 19502 14328
rect 18601 14291 18659 14297
rect 19490 14297 19502 14300
rect 19536 14297 19548 14331
rect 19490 14291 19548 14297
rect 21008 14272 21036 14368
rect 31128 14340 31156 14427
rect 31662 14424 31668 14476
rect 31720 14424 31726 14476
rect 31570 14356 31576 14408
rect 31628 14356 31634 14408
rect 31754 14356 31760 14408
rect 31812 14396 31818 14408
rect 31921 14399 31979 14405
rect 31921 14396 31933 14399
rect 31812 14368 31933 14396
rect 31812 14356 31818 14368
rect 31921 14365 31933 14368
rect 31967 14365 31979 14399
rect 31921 14359 31979 14365
rect 31110 14288 31116 14340
rect 31168 14288 31174 14340
rect 2866 14220 2872 14272
rect 2924 14220 2930 14272
rect 11974 14220 11980 14272
rect 12032 14220 12038 14272
rect 20990 14220 20996 14272
rect 21048 14220 21054 14272
rect 31018 14220 31024 14272
rect 31076 14260 31082 14272
rect 33045 14263 33103 14269
rect 33045 14260 33057 14263
rect 31076 14232 33057 14260
rect 31076 14220 31082 14232
rect 33045 14229 33057 14232
rect 33091 14229 33103 14263
rect 33045 14223 33103 14229
rect 1104 14170 34016 14192
rect 1104 14118 9138 14170
rect 9190 14118 9202 14170
rect 9254 14118 9266 14170
rect 9318 14118 9330 14170
rect 9382 14118 9394 14170
rect 9446 14118 17326 14170
rect 17378 14118 17390 14170
rect 17442 14118 17454 14170
rect 17506 14118 17518 14170
rect 17570 14118 17582 14170
rect 17634 14118 25514 14170
rect 25566 14118 25578 14170
rect 25630 14118 25642 14170
rect 25694 14118 25706 14170
rect 25758 14118 25770 14170
rect 25822 14118 33702 14170
rect 33754 14118 33766 14170
rect 33818 14118 33830 14170
rect 33882 14118 33894 14170
rect 33946 14118 33958 14170
rect 34010 14118 34016 14170
rect 1104 14096 34016 14118
rect 2590 14016 2596 14068
rect 2648 14016 2654 14068
rect 2958 14056 2964 14068
rect 2700 14028 2964 14056
rect 2317 13991 2375 13997
rect 2317 13957 2329 13991
rect 2363 13988 2375 13991
rect 2608 13988 2636 14016
rect 2363 13960 2636 13988
rect 2363 13957 2375 13960
rect 2317 13951 2375 13957
rect 2700 13929 2728 14028
rect 2958 14016 2964 14028
rect 3016 14016 3022 14068
rect 18877 14059 18935 14065
rect 18877 14025 18889 14059
rect 18923 14056 18935 14059
rect 19334 14056 19340 14068
rect 18923 14028 19340 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 19794 14016 19800 14068
rect 19852 14016 19858 14068
rect 30558 14016 30564 14068
rect 30616 14016 30622 14068
rect 19812 13988 19840 14016
rect 19990 13991 20048 13997
rect 19990 13988 20002 13991
rect 19812 13960 20002 13988
rect 19990 13957 20002 13960
rect 20036 13957 20048 13991
rect 19990 13951 20048 13957
rect 31570 13948 31576 14000
rect 31628 13988 31634 14000
rect 32585 13991 32643 13997
rect 32585 13988 32597 13991
rect 31628 13960 32597 13988
rect 31628 13948 31634 13960
rect 32585 13957 32597 13960
rect 32631 13957 32643 13991
rect 32585 13951 32643 13957
rect 2685 13923 2743 13929
rect 2685 13889 2697 13923
rect 2731 13889 2743 13923
rect 2685 13883 2743 13889
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 2869 13923 2927 13929
rect 2869 13920 2881 13923
rect 2832 13892 2881 13920
rect 2832 13880 2838 13892
rect 2869 13889 2881 13892
rect 2915 13889 2927 13923
rect 2869 13883 2927 13889
rect 20257 13923 20315 13929
rect 20257 13889 20269 13923
rect 20303 13920 20315 13923
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20303 13892 20637 13920
rect 20303 13889 20315 13892
rect 20257 13883 20315 13889
rect 20625 13889 20637 13892
rect 20671 13920 20683 13923
rect 20990 13920 20996 13932
rect 20671 13892 20996 13920
rect 20671 13889 20683 13892
rect 20625 13883 20683 13889
rect 20990 13880 20996 13892
rect 21048 13920 21054 13932
rect 22002 13920 22008 13932
rect 21048 13892 22008 13920
rect 21048 13880 21054 13892
rect 22002 13880 22008 13892
rect 22060 13920 22066 13932
rect 26510 13920 26516 13932
rect 22060 13892 26516 13920
rect 22060 13880 22066 13892
rect 26510 13880 26516 13892
rect 26568 13920 26574 13932
rect 31202 13920 31208 13932
rect 26568 13892 31208 13920
rect 26568 13880 26574 13892
rect 31202 13880 31208 13892
rect 31260 13880 31266 13932
rect 31941 13923 31999 13929
rect 31941 13889 31953 13923
rect 31987 13920 31999 13923
rect 32217 13923 32275 13929
rect 32217 13920 32229 13923
rect 31987 13892 32229 13920
rect 31987 13889 31999 13892
rect 31941 13883 31999 13889
rect 32217 13889 32229 13892
rect 32263 13889 32275 13923
rect 32217 13883 32275 13889
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 3329 13855 3387 13861
rect 3329 13852 3341 13855
rect 1360 13824 3341 13852
rect 1360 13812 1366 13824
rect 3329 13821 3341 13824
rect 3375 13821 3387 13855
rect 3329 13815 3387 13821
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 4433 13787 4491 13793
rect 4433 13784 4445 13787
rect 3476 13756 4445 13784
rect 3476 13744 3482 13756
rect 4433 13753 4445 13756
rect 4479 13753 4491 13787
rect 4433 13747 4491 13753
rect 4816 13728 4844 13815
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 15930 13852 15936 13864
rect 13688 13824 15936 13852
rect 13688 13812 13694 13824
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 29917 13855 29975 13861
rect 29917 13821 29929 13855
rect 29963 13852 29975 13855
rect 30006 13852 30012 13864
rect 29963 13824 30012 13852
rect 29963 13821 29975 13824
rect 29917 13815 29975 13821
rect 30006 13812 30012 13824
rect 30064 13852 30070 13864
rect 30558 13852 30564 13864
rect 30064 13824 30564 13852
rect 30064 13812 30070 13824
rect 30558 13812 30564 13824
rect 30616 13812 30622 13864
rect 31018 13812 31024 13864
rect 31076 13852 31082 13864
rect 31113 13855 31171 13861
rect 31113 13852 31125 13855
rect 31076 13824 31125 13852
rect 31076 13812 31082 13824
rect 31113 13821 31125 13824
rect 31159 13821 31171 13855
rect 31294 13852 31300 13864
rect 31255 13824 31300 13852
rect 31113 13815 31171 13821
rect 31294 13812 31300 13824
rect 31352 13812 31358 13864
rect 30377 13787 30435 13793
rect 30377 13753 30389 13787
rect 30423 13784 30435 13787
rect 31312 13784 31340 13812
rect 30423 13756 31340 13784
rect 30423 13753 30435 13756
rect 30377 13747 30435 13753
rect 4338 13676 4344 13728
rect 4396 13676 4402 13728
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 5077 13719 5135 13725
rect 5077 13716 5089 13719
rect 4856 13688 5089 13716
rect 4856 13676 4862 13688
rect 5077 13685 5089 13688
rect 5123 13685 5135 13719
rect 5077 13679 5135 13685
rect 30469 13719 30527 13725
rect 30469 13685 30481 13719
rect 30515 13716 30527 13719
rect 31754 13716 31760 13728
rect 30515 13688 31760 13716
rect 30515 13685 30527 13688
rect 30469 13679 30527 13685
rect 31754 13676 31760 13688
rect 31812 13676 31818 13728
rect 1104 13626 33856 13648
rect 1104 13574 5044 13626
rect 5096 13574 5108 13626
rect 5160 13574 5172 13626
rect 5224 13574 5236 13626
rect 5288 13574 5300 13626
rect 5352 13574 13232 13626
rect 13284 13574 13296 13626
rect 13348 13574 13360 13626
rect 13412 13574 13424 13626
rect 13476 13574 13488 13626
rect 13540 13574 21420 13626
rect 21472 13574 21484 13626
rect 21536 13574 21548 13626
rect 21600 13574 21612 13626
rect 21664 13574 21676 13626
rect 21728 13574 29608 13626
rect 29660 13574 29672 13626
rect 29724 13574 29736 13626
rect 29788 13574 29800 13626
rect 29852 13574 29864 13626
rect 29916 13574 33856 13626
rect 1104 13552 33856 13574
rect 33045 13515 33103 13521
rect 33045 13512 33057 13515
rect 31036 13484 33057 13512
rect 10594 13404 10600 13456
rect 10652 13404 10658 13456
rect 2409 13379 2467 13385
rect 2409 13345 2421 13379
rect 2455 13376 2467 13379
rect 2774 13376 2780 13388
rect 2455 13348 2780 13376
rect 2455 13345 2467 13348
rect 2409 13339 2467 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 4430 13336 4436 13388
rect 4488 13336 4494 13388
rect 31036 13385 31064 13484
rect 33045 13481 33057 13484
rect 33091 13481 33103 13515
rect 33045 13475 33103 13481
rect 31021 13379 31079 13385
rect 31021 13345 31033 13379
rect 31067 13345 31079 13379
rect 31021 13339 31079 13345
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13308 2743 13311
rect 2866 13308 2872 13320
rect 2731 13280 2872 13308
rect 2731 13277 2743 13280
rect 2685 13271 2743 13277
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 4246 13308 4252 13320
rect 3559 13280 4252 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 4246 13268 4252 13280
rect 4304 13268 4310 13320
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 19702 13308 19708 13320
rect 19484 13280 19708 13308
rect 19484 13268 19490 13280
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 30285 13311 30343 13317
rect 30285 13277 30297 13311
rect 30331 13308 30343 13311
rect 30926 13308 30932 13320
rect 30331 13280 30932 13308
rect 30331 13277 30343 13280
rect 30285 13271 30343 13277
rect 30926 13268 30932 13280
rect 30984 13268 30990 13320
rect 31202 13268 31208 13320
rect 31260 13308 31266 13320
rect 31665 13311 31723 13317
rect 31665 13308 31677 13311
rect 31260 13280 31677 13308
rect 31260 13268 31266 13280
rect 31665 13277 31677 13280
rect 31711 13277 31723 13311
rect 31665 13271 31723 13277
rect 31754 13268 31760 13320
rect 31812 13308 31818 13320
rect 31921 13311 31979 13317
rect 31921 13308 31933 13311
rect 31812 13280 31933 13308
rect 31812 13268 31818 13280
rect 31921 13277 31933 13280
rect 31967 13277 31979 13311
rect 31921 13271 31979 13277
rect 10965 13243 11023 13249
rect 10965 13209 10977 13243
rect 11011 13240 11023 13243
rect 11011 13212 11376 13240
rect 11011 13209 11023 13212
rect 10965 13203 11023 13209
rect 2866 13132 2872 13184
rect 2924 13132 2930 13184
rect 3418 13132 3424 13184
rect 3476 13172 3482 13184
rect 3789 13175 3847 13181
rect 3789 13172 3801 13175
rect 3476 13144 3801 13172
rect 3476 13132 3482 13144
rect 3789 13141 3801 13144
rect 3835 13141 3847 13175
rect 3789 13135 3847 13141
rect 10505 13175 10563 13181
rect 10505 13141 10517 13175
rect 10551 13172 10563 13175
rect 11146 13172 11152 13184
rect 10551 13144 11152 13172
rect 10551 13141 10563 13144
rect 10505 13135 10563 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11348 13181 11376 13212
rect 11333 13175 11391 13181
rect 11333 13141 11345 13175
rect 11379 13172 11391 13175
rect 11974 13172 11980 13184
rect 11379 13144 11980 13172
rect 11379 13141 11391 13144
rect 11333 13135 11391 13141
rect 11974 13132 11980 13144
rect 12032 13172 12038 13184
rect 13630 13172 13636 13184
rect 12032 13144 13636 13172
rect 12032 13132 12038 13144
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13172 20039 13175
rect 20346 13172 20352 13184
rect 20027 13144 20352 13172
rect 20027 13141 20039 13144
rect 19981 13135 20039 13141
rect 20346 13132 20352 13144
rect 20404 13132 20410 13184
rect 30834 13132 30840 13184
rect 30892 13132 30898 13184
rect 31570 13132 31576 13184
rect 31628 13132 31634 13184
rect 1104 13082 34016 13104
rect 1104 13030 9138 13082
rect 9190 13030 9202 13082
rect 9254 13030 9266 13082
rect 9318 13030 9330 13082
rect 9382 13030 9394 13082
rect 9446 13030 17326 13082
rect 17378 13030 17390 13082
rect 17442 13030 17454 13082
rect 17506 13030 17518 13082
rect 17570 13030 17582 13082
rect 17634 13030 25514 13082
rect 25566 13030 25578 13082
rect 25630 13030 25642 13082
rect 25694 13030 25706 13082
rect 25758 13030 25770 13082
rect 25822 13030 33702 13082
rect 33754 13030 33766 13082
rect 33818 13030 33830 13082
rect 33882 13030 33894 13082
rect 33946 13030 33958 13082
rect 34010 13030 34016 13082
rect 1104 13008 34016 13030
rect 4246 12928 4252 12980
rect 4304 12968 4310 12980
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 4304 12940 4629 12968
rect 4304 12928 4310 12940
rect 4617 12937 4629 12940
rect 4663 12937 4675 12971
rect 4617 12931 4675 12937
rect 23474 12928 23480 12980
rect 23532 12928 23538 12980
rect 31202 12928 31208 12980
rect 31260 12928 31266 12980
rect 2032 12903 2090 12909
rect 2032 12869 2044 12903
rect 2078 12900 2090 12903
rect 4338 12900 4344 12912
rect 2078 12872 4344 12900
rect 2078 12869 2090 12872
rect 2032 12863 2090 12869
rect 4338 12860 4344 12872
rect 4396 12860 4402 12912
rect 4430 12860 4436 12912
rect 4488 12860 4494 12912
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12832 3387 12835
rect 3510 12832 3516 12844
rect 3375 12804 3516 12832
rect 3375 12801 3387 12804
rect 3329 12795 3387 12801
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 3881 12835 3939 12841
rect 3881 12801 3893 12835
rect 3927 12832 3939 12835
rect 4448 12832 4476 12860
rect 23492 12841 23520 12928
rect 30852 12872 32260 12900
rect 30852 12844 30880 12872
rect 3927 12804 4476 12832
rect 23477 12835 23535 12841
rect 3927 12801 3939 12804
rect 3881 12795 3939 12801
rect 23477 12801 23489 12835
rect 23523 12832 23535 12835
rect 26970 12832 26976 12844
rect 23523 12804 26976 12832
rect 23523 12801 23535 12804
rect 23477 12795 23535 12801
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 30834 12792 30840 12844
rect 30892 12792 30898 12844
rect 30926 12792 30932 12844
rect 30984 12832 30990 12844
rect 31297 12835 31355 12841
rect 31297 12832 31309 12835
rect 30984 12804 31309 12832
rect 30984 12792 30990 12804
rect 31297 12801 31309 12804
rect 31343 12801 31355 12835
rect 31297 12795 31355 12801
rect 31570 12792 31576 12844
rect 31628 12832 31634 12844
rect 32232 12841 32260 12872
rect 31849 12835 31907 12841
rect 31849 12832 31861 12835
rect 31628 12804 31861 12832
rect 31628 12792 31634 12804
rect 31849 12801 31861 12804
rect 31895 12801 31907 12835
rect 31849 12795 31907 12801
rect 32217 12835 32275 12841
rect 32217 12801 32229 12835
rect 32263 12801 32275 12835
rect 32217 12795 32275 12801
rect 1762 12724 1768 12776
rect 1820 12724 1826 12776
rect 3970 12724 3976 12776
rect 4028 12724 4034 12776
rect 32490 12724 32496 12776
rect 32548 12724 32554 12776
rect 3142 12588 3148 12640
rect 3200 12588 3206 12640
rect 4798 12588 4804 12640
rect 4856 12628 4862 12640
rect 5077 12631 5135 12637
rect 5077 12628 5089 12631
rect 4856 12600 5089 12628
rect 4856 12588 4862 12600
rect 5077 12597 5089 12600
rect 5123 12597 5135 12631
rect 5077 12591 5135 12597
rect 23658 12588 23664 12640
rect 23716 12588 23722 12640
rect 1104 12538 33856 12560
rect 1104 12486 5044 12538
rect 5096 12486 5108 12538
rect 5160 12486 5172 12538
rect 5224 12486 5236 12538
rect 5288 12486 5300 12538
rect 5352 12486 13232 12538
rect 13284 12486 13296 12538
rect 13348 12486 13360 12538
rect 13412 12486 13424 12538
rect 13476 12486 13488 12538
rect 13540 12486 21420 12538
rect 21472 12486 21484 12538
rect 21536 12486 21548 12538
rect 21600 12486 21612 12538
rect 21664 12486 21676 12538
rect 21728 12486 29608 12538
rect 29660 12486 29672 12538
rect 29724 12486 29736 12538
rect 29788 12486 29800 12538
rect 29852 12486 29864 12538
rect 29916 12486 33856 12538
rect 1104 12464 33856 12486
rect 3513 12427 3571 12433
rect 3513 12393 3525 12427
rect 3559 12424 3571 12427
rect 3970 12424 3976 12436
rect 3559 12396 3976 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 3970 12384 3976 12396
rect 4028 12384 4034 12436
rect 30558 12384 30564 12436
rect 30616 12424 30622 12436
rect 30653 12427 30711 12433
rect 30653 12424 30665 12427
rect 30616 12396 30665 12424
rect 30616 12384 30622 12396
rect 30653 12393 30665 12396
rect 30699 12393 30711 12427
rect 30653 12387 30711 12393
rect 4246 12316 4252 12368
rect 4304 12356 4310 12368
rect 4617 12359 4675 12365
rect 4617 12356 4629 12359
rect 4304 12328 4629 12356
rect 4304 12316 4310 12328
rect 4617 12325 4629 12328
rect 4663 12325 4675 12359
rect 4617 12319 4675 12325
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12288 3019 12291
rect 3142 12288 3148 12300
rect 3007 12260 3148 12288
rect 3007 12257 3019 12260
rect 2961 12251 3019 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 5442 12248 5448 12300
rect 5500 12248 5506 12300
rect 24394 12248 24400 12300
rect 24452 12248 24458 12300
rect 30668 12288 30696 12387
rect 30926 12316 30932 12368
rect 30984 12356 30990 12368
rect 31113 12359 31171 12365
rect 31113 12356 31125 12359
rect 30984 12328 31125 12356
rect 30984 12316 30990 12328
rect 31113 12325 31125 12328
rect 31159 12325 31171 12359
rect 31113 12319 31171 12325
rect 30837 12291 30895 12297
rect 30837 12288 30849 12291
rect 30668 12260 30849 12288
rect 30837 12257 30849 12260
rect 30883 12257 30895 12291
rect 30837 12251 30895 12257
rect 33318 12248 33324 12300
rect 33376 12248 33382 12300
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 2866 12220 2872 12232
rect 2731 12192 2872 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3786 12180 3792 12232
rect 3844 12180 3850 12232
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 11422 12220 11428 12232
rect 9548 12192 11428 12220
rect 9548 12180 9554 12192
rect 11422 12180 11428 12192
rect 11480 12180 11486 12232
rect 32030 12180 32036 12232
rect 32088 12180 32094 12232
rect 32309 12223 32367 12229
rect 32309 12189 32321 12223
rect 32355 12220 32367 12223
rect 32490 12220 32496 12232
rect 32355 12192 32496 12220
rect 32355 12189 32367 12192
rect 32309 12183 32367 12189
rect 32490 12180 32496 12192
rect 32548 12180 32554 12232
rect 2317 12155 2375 12161
rect 2317 12121 2329 12155
rect 2363 12152 2375 12155
rect 2363 12124 2636 12152
rect 2363 12121 2375 12124
rect 2317 12115 2375 12121
rect 2608 12096 2636 12124
rect 4798 12112 4804 12164
rect 4856 12152 4862 12164
rect 4985 12155 5043 12161
rect 4985 12152 4997 12155
rect 4856 12124 4997 12152
rect 4856 12112 4862 12124
rect 4985 12121 4997 12124
rect 5031 12121 5043 12155
rect 4985 12115 5043 12121
rect 2590 12044 2596 12096
rect 2648 12044 2654 12096
rect 4430 12044 4436 12096
rect 4488 12044 4494 12096
rect 4522 12044 4528 12096
rect 4580 12044 4586 12096
rect 5994 12044 6000 12096
rect 6052 12044 6058 12096
rect 8938 12044 8944 12096
rect 8996 12044 9002 12096
rect 25038 12044 25044 12096
rect 25096 12044 25102 12096
rect 31294 12044 31300 12096
rect 31352 12044 31358 12096
rect 31386 12044 31392 12096
rect 31444 12044 31450 12096
rect 1104 11994 34016 12016
rect 1104 11942 9138 11994
rect 9190 11942 9202 11994
rect 9254 11942 9266 11994
rect 9318 11942 9330 11994
rect 9382 11942 9394 11994
rect 9446 11942 17326 11994
rect 17378 11942 17390 11994
rect 17442 11942 17454 11994
rect 17506 11942 17518 11994
rect 17570 11942 17582 11994
rect 17634 11942 25514 11994
rect 25566 11942 25578 11994
rect 25630 11942 25642 11994
rect 25694 11942 25706 11994
rect 25758 11942 25770 11994
rect 25822 11942 33702 11994
rect 33754 11942 33766 11994
rect 33818 11942 33830 11994
rect 33882 11942 33894 11994
rect 33946 11942 33958 11994
rect 34010 11942 34016 11994
rect 1104 11920 34016 11942
rect 4430 11840 4436 11892
rect 4488 11840 4494 11892
rect 32030 11840 32036 11892
rect 32088 11880 32094 11892
rect 33505 11883 33563 11889
rect 33505 11880 33517 11883
rect 32088 11852 33517 11880
rect 32088 11840 32094 11852
rect 33505 11849 33517 11852
rect 33551 11849 33563 11883
rect 33505 11843 33563 11849
rect 1578 11772 1584 11824
rect 1636 11772 1642 11824
rect 2590 11704 2596 11756
rect 2648 11704 2654 11756
rect 2866 11704 2872 11756
rect 2924 11704 2930 11756
rect 4448 11744 4476 11840
rect 11146 11772 11152 11824
rect 11204 11812 11210 11824
rect 12866 11815 12924 11821
rect 12866 11812 12878 11815
rect 11204 11784 12878 11812
rect 11204 11772 11210 11784
rect 12866 11781 12878 11784
rect 12912 11781 12924 11815
rect 12866 11775 12924 11781
rect 31294 11772 31300 11824
rect 31352 11812 31358 11824
rect 32370 11815 32428 11821
rect 32370 11812 32382 11815
rect 31352 11784 32382 11812
rect 31352 11772 31358 11784
rect 32370 11781 32382 11784
rect 32416 11781 32428 11815
rect 32370 11775 32428 11781
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4448 11716 4905 11744
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 12710 11744 12716 11756
rect 12667 11716 12716 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 12710 11704 12716 11716
rect 12768 11704 12774 11756
rect 19334 11704 19340 11756
rect 19392 11704 19398 11756
rect 31662 11704 31668 11756
rect 31720 11704 31726 11756
rect 31938 11704 31944 11756
rect 31996 11704 32002 11756
rect 1302 11636 1308 11688
rect 1360 11676 1366 11688
rect 3329 11679 3387 11685
rect 3329 11676 3341 11679
rect 1360 11648 3341 11676
rect 1360 11636 1366 11648
rect 3329 11645 3341 11648
rect 3375 11645 3387 11679
rect 3329 11639 3387 11645
rect 31478 11636 31484 11688
rect 31536 11636 31542 11688
rect 31680 11676 31708 11704
rect 32125 11679 32183 11685
rect 32125 11676 32137 11679
rect 31680 11648 32137 11676
rect 32125 11645 32137 11648
rect 32171 11645 32183 11679
rect 32125 11639 32183 11645
rect 4338 11500 4344 11552
rect 4396 11500 4402 11552
rect 14001 11543 14059 11549
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 15470 11540 15476 11552
rect 14047 11512 15476 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 19978 11500 19984 11552
rect 20036 11500 20042 11552
rect 1104 11450 33856 11472
rect 1104 11398 5044 11450
rect 5096 11398 5108 11450
rect 5160 11398 5172 11450
rect 5224 11398 5236 11450
rect 5288 11398 5300 11450
rect 5352 11398 13232 11450
rect 13284 11398 13296 11450
rect 13348 11398 13360 11450
rect 13412 11398 13424 11450
rect 13476 11398 13488 11450
rect 13540 11398 21420 11450
rect 21472 11398 21484 11450
rect 21536 11398 21548 11450
rect 21600 11398 21612 11450
rect 21664 11398 21676 11450
rect 21728 11398 29608 11450
rect 29660 11398 29672 11450
rect 29724 11398 29736 11450
rect 29788 11398 29800 11450
rect 29852 11398 29864 11450
rect 29916 11398 33856 11450
rect 1104 11376 33856 11398
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3786 11336 3792 11348
rect 3191 11308 3792 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4522 11296 4528 11348
rect 4580 11296 4586 11348
rect 30558 11296 30564 11348
rect 30616 11296 30622 11348
rect 31938 11296 31944 11348
rect 31996 11336 32002 11348
rect 31996 11308 32536 11336
rect 31996 11296 32002 11308
rect 4338 11160 4344 11212
rect 4396 11160 4402 11212
rect 1762 11092 1768 11144
rect 1820 11092 1826 11144
rect 2032 11135 2090 11141
rect 2032 11101 2044 11135
rect 2078 11132 2090 11135
rect 4540 11132 4568 11296
rect 31386 11160 31392 11212
rect 31444 11200 31450 11212
rect 32508 11209 32536 11308
rect 31941 11203 31999 11209
rect 31941 11200 31953 11203
rect 31444 11172 31953 11200
rect 31444 11160 31450 11172
rect 31941 11169 31953 11172
rect 31987 11169 31999 11203
rect 31941 11163 31999 11169
rect 32493 11203 32551 11209
rect 32493 11169 32505 11203
rect 32539 11169 32551 11203
rect 32493 11163 32551 11169
rect 2078 11104 4568 11132
rect 2078 11101 2090 11104
rect 2032 11095 2090 11101
rect 32214 11092 32220 11144
rect 32272 11092 32278 11144
rect 3786 10956 3792 11008
rect 3844 10956 3850 11008
rect 31386 10956 31392 11008
rect 31444 10956 31450 11008
rect 1104 10906 34016 10928
rect 1104 10854 9138 10906
rect 9190 10854 9202 10906
rect 9254 10854 9266 10906
rect 9318 10854 9330 10906
rect 9382 10854 9394 10906
rect 9446 10854 17326 10906
rect 17378 10854 17390 10906
rect 17442 10854 17454 10906
rect 17506 10854 17518 10906
rect 17570 10854 17582 10906
rect 17634 10854 25514 10906
rect 25566 10854 25578 10906
rect 25630 10854 25642 10906
rect 25694 10854 25706 10906
rect 25758 10854 25770 10906
rect 25822 10854 33702 10906
rect 33754 10854 33766 10906
rect 33818 10854 33830 10906
rect 33882 10854 33894 10906
rect 33946 10854 33958 10906
rect 34010 10854 34016 10906
rect 1104 10832 34016 10854
rect 9953 10795 10011 10801
rect 9953 10761 9965 10795
rect 9999 10792 10011 10795
rect 10318 10792 10324 10804
rect 9999 10764 10324 10792
rect 9999 10761 10011 10764
rect 9953 10755 10011 10761
rect 2317 10727 2375 10733
rect 2317 10693 2329 10727
rect 2363 10724 2375 10727
rect 2866 10724 2872 10736
rect 2363 10696 2872 10724
rect 2363 10693 2375 10696
rect 2317 10687 2375 10693
rect 2866 10684 2872 10696
rect 2924 10684 2930 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 9968 10724 9996 10755
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 31941 10795 31999 10801
rect 31941 10761 31953 10795
rect 31987 10792 31999 10795
rect 32214 10792 32220 10804
rect 31987 10764 32220 10792
rect 31987 10761 31999 10764
rect 31941 10755 31999 10761
rect 32214 10752 32220 10764
rect 32272 10752 32278 10804
rect 7892 10696 9996 10724
rect 30377 10727 30435 10733
rect 7892 10684 7898 10696
rect 30377 10693 30389 10727
rect 30423 10724 30435 10727
rect 31662 10724 31668 10736
rect 30423 10696 31668 10724
rect 30423 10693 30435 10696
rect 30377 10687 30435 10693
rect 31662 10684 31668 10696
rect 31720 10684 31726 10736
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 3786 10656 3792 10668
rect 2731 10628 3792 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 4614 10656 4620 10668
rect 4080 10628 4620 10656
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10588 3663 10591
rect 4080 10588 4108 10628
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 28629 10659 28687 10665
rect 28629 10656 28641 10659
rect 28460 10628 28641 10656
rect 3651 10560 4108 10588
rect 4157 10591 4215 10597
rect 3651 10557 3663 10560
rect 3605 10551 3663 10557
rect 4157 10557 4169 10591
rect 4203 10588 4215 10591
rect 4798 10588 4804 10600
rect 4203 10560 4804 10588
rect 4203 10557 4215 10560
rect 4157 10551 4215 10557
rect 3881 10523 3939 10529
rect 3881 10489 3893 10523
rect 3927 10520 3939 10523
rect 4338 10520 4344 10532
rect 3927 10492 4344 10520
rect 3927 10489 3939 10492
rect 3881 10483 3939 10489
rect 4338 10480 4344 10492
rect 4396 10480 4402 10532
rect 4448 10464 4476 10560
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 12710 10588 12716 10600
rect 9640 10560 12716 10588
rect 9640 10548 9646 10560
rect 12710 10548 12716 10560
rect 12768 10548 12774 10600
rect 2958 10412 2964 10464
rect 3016 10412 3022 10464
rect 3694 10412 3700 10464
rect 3752 10412 3758 10464
rect 4430 10412 4436 10464
rect 4488 10412 4494 10464
rect 27798 10412 27804 10464
rect 27856 10452 27862 10464
rect 28460 10461 28488 10628
rect 28629 10625 28641 10628
rect 28675 10625 28687 10659
rect 30558 10656 30564 10668
rect 28629 10619 28687 10625
rect 30346 10628 30564 10656
rect 30006 10548 30012 10600
rect 30064 10588 30070 10600
rect 30346 10588 30374 10628
rect 30558 10616 30564 10628
rect 30616 10656 30622 10668
rect 30745 10659 30803 10665
rect 30745 10656 30757 10659
rect 30616 10628 30757 10656
rect 30616 10616 30622 10628
rect 30745 10625 30757 10628
rect 30791 10625 30803 10659
rect 30745 10619 30803 10625
rect 31386 10616 31392 10668
rect 31444 10616 31450 10668
rect 32306 10616 32312 10668
rect 32364 10616 32370 10668
rect 30064 10560 30374 10588
rect 30064 10548 30070 10560
rect 31113 10523 31171 10529
rect 31113 10489 31125 10523
rect 31159 10520 31171 10523
rect 31404 10520 31432 10616
rect 33318 10548 33324 10600
rect 33376 10548 33382 10600
rect 31159 10492 31432 10520
rect 31159 10489 31171 10492
rect 31113 10483 31171 10489
rect 28445 10455 28503 10461
rect 28445 10452 28457 10455
rect 27856 10424 28457 10452
rect 27856 10412 27862 10424
rect 28445 10421 28457 10424
rect 28491 10421 28503 10455
rect 28445 10415 28503 10421
rect 31202 10412 31208 10464
rect 31260 10412 31266 10464
rect 1104 10362 33856 10384
rect 1104 10310 5044 10362
rect 5096 10310 5108 10362
rect 5160 10310 5172 10362
rect 5224 10310 5236 10362
rect 5288 10310 5300 10362
rect 5352 10310 13232 10362
rect 13284 10310 13296 10362
rect 13348 10310 13360 10362
rect 13412 10310 13424 10362
rect 13476 10310 13488 10362
rect 13540 10310 21420 10362
rect 21472 10310 21484 10362
rect 21536 10310 21548 10362
rect 21600 10310 21612 10362
rect 21664 10310 21676 10362
rect 21728 10310 29608 10362
rect 29660 10310 29672 10362
rect 29724 10310 29736 10362
rect 29788 10310 29800 10362
rect 29852 10310 29864 10362
rect 29916 10310 33856 10362
rect 1104 10288 33856 10310
rect 7377 10251 7435 10257
rect 7377 10217 7389 10251
rect 7423 10248 7435 10251
rect 7834 10248 7840 10260
rect 7423 10220 7840 10248
rect 7423 10217 7435 10220
rect 7377 10211 7435 10217
rect 5261 10115 5319 10121
rect 5261 10112 5273 10115
rect 2792 10084 5273 10112
rect 1762 10004 1768 10056
rect 1820 10044 1826 10056
rect 2792 10044 2820 10084
rect 5261 10081 5273 10084
rect 5307 10081 5319 10115
rect 5261 10075 5319 10081
rect 1820 10016 2820 10044
rect 1820 10004 1826 10016
rect 3694 10004 3700 10056
rect 3752 10004 3758 10056
rect 4338 10004 4344 10056
rect 4396 10004 4402 10056
rect 7009 10047 7067 10053
rect 7009 10013 7021 10047
rect 7055 10044 7067 10047
rect 7392 10044 7420 10211
rect 7834 10208 7840 10220
rect 7892 10208 7898 10260
rect 25866 10208 25872 10260
rect 25924 10208 25930 10260
rect 26510 10208 26516 10260
rect 26568 10208 26574 10260
rect 15470 10072 15476 10124
rect 15528 10072 15534 10124
rect 7055 10016 7420 10044
rect 25884 10044 25912 10208
rect 30193 10115 30251 10121
rect 30193 10081 30205 10115
rect 30239 10112 30251 10115
rect 30374 10112 30380 10124
rect 30239 10084 30380 10112
rect 30239 10081 30251 10084
rect 30193 10075 30251 10081
rect 30374 10072 30380 10084
rect 30432 10112 30438 10124
rect 30929 10115 30987 10121
rect 30929 10112 30941 10115
rect 30432 10084 30941 10112
rect 30432 10072 30438 10084
rect 30929 10081 30941 10084
rect 30975 10081 30987 10115
rect 30929 10075 30987 10081
rect 31662 10072 31668 10124
rect 31720 10072 31726 10124
rect 27798 10044 27804 10056
rect 25884 10016 27804 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 27798 10004 27804 10016
rect 27856 10004 27862 10056
rect 30834 10004 30840 10056
rect 30892 10004 30898 10056
rect 31202 10004 31208 10056
rect 31260 10044 31266 10056
rect 31921 10047 31979 10053
rect 31921 10044 31933 10047
rect 31260 10016 31933 10044
rect 31260 10004 31266 10016
rect 31921 10013 31933 10016
rect 31967 10013 31979 10047
rect 31921 10007 31979 10013
rect 2032 9979 2090 9985
rect 2032 9945 2044 9979
rect 2078 9976 2090 9979
rect 3712 9976 3740 10004
rect 2078 9948 3740 9976
rect 2078 9945 2090 9948
rect 2032 9939 2090 9945
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 3786 9868 3792 9920
rect 3844 9868 3850 9920
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16942 9908 16948 9920
rect 16163 9880 16948 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 31570 9868 31576 9920
rect 31628 9868 31634 9920
rect 33042 9868 33048 9920
rect 33100 9868 33106 9920
rect 1104 9818 34016 9840
rect 1104 9766 9138 9818
rect 9190 9766 9202 9818
rect 9254 9766 9266 9818
rect 9318 9766 9330 9818
rect 9382 9766 9394 9818
rect 9446 9766 17326 9818
rect 17378 9766 17390 9818
rect 17442 9766 17454 9818
rect 17506 9766 17518 9818
rect 17570 9766 17582 9818
rect 17634 9766 25514 9818
rect 25566 9766 25578 9818
rect 25630 9766 25642 9818
rect 25694 9766 25706 9818
rect 25758 9766 25770 9818
rect 25822 9766 33702 9818
rect 33754 9766 33766 9818
rect 33818 9766 33830 9818
rect 33882 9766 33894 9818
rect 33946 9766 33958 9818
rect 34010 9766 34016 9818
rect 1104 9744 34016 9766
rect 26970 9664 26976 9716
rect 27028 9664 27034 9716
rect 30834 9664 30840 9716
rect 30892 9704 30898 9716
rect 31297 9707 31355 9713
rect 31297 9704 31309 9707
rect 30892 9676 31309 9704
rect 30892 9664 30898 9676
rect 31297 9673 31309 9676
rect 31343 9673 31355 9707
rect 31297 9667 31355 9673
rect 1578 9596 1584 9648
rect 1636 9596 1642 9648
rect 32306 9596 32312 9648
rect 32364 9636 32370 9648
rect 32585 9639 32643 9645
rect 32585 9636 32597 9639
rect 32364 9608 32597 9636
rect 32364 9596 32370 9608
rect 32585 9605 32597 9608
rect 32631 9605 32643 9639
rect 32585 9599 32643 9605
rect 2590 9528 2596 9580
rect 2648 9528 2654 9580
rect 3142 9528 3148 9580
rect 3200 9568 3206 9580
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 3200 9540 3433 9568
rect 3200 9528 3206 9540
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4111 9540 4476 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4338 9460 4344 9512
rect 4396 9460 4402 9512
rect 3789 9435 3847 9441
rect 3789 9401 3801 9435
rect 3835 9432 3847 9435
rect 4356 9432 4384 9460
rect 3835 9404 4384 9432
rect 3835 9401 3847 9404
rect 3789 9395 3847 9401
rect 4448 9376 4476 9540
rect 24946 9528 24952 9580
rect 25004 9528 25010 9580
rect 25038 9528 25044 9580
rect 25096 9568 25102 9580
rect 27525 9571 27583 9577
rect 27525 9568 27537 9571
rect 25096 9540 27537 9568
rect 25096 9528 25102 9540
rect 27525 9537 27537 9540
rect 27571 9537 27583 9571
rect 27525 9531 27583 9537
rect 31570 9528 31576 9580
rect 31628 9568 31634 9580
rect 32217 9571 32275 9577
rect 32217 9568 32229 9571
rect 31628 9540 32229 9568
rect 31628 9528 31634 9540
rect 32217 9537 32229 9540
rect 32263 9537 32275 9571
rect 32217 9531 32275 9537
rect 33042 9528 33048 9580
rect 33100 9528 33106 9580
rect 15194 9460 15200 9512
rect 15252 9500 15258 9512
rect 18874 9500 18880 9512
rect 15252 9472 18880 9500
rect 15252 9460 15258 9472
rect 18874 9460 18880 9472
rect 18932 9460 18938 9512
rect 30006 9500 30012 9512
rect 29840 9472 30012 9500
rect 2866 9324 2872 9376
rect 2924 9324 2930 9376
rect 3602 9324 3608 9376
rect 3660 9324 3666 9376
rect 4430 9324 4436 9376
rect 4488 9324 4494 9376
rect 13906 9324 13912 9376
rect 13964 9364 13970 9376
rect 14645 9367 14703 9373
rect 14645 9364 14657 9367
rect 13964 9336 14657 9364
rect 13964 9324 13970 9336
rect 14645 9333 14657 9336
rect 14691 9333 14703 9367
rect 14645 9327 14703 9333
rect 23658 9324 23664 9376
rect 23716 9364 23722 9376
rect 24305 9367 24363 9373
rect 24305 9364 24317 9367
rect 23716 9336 24317 9364
rect 23716 9324 23722 9336
rect 24305 9333 24317 9336
rect 24351 9333 24363 9367
rect 24305 9327 24363 9333
rect 27614 9324 27620 9376
rect 27672 9364 27678 9376
rect 29840 9373 29868 9472
rect 30006 9460 30012 9472
rect 30064 9460 30070 9512
rect 31110 9460 31116 9512
rect 31168 9460 31174 9512
rect 31941 9503 31999 9509
rect 31941 9469 31953 9503
rect 31987 9500 31999 9503
rect 33060 9500 33088 9528
rect 31987 9472 33088 9500
rect 31987 9469 31999 9472
rect 31941 9463 31999 9469
rect 30374 9392 30380 9444
rect 30432 9392 30438 9444
rect 29825 9367 29883 9373
rect 29825 9364 29837 9367
rect 27672 9336 29837 9364
rect 27672 9324 27678 9336
rect 29825 9333 29837 9336
rect 29871 9333 29883 9367
rect 29825 9327 29883 9333
rect 30466 9324 30472 9376
rect 30524 9324 30530 9376
rect 30558 9324 30564 9376
rect 30616 9324 30622 9376
rect 1104 9274 33856 9296
rect 1104 9222 5044 9274
rect 5096 9222 5108 9274
rect 5160 9222 5172 9274
rect 5224 9222 5236 9274
rect 5288 9222 5300 9274
rect 5352 9222 13232 9274
rect 13284 9222 13296 9274
rect 13348 9222 13360 9274
rect 13412 9222 13424 9274
rect 13476 9222 13488 9274
rect 13540 9222 21420 9274
rect 21472 9222 21484 9274
rect 21536 9222 21548 9274
rect 21600 9222 21612 9274
rect 21664 9222 21676 9274
rect 21728 9222 29608 9274
rect 29660 9222 29672 9274
rect 29724 9222 29736 9274
rect 29788 9222 29800 9274
rect 29852 9222 29864 9274
rect 29916 9222 33856 9274
rect 1104 9200 33856 9222
rect 2590 9120 2596 9172
rect 2648 9120 2654 9172
rect 2866 9120 2872 9172
rect 2924 9120 2930 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 4338 9160 4344 9172
rect 3559 9132 4344 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 6181 9163 6239 9169
rect 6181 9129 6193 9163
rect 6227 9160 6239 9163
rect 9490 9160 9496 9172
rect 6227 9132 9496 9160
rect 6227 9129 6239 9132
rect 6181 9123 6239 9129
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 19702 9120 19708 9172
rect 19760 9120 19766 9172
rect 2409 9027 2467 9033
rect 2409 8993 2421 9027
rect 2455 9024 2467 9027
rect 2608 9024 2636 9120
rect 2884 9033 2912 9120
rect 2455 8996 2636 9024
rect 2869 9027 2927 9033
rect 2455 8993 2467 8996
rect 2409 8987 2467 8993
rect 2869 8993 2881 9027
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 5994 9024 6000 9036
rect 5675 8996 6000 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 5994 8984 6000 8996
rect 6052 8984 6058 9036
rect 19978 8984 19984 9036
rect 20036 9024 20042 9036
rect 20257 9027 20315 9033
rect 20257 9024 20269 9027
rect 20036 8996 20269 9024
rect 20036 8984 20042 8996
rect 20257 8993 20269 8996
rect 20303 8993 20315 9027
rect 20257 8987 20315 8993
rect 31021 9027 31079 9033
rect 31021 8993 31033 9027
rect 31067 8993 31079 9027
rect 31021 8987 31079 8993
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 3786 8956 3792 8968
rect 2731 8928 3792 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 4338 8916 4344 8968
rect 4396 8916 4402 8968
rect 30466 8916 30472 8968
rect 30524 8916 30530 8968
rect 31036 8956 31064 8987
rect 31662 8984 31668 9036
rect 31720 8984 31726 9036
rect 31294 8956 31300 8968
rect 31036 8928 31300 8956
rect 31294 8916 31300 8928
rect 31352 8916 31358 8968
rect 31570 8916 31576 8968
rect 31628 8916 31634 8968
rect 30484 8888 30512 8916
rect 31910 8891 31968 8897
rect 31910 8888 31922 8891
rect 30484 8860 31922 8888
rect 31910 8857 31922 8860
rect 31956 8857 31968 8891
rect 31910 8851 31968 8857
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3200 8792 3801 8820
rect 3200 8780 3206 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 31202 8780 31208 8832
rect 31260 8820 31266 8832
rect 33045 8823 33103 8829
rect 33045 8820 33057 8823
rect 31260 8792 33057 8820
rect 31260 8780 31266 8792
rect 33045 8789 33057 8792
rect 33091 8789 33103 8823
rect 33045 8783 33103 8789
rect 1104 8730 34016 8752
rect 1104 8678 9138 8730
rect 9190 8678 9202 8730
rect 9254 8678 9266 8730
rect 9318 8678 9330 8730
rect 9382 8678 9394 8730
rect 9446 8678 17326 8730
rect 17378 8678 17390 8730
rect 17442 8678 17454 8730
rect 17506 8678 17518 8730
rect 17570 8678 17582 8730
rect 17634 8678 25514 8730
rect 25566 8678 25578 8730
rect 25630 8678 25642 8730
rect 25694 8678 25706 8730
rect 25758 8678 25770 8730
rect 25822 8678 33702 8730
rect 33754 8678 33766 8730
rect 33818 8678 33830 8730
rect 33882 8678 33894 8730
rect 33946 8678 33958 8730
rect 34010 8678 34016 8730
rect 1104 8656 34016 8678
rect 3602 8616 3608 8628
rect 2047 8588 3608 8616
rect 2047 8557 2075 8588
rect 3602 8576 3608 8588
rect 3660 8576 3666 8628
rect 30561 8619 30619 8625
rect 30561 8585 30573 8619
rect 30607 8616 30619 8619
rect 31110 8616 31116 8628
rect 30607 8588 31116 8616
rect 30607 8585 30619 8588
rect 30561 8579 30619 8585
rect 31110 8576 31116 8588
rect 31168 8576 31174 8628
rect 2032 8551 2090 8557
rect 2032 8517 2044 8551
rect 2078 8517 2090 8551
rect 2032 8511 2090 8517
rect 31570 8508 31576 8560
rect 31628 8548 31634 8560
rect 32585 8551 32643 8557
rect 32585 8548 32597 8551
rect 31628 8520 32597 8548
rect 31628 8508 31634 8520
rect 32585 8517 32597 8520
rect 32631 8517 32643 8551
rect 32585 8511 32643 8517
rect 31941 8483 31999 8489
rect 31941 8449 31953 8483
rect 31987 8480 31999 8483
rect 32217 8483 32275 8489
rect 32217 8480 32229 8483
rect 31987 8452 32229 8480
rect 31987 8449 31999 8452
rect 31941 8443 31999 8449
rect 32217 8449 32229 8452
rect 32263 8449 32275 8483
rect 32217 8443 32275 8449
rect 1762 8372 1768 8424
rect 1820 8372 1826 8424
rect 3789 8415 3847 8421
rect 3789 8412 3801 8415
rect 3160 8384 3801 8412
rect 3160 8353 3188 8384
rect 3789 8381 3801 8384
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 4488 8384 4844 8412
rect 4488 8372 4494 8384
rect 3145 8347 3203 8353
rect 3145 8313 3157 8347
rect 3191 8313 3203 8347
rect 3145 8307 3203 8313
rect 3970 8304 3976 8356
rect 4028 8304 4034 8356
rect 4157 8347 4215 8353
rect 4157 8313 4169 8347
rect 4203 8344 4215 8347
rect 4338 8344 4344 8356
rect 4203 8316 4344 8344
rect 4203 8313 4215 8316
rect 4157 8307 4215 8313
rect 4338 8304 4344 8316
rect 4396 8304 4402 8356
rect 4816 8288 4844 8384
rect 30098 8372 30104 8424
rect 30156 8412 30162 8424
rect 30377 8415 30435 8421
rect 30377 8412 30389 8415
rect 30156 8384 30389 8412
rect 30156 8372 30162 8384
rect 30377 8381 30389 8384
rect 30423 8381 30435 8415
rect 30377 8375 30435 8381
rect 31202 8372 31208 8424
rect 31260 8372 31266 8424
rect 31294 8372 31300 8424
rect 31352 8372 31358 8424
rect 28994 8304 29000 8356
rect 29052 8344 29058 8356
rect 29825 8347 29883 8353
rect 29825 8344 29837 8347
rect 29052 8316 29837 8344
rect 29052 8304 29058 8316
rect 29825 8313 29837 8316
rect 29871 8313 29883 8347
rect 29825 8307 29883 8313
rect 3234 8236 3240 8288
rect 3292 8236 3298 8288
rect 4798 8236 4804 8288
rect 4856 8236 4862 8288
rect 29454 8236 29460 8288
rect 29512 8236 29518 8288
rect 1104 8186 33856 8208
rect 1104 8134 5044 8186
rect 5096 8134 5108 8186
rect 5160 8134 5172 8186
rect 5224 8134 5236 8186
rect 5288 8134 5300 8186
rect 5352 8134 13232 8186
rect 13284 8134 13296 8186
rect 13348 8134 13360 8186
rect 13412 8134 13424 8186
rect 13476 8134 13488 8186
rect 13540 8134 21420 8186
rect 21472 8134 21484 8186
rect 21536 8134 21548 8186
rect 21600 8134 21612 8186
rect 21664 8134 21676 8186
rect 21728 8134 29608 8186
rect 29660 8134 29672 8186
rect 29724 8134 29736 8186
rect 29788 8134 29800 8186
rect 29852 8134 29864 8186
rect 29916 8134 33856 8186
rect 1104 8112 33856 8134
rect 3513 8075 3571 8081
rect 3513 8041 3525 8075
rect 3559 8072 3571 8075
rect 4338 8072 4344 8084
rect 3559 8044 4344 8072
rect 3559 8041 3571 8044
rect 3513 8035 3571 8041
rect 4338 8032 4344 8044
rect 4396 8032 4402 8084
rect 29365 8075 29423 8081
rect 29365 8041 29377 8075
rect 29411 8072 29423 8075
rect 32030 8072 32036 8084
rect 29411 8044 32036 8072
rect 29411 8041 29423 8044
rect 29365 8035 29423 8041
rect 32030 8032 32036 8044
rect 32088 8032 32094 8084
rect 4706 7964 4712 8016
rect 4764 7964 4770 8016
rect 29273 8007 29331 8013
rect 29273 7973 29285 8007
rect 29319 7973 29331 8007
rect 29273 7967 29331 7973
rect 30009 8007 30067 8013
rect 30009 7973 30021 8007
rect 30055 8004 30067 8007
rect 30558 8004 30564 8016
rect 30055 7976 30564 8004
rect 30055 7973 30067 7976
rect 30009 7967 30067 7973
rect 1578 7896 1584 7948
rect 1636 7896 1642 7948
rect 2961 7939 3019 7945
rect 2961 7905 2973 7939
rect 3007 7936 3019 7939
rect 3234 7936 3240 7948
rect 3007 7908 3240 7936
rect 3007 7905 3019 7908
rect 2961 7899 3019 7905
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4525 7939 4583 7945
rect 4525 7936 4537 7939
rect 4212 7908 4537 7936
rect 4212 7896 4218 7908
rect 4525 7905 4537 7908
rect 4571 7905 4583 7939
rect 29288 7936 29316 7967
rect 30558 7964 30564 7976
rect 30616 8004 30622 8016
rect 31294 8004 31300 8016
rect 30616 7976 31300 8004
rect 30616 7964 30622 7976
rect 31294 7964 31300 7976
rect 31352 7964 31358 8016
rect 29822 7936 29828 7948
rect 29288 7908 29828 7936
rect 4525 7899 4583 7905
rect 29822 7896 29828 7908
rect 29880 7936 29886 7948
rect 30193 7939 30251 7945
rect 30193 7936 30205 7939
rect 29880 7908 30205 7936
rect 29880 7896 29886 7908
rect 30193 7905 30205 7908
rect 30239 7905 30251 7939
rect 30193 7899 30251 7905
rect 31662 7896 31668 7948
rect 31720 7896 31726 7948
rect 2590 7828 2596 7880
rect 2648 7828 2654 7880
rect 3786 7828 3792 7880
rect 3844 7828 3850 7880
rect 30837 7871 30895 7877
rect 30837 7837 30849 7871
rect 30883 7868 30895 7871
rect 30929 7871 30987 7877
rect 30929 7868 30941 7871
rect 30883 7840 30941 7868
rect 30883 7837 30895 7840
rect 30837 7831 30895 7837
rect 30929 7837 30941 7840
rect 30975 7837 30987 7871
rect 30929 7831 30987 7837
rect 31573 7871 31631 7877
rect 31573 7837 31585 7871
rect 31619 7868 31631 7871
rect 31619 7840 33088 7868
rect 31619 7837 31631 7840
rect 31573 7831 31631 7837
rect 4338 7760 4344 7812
rect 4396 7800 4402 7812
rect 4798 7800 4804 7812
rect 4396 7772 4804 7800
rect 4396 7760 4402 7772
rect 4798 7760 4804 7772
rect 4856 7800 4862 7812
rect 4985 7803 5043 7809
rect 4985 7800 4997 7803
rect 4856 7772 4997 7800
rect 4856 7760 4862 7772
rect 4985 7769 4997 7772
rect 5031 7800 5043 7803
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 5031 7772 5273 7800
rect 5031 7769 5043 7772
rect 4985 7763 5043 7769
rect 5261 7769 5273 7772
rect 5307 7769 5319 7803
rect 28905 7803 28963 7809
rect 28905 7800 28917 7803
rect 5261 7763 5319 7769
rect 28736 7772 28917 7800
rect 4430 7692 4436 7744
rect 4488 7692 4494 7744
rect 27246 7692 27252 7744
rect 27304 7732 27310 7744
rect 28736 7741 28764 7772
rect 28905 7769 28917 7772
rect 28951 7800 28963 7803
rect 29454 7800 29460 7812
rect 28951 7772 29460 7800
rect 28951 7769 28963 7772
rect 28905 7763 28963 7769
rect 29454 7760 29460 7772
rect 29512 7800 29518 7812
rect 29641 7803 29699 7809
rect 29641 7800 29653 7803
rect 29512 7772 29653 7800
rect 29512 7760 29518 7772
rect 29641 7769 29653 7772
rect 29687 7769 29699 7803
rect 31910 7803 31968 7809
rect 31910 7800 31922 7803
rect 29641 7763 29699 7769
rect 30116 7772 31922 7800
rect 30116 7741 30144 7772
rect 31910 7769 31922 7772
rect 31956 7769 31968 7803
rect 31910 7763 31968 7769
rect 33060 7741 33088 7840
rect 28721 7735 28779 7741
rect 28721 7732 28733 7735
rect 27304 7704 28733 7732
rect 27304 7692 27310 7704
rect 28721 7701 28733 7704
rect 28767 7701 28779 7735
rect 28721 7695 28779 7701
rect 30101 7735 30159 7741
rect 30101 7701 30113 7735
rect 30147 7701 30159 7735
rect 30101 7695 30159 7701
rect 33045 7735 33103 7741
rect 33045 7701 33057 7735
rect 33091 7701 33103 7735
rect 33045 7695 33103 7701
rect 1104 7642 34016 7664
rect 1104 7590 9138 7642
rect 9190 7590 9202 7642
rect 9254 7590 9266 7642
rect 9318 7590 9330 7642
rect 9382 7590 9394 7642
rect 9446 7590 17326 7642
rect 17378 7590 17390 7642
rect 17442 7590 17454 7642
rect 17506 7590 17518 7642
rect 17570 7590 17582 7642
rect 17634 7590 25514 7642
rect 25566 7590 25578 7642
rect 25630 7590 25642 7642
rect 25694 7590 25706 7642
rect 25758 7590 25770 7642
rect 25822 7590 33702 7642
rect 33754 7590 33766 7642
rect 33818 7590 33830 7642
rect 33882 7590 33894 7642
rect 33946 7590 33958 7642
rect 34010 7590 34016 7642
rect 1104 7568 34016 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 1820 7500 4200 7528
rect 1820 7488 1826 7500
rect 2317 7463 2375 7469
rect 2317 7429 2329 7463
rect 2363 7460 2375 7463
rect 2590 7460 2596 7472
rect 2363 7432 2596 7460
rect 2363 7429 2375 7432
rect 2317 7423 2375 7429
rect 2590 7420 2596 7432
rect 2648 7420 2654 7472
rect 2685 7395 2743 7401
rect 2685 7361 2697 7395
rect 2731 7392 2743 7395
rect 3142 7392 3148 7404
rect 2731 7364 3148 7392
rect 2731 7361 2743 7364
rect 2685 7355 2743 7361
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3602 7352 3608 7404
rect 3660 7392 3666 7404
rect 3982 7395 4040 7401
rect 3982 7392 3994 7395
rect 3660 7364 3994 7392
rect 3660 7352 3666 7364
rect 3982 7361 3994 7364
rect 4028 7361 4040 7395
rect 4172 7392 4200 7500
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 4448 7401 4476 7488
rect 30469 7463 30527 7469
rect 30469 7429 30481 7463
rect 30515 7460 30527 7463
rect 30515 7432 31754 7460
rect 30515 7429 30527 7432
rect 30469 7423 30527 7429
rect 4249 7395 4307 7401
rect 4249 7392 4261 7395
rect 4172 7364 4261 7392
rect 3982 7355 4040 7361
rect 4249 7361 4261 7364
rect 4295 7361 4307 7395
rect 4249 7355 4307 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17313 7395 17371 7401
rect 17313 7392 17325 7395
rect 17000 7364 17325 7392
rect 17000 7352 17006 7364
rect 17313 7361 17325 7364
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 28994 7352 29000 7404
rect 29052 7352 29058 7404
rect 29822 7352 29828 7404
rect 29880 7352 29886 7404
rect 30745 7395 30803 7401
rect 30745 7361 30757 7395
rect 30791 7392 30803 7395
rect 31018 7392 31024 7404
rect 30791 7364 31024 7392
rect 30791 7361 30803 7364
rect 30745 7355 30803 7361
rect 31018 7352 31024 7364
rect 31076 7352 31082 7404
rect 31726 7392 31754 7432
rect 32217 7395 32275 7401
rect 32217 7392 32229 7395
rect 31726 7364 32229 7392
rect 32217 7361 32229 7364
rect 32263 7361 32275 7395
rect 32217 7355 32275 7361
rect 27338 7284 27344 7336
rect 27396 7324 27402 7336
rect 29641 7327 29699 7333
rect 29641 7324 29653 7327
rect 27396 7296 29653 7324
rect 27396 7284 27402 7296
rect 29641 7293 29653 7296
rect 29687 7293 29699 7327
rect 29641 7287 29699 7293
rect 31202 7284 31208 7336
rect 31260 7284 31266 7336
rect 32490 7284 32496 7336
rect 32548 7284 32554 7336
rect 2866 7148 2872 7200
rect 2924 7148 2930 7200
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 4706 7188 4712 7200
rect 4488 7160 4712 7188
rect 4488 7148 4494 7160
rect 4706 7148 4712 7160
rect 4764 7188 4770 7200
rect 4985 7191 5043 7197
rect 4985 7188 4997 7191
rect 4764 7160 4997 7188
rect 4764 7148 4770 7160
rect 4985 7157 4997 7160
rect 5031 7157 5043 7191
rect 4985 7151 5043 7157
rect 16758 7148 16764 7200
rect 16816 7148 16822 7200
rect 27522 7148 27528 7200
rect 27580 7188 27586 7200
rect 27985 7191 28043 7197
rect 27985 7188 27997 7191
rect 27580 7160 27997 7188
rect 27580 7148 27586 7160
rect 27985 7157 27997 7160
rect 28031 7157 28043 7191
rect 27985 7151 28043 7157
rect 28350 7148 28356 7200
rect 28408 7148 28414 7200
rect 29086 7148 29092 7200
rect 29144 7148 29150 7200
rect 1104 7098 33856 7120
rect 1104 7046 5044 7098
rect 5096 7046 5108 7098
rect 5160 7046 5172 7098
rect 5224 7046 5236 7098
rect 5288 7046 5300 7098
rect 5352 7046 13232 7098
rect 13284 7046 13296 7098
rect 13348 7046 13360 7098
rect 13412 7046 13424 7098
rect 13476 7046 13488 7098
rect 13540 7046 21420 7098
rect 21472 7046 21484 7098
rect 21536 7046 21548 7098
rect 21600 7046 21612 7098
rect 21664 7046 21676 7098
rect 21728 7046 29608 7098
rect 29660 7046 29672 7098
rect 29724 7046 29736 7098
rect 29788 7046 29800 7098
rect 29852 7046 29864 7098
rect 29916 7046 33856 7098
rect 1104 7024 33856 7046
rect 3145 6987 3203 6993
rect 3145 6953 3157 6987
rect 3191 6984 3203 6987
rect 3786 6984 3792 6996
rect 3191 6956 3792 6984
rect 3191 6953 3203 6956
rect 3145 6947 3203 6953
rect 3786 6944 3792 6956
rect 3844 6944 3850 6996
rect 26234 6876 26240 6928
rect 26292 6916 26298 6928
rect 28721 6919 28779 6925
rect 28721 6916 28733 6919
rect 26292 6888 28733 6916
rect 26292 6876 26298 6888
rect 28721 6885 28733 6888
rect 28767 6885 28779 6919
rect 28721 6879 28779 6885
rect 1762 6808 1768 6860
rect 1820 6808 1826 6860
rect 4430 6808 4436 6860
rect 4488 6808 4494 6860
rect 28074 6808 28080 6860
rect 28132 6848 28138 6860
rect 29086 6848 29092 6860
rect 28132 6820 29092 6848
rect 28132 6808 28138 6820
rect 29086 6808 29092 6820
rect 29144 6808 29150 6860
rect 33318 6808 33324 6860
rect 33376 6808 33382 6860
rect 2032 6783 2090 6789
rect 2032 6749 2044 6783
rect 2078 6780 2090 6783
rect 3970 6780 3976 6792
rect 2078 6752 3976 6780
rect 2078 6749 2090 6752
rect 2032 6743 2090 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4522 6740 4528 6792
rect 4580 6780 4586 6792
rect 5077 6783 5135 6789
rect 5077 6780 5089 6783
rect 4580 6752 5089 6780
rect 4580 6740 4586 6752
rect 5077 6749 5089 6752
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 28629 6783 28687 6789
rect 28629 6749 28641 6783
rect 28675 6780 28687 6783
rect 29178 6780 29184 6792
rect 28675 6752 29184 6780
rect 28675 6749 28687 6752
rect 28629 6743 28687 6749
rect 29178 6740 29184 6752
rect 29236 6740 29242 6792
rect 29365 6783 29423 6789
rect 29365 6749 29377 6783
rect 29411 6749 29423 6783
rect 29365 6743 29423 6749
rect 27522 6672 27528 6724
rect 27580 6672 27586 6724
rect 29380 6712 29408 6743
rect 30558 6740 30564 6792
rect 30616 6740 30622 6792
rect 30742 6740 30748 6792
rect 30800 6740 30806 6792
rect 31018 6740 31024 6792
rect 31076 6780 31082 6792
rect 31113 6783 31171 6789
rect 31113 6780 31125 6783
rect 31076 6752 31125 6780
rect 31076 6740 31082 6752
rect 31113 6749 31125 6752
rect 31159 6749 31171 6783
rect 31113 6743 31171 6749
rect 32309 6783 32367 6789
rect 32309 6749 32321 6783
rect 32355 6780 32367 6783
rect 32490 6780 32496 6792
rect 32355 6752 32496 6780
rect 32355 6749 32367 6752
rect 32309 6743 32367 6749
rect 32490 6740 32496 6752
rect 32548 6740 32554 6792
rect 32582 6712 32588 6724
rect 29380 6684 32588 6712
rect 32582 6672 32588 6684
rect 32640 6672 32646 6724
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 3789 6647 3847 6653
rect 3789 6644 3801 6647
rect 2832 6616 3801 6644
rect 2832 6604 2838 6616
rect 3789 6613 3801 6616
rect 3835 6613 3847 6647
rect 3789 6607 3847 6613
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4525 6647 4583 6653
rect 4525 6644 4537 6647
rect 4304 6616 4537 6644
rect 4304 6604 4310 6616
rect 4525 6613 4537 6616
rect 4571 6613 4583 6647
rect 4525 6607 4583 6613
rect 27614 6604 27620 6656
rect 27672 6604 27678 6656
rect 29917 6647 29975 6653
rect 29917 6613 29929 6647
rect 29963 6644 29975 6647
rect 30466 6644 30472 6656
rect 29963 6616 30472 6644
rect 29963 6613 29975 6616
rect 29917 6607 29975 6613
rect 30466 6604 30472 6616
rect 30524 6604 30530 6656
rect 1104 6554 34016 6576
rect 1104 6502 9138 6554
rect 9190 6502 9202 6554
rect 9254 6502 9266 6554
rect 9318 6502 9330 6554
rect 9382 6502 9394 6554
rect 9446 6502 17326 6554
rect 17378 6502 17390 6554
rect 17442 6502 17454 6554
rect 17506 6502 17518 6554
rect 17570 6502 17582 6554
rect 17634 6502 25514 6554
rect 25566 6502 25578 6554
rect 25630 6502 25642 6554
rect 25694 6502 25706 6554
rect 25758 6502 25770 6554
rect 25822 6502 33702 6554
rect 33754 6502 33766 6554
rect 33818 6502 33830 6554
rect 33882 6502 33894 6554
rect 33946 6502 33958 6554
rect 34010 6502 34016 6554
rect 1104 6480 34016 6502
rect 4706 6400 4712 6452
rect 4764 6400 4770 6452
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 27246 6440 27252 6452
rect 25280 6412 27252 6440
rect 25280 6400 25286 6412
rect 27246 6400 27252 6412
rect 27304 6400 27310 6452
rect 28997 6443 29055 6449
rect 28997 6409 29009 6443
rect 29043 6440 29055 6443
rect 30742 6440 30748 6452
rect 29043 6412 30748 6440
rect 29043 6409 29055 6412
rect 28997 6403 29055 6409
rect 30742 6400 30748 6412
rect 30800 6400 30806 6452
rect 33505 6443 33563 6449
rect 33505 6440 33517 6443
rect 31726 6412 33517 6440
rect 2032 6375 2090 6381
rect 2032 6341 2044 6375
rect 2078 6372 2090 6375
rect 4154 6372 4160 6384
rect 2078 6344 4160 6372
rect 2078 6341 2090 6344
rect 2032 6335 2090 6341
rect 4154 6332 4160 6344
rect 4212 6332 4218 6384
rect 26789 6375 26847 6381
rect 26789 6341 26801 6375
rect 26835 6372 26847 6375
rect 27157 6375 27215 6381
rect 27157 6372 27169 6375
rect 26835 6344 27169 6372
rect 26835 6341 26847 6344
rect 26789 6335 26847 6341
rect 27157 6341 27169 6344
rect 27203 6372 27215 6375
rect 27614 6372 27620 6384
rect 27203 6344 27620 6372
rect 27203 6341 27215 6344
rect 27157 6335 27215 6341
rect 27614 6332 27620 6344
rect 27672 6332 27678 6384
rect 30558 6332 30564 6384
rect 30616 6372 30622 6384
rect 31726 6372 31754 6412
rect 33505 6409 33517 6412
rect 33551 6409 33563 6443
rect 33505 6403 33563 6409
rect 30616 6344 31754 6372
rect 30616 6332 30622 6344
rect 32030 6332 32036 6384
rect 32088 6372 32094 6384
rect 32370 6375 32428 6381
rect 32370 6372 32382 6375
rect 32088 6344 32382 6372
rect 32088 6332 32094 6344
rect 32370 6341 32382 6344
rect 32416 6341 32428 6375
rect 32370 6335 32428 6341
rect 1762 6264 1768 6316
rect 1820 6264 1826 6316
rect 3234 6264 3240 6316
rect 3292 6264 3298 6316
rect 30469 6307 30527 6313
rect 30469 6273 30481 6307
rect 30515 6304 30527 6307
rect 30926 6304 30932 6316
rect 30515 6276 30932 6304
rect 30515 6273 30527 6276
rect 30469 6267 30527 6273
rect 30926 6264 30932 6276
rect 30984 6264 30990 6316
rect 31662 6264 31668 6316
rect 31720 6264 31726 6316
rect 31938 6264 31944 6316
rect 31996 6264 32002 6316
rect 3697 6239 3755 6245
rect 3697 6205 3709 6239
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3712 6168 3740 6199
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 4396 6208 5273 6236
rect 4396 6196 4402 6208
rect 5261 6205 5273 6208
rect 5307 6205 5319 6239
rect 5261 6199 5319 6205
rect 9585 6239 9643 6245
rect 9585 6205 9597 6239
rect 9631 6236 9643 6239
rect 9631 6208 10456 6236
rect 9631 6205 9643 6208
rect 9585 6199 9643 6205
rect 2700 6140 3740 6168
rect 1302 6060 1308 6112
rect 1360 6100 1366 6112
rect 2700 6100 2728 6140
rect 9858 6128 9864 6180
rect 9916 6128 9922 6180
rect 10428 6112 10456 6208
rect 27614 6196 27620 6248
rect 27672 6196 27678 6248
rect 28445 6239 28503 6245
rect 28445 6205 28457 6239
rect 28491 6236 28503 6239
rect 28810 6236 28816 6248
rect 28491 6208 28816 6236
rect 28491 6205 28503 6208
rect 28445 6199 28503 6205
rect 28810 6196 28816 6208
rect 28868 6196 28874 6248
rect 30009 6239 30067 6245
rect 30009 6205 30021 6239
rect 30055 6205 30067 6239
rect 30009 6199 30067 6205
rect 1360 6072 2728 6100
rect 1360 6060 1366 6072
rect 3142 6060 3148 6112
rect 3200 6060 3206 6112
rect 10045 6103 10103 6109
rect 10045 6069 10057 6103
rect 10091 6100 10103 6103
rect 10226 6100 10232 6112
rect 10091 6072 10232 6100
rect 10091 6069 10103 6072
rect 10045 6063 10103 6069
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10410 6060 10416 6112
rect 10468 6060 10474 6112
rect 28261 6103 28319 6109
rect 28261 6069 28273 6103
rect 28307 6100 28319 6103
rect 29086 6100 29092 6112
rect 28307 6072 29092 6100
rect 28307 6069 28319 6072
rect 28261 6063 28319 6069
rect 29086 6060 29092 6072
rect 29144 6060 29150 6112
rect 30024 6100 30052 6199
rect 31478 6196 31484 6248
rect 31536 6196 31542 6248
rect 31680 6236 31708 6264
rect 32122 6236 32128 6248
rect 31680 6208 32128 6236
rect 32122 6196 32128 6208
rect 32180 6196 32186 6248
rect 34054 6100 34060 6112
rect 30024 6072 34060 6100
rect 34054 6060 34060 6072
rect 34112 6060 34118 6112
rect 1104 6010 33856 6032
rect 1104 5958 5044 6010
rect 5096 5958 5108 6010
rect 5160 5958 5172 6010
rect 5224 5958 5236 6010
rect 5288 5958 5300 6010
rect 5352 5958 13232 6010
rect 13284 5958 13296 6010
rect 13348 5958 13360 6010
rect 13412 5958 13424 6010
rect 13476 5958 13488 6010
rect 13540 5958 21420 6010
rect 21472 5958 21484 6010
rect 21536 5958 21548 6010
rect 21600 5958 21612 6010
rect 21664 5958 21676 6010
rect 21728 5958 29608 6010
rect 29660 5958 29672 6010
rect 29724 5958 29736 6010
rect 29788 5958 29800 6010
rect 29852 5958 29864 6010
rect 29916 5958 33856 6010
rect 1104 5936 33856 5958
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 4338 5896 4344 5908
rect 3559 5868 4344 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 4522 5896 4528 5908
rect 4479 5868 4528 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 10413 5899 10471 5905
rect 10413 5865 10425 5899
rect 10459 5896 10471 5899
rect 15194 5896 15200 5908
rect 10459 5868 15200 5896
rect 10459 5865 10471 5868
rect 10413 5859 10471 5865
rect 15194 5856 15200 5868
rect 15252 5856 15258 5908
rect 24949 5899 25007 5905
rect 24949 5865 24961 5899
rect 24995 5896 25007 5899
rect 26142 5896 26148 5908
rect 24995 5868 26148 5896
rect 24995 5865 25007 5868
rect 24949 5859 25007 5865
rect 26142 5856 26148 5868
rect 26200 5896 26206 5908
rect 26510 5896 26516 5908
rect 26200 5868 26516 5896
rect 26200 5856 26206 5868
rect 26510 5856 26516 5868
rect 26568 5856 26574 5908
rect 27338 5856 27344 5908
rect 27396 5856 27402 5908
rect 27433 5899 27491 5905
rect 27433 5865 27445 5899
rect 27479 5896 27491 5899
rect 27614 5896 27620 5908
rect 27479 5868 27620 5896
rect 27479 5865 27491 5868
rect 27433 5859 27491 5865
rect 27614 5856 27620 5868
rect 27672 5856 27678 5908
rect 31754 5896 31760 5908
rect 29012 5868 31760 5896
rect 11698 5788 11704 5840
rect 11756 5788 11762 5840
rect 25222 5788 25228 5840
rect 25280 5828 25286 5840
rect 25777 5831 25835 5837
rect 25777 5828 25789 5831
rect 25280 5800 25789 5828
rect 25280 5788 25286 5800
rect 25777 5797 25789 5800
rect 25823 5797 25835 5831
rect 25777 5791 25835 5797
rect 26605 5831 26663 5837
rect 26605 5797 26617 5831
rect 26651 5828 26663 5831
rect 29012 5828 29040 5868
rect 31754 5856 31760 5868
rect 31812 5856 31818 5908
rect 26651 5800 29040 5828
rect 26651 5797 26663 5800
rect 26605 5791 26663 5797
rect 29086 5788 29092 5840
rect 29144 5828 29150 5840
rect 30374 5828 30380 5840
rect 29144 5800 30380 5828
rect 29144 5788 29150 5800
rect 30374 5788 30380 5800
rect 30432 5788 30438 5840
rect 1578 5720 1584 5772
rect 1636 5720 1642 5772
rect 2866 5720 2872 5772
rect 2924 5720 2930 5772
rect 8846 5720 8852 5772
rect 8904 5760 8910 5772
rect 11517 5763 11575 5769
rect 11517 5760 11529 5763
rect 8904 5732 11529 5760
rect 8904 5720 8910 5732
rect 11517 5729 11529 5732
rect 11563 5729 11575 5763
rect 11517 5723 11575 5729
rect 26053 5763 26111 5769
rect 26053 5729 26065 5763
rect 26099 5760 26111 5763
rect 26786 5760 26792 5772
rect 26099 5732 26792 5760
rect 26099 5729 26111 5732
rect 26053 5723 26111 5729
rect 26786 5720 26792 5732
rect 26844 5760 26850 5772
rect 28350 5760 28356 5772
rect 26844 5732 28356 5760
rect 26844 5720 26850 5732
rect 28350 5720 28356 5732
rect 28408 5720 28414 5772
rect 29365 5763 29423 5769
rect 29365 5729 29377 5763
rect 29411 5760 29423 5763
rect 29454 5760 29460 5772
rect 29411 5732 29460 5760
rect 29411 5729 29423 5732
rect 29365 5723 29423 5729
rect 29454 5720 29460 5732
rect 29512 5760 29518 5772
rect 29733 5763 29791 5769
rect 29733 5760 29745 5763
rect 29512 5732 29745 5760
rect 29512 5720 29518 5732
rect 29733 5729 29745 5732
rect 29779 5729 29791 5763
rect 29733 5723 29791 5729
rect 30466 5720 30472 5772
rect 30524 5720 30530 5772
rect 31573 5763 31631 5769
rect 31573 5729 31585 5763
rect 31619 5729 31631 5763
rect 31573 5723 31631 5729
rect 2590 5652 2596 5704
rect 2648 5652 2654 5704
rect 3510 5652 3516 5704
rect 3568 5692 3574 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3568 5664 3801 5692
rect 3568 5652 3574 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 10042 5652 10048 5704
rect 10100 5652 10106 5704
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5692 10287 5695
rect 10686 5692 10692 5704
rect 10275 5664 10692 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 26694 5652 26700 5704
rect 26752 5652 26758 5704
rect 28077 5695 28135 5701
rect 28077 5661 28089 5695
rect 28123 5661 28135 5695
rect 28077 5655 28135 5661
rect 8754 5584 8760 5636
rect 8812 5624 8818 5636
rect 10410 5624 10416 5636
rect 8812 5596 10416 5624
rect 8812 5584 8818 5596
rect 10410 5584 10416 5596
rect 10468 5624 10474 5636
rect 11977 5627 12035 5633
rect 11977 5624 11989 5627
rect 10468 5596 11989 5624
rect 10468 5584 10474 5596
rect 11977 5593 11989 5596
rect 12023 5593 12035 5627
rect 28092 5624 28120 5655
rect 28166 5652 28172 5704
rect 28224 5652 28230 5704
rect 28813 5695 28871 5701
rect 28813 5661 28825 5695
rect 28859 5692 28871 5695
rect 31110 5692 31116 5704
rect 28859 5664 31116 5692
rect 28859 5661 28871 5664
rect 28813 5655 28871 5661
rect 31110 5652 31116 5664
rect 31168 5652 31174 5704
rect 31588 5636 31616 5723
rect 31938 5720 31944 5772
rect 31996 5760 32002 5772
rect 33137 5763 33195 5769
rect 33137 5760 33149 5763
rect 31996 5732 33149 5760
rect 31996 5720 32002 5732
rect 33137 5729 33149 5732
rect 33183 5729 33195 5763
rect 33137 5723 33195 5729
rect 32030 5652 32036 5704
rect 32088 5652 32094 5704
rect 32858 5652 32864 5704
rect 32916 5652 32922 5704
rect 29270 5624 29276 5636
rect 28092 5596 29276 5624
rect 11977 5587 12035 5593
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9493 5559 9551 5565
rect 9493 5556 9505 5559
rect 9088 5528 9505 5556
rect 9088 5516 9094 5528
rect 9493 5525 9505 5528
rect 9539 5525 9551 5559
rect 11992 5556 12020 5587
rect 29270 5584 29276 5596
rect 29328 5584 29334 5636
rect 31570 5584 31576 5636
rect 31628 5584 31634 5636
rect 12345 5559 12403 5565
rect 12345 5556 12357 5559
rect 11992 5528 12357 5556
rect 9493 5519 9551 5525
rect 12345 5525 12357 5528
rect 12391 5556 12403 5559
rect 12526 5556 12532 5568
rect 12391 5528 12532 5556
rect 12391 5525 12403 5528
rect 12345 5519 12403 5525
rect 12526 5516 12532 5528
rect 12584 5556 12590 5568
rect 13722 5556 13728 5568
rect 12584 5528 13728 5556
rect 12584 5516 12590 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 28902 5516 28908 5568
rect 28960 5516 28966 5568
rect 29914 5516 29920 5568
rect 29972 5516 29978 5568
rect 1104 5466 34016 5488
rect 1104 5414 9138 5466
rect 9190 5414 9202 5466
rect 9254 5414 9266 5466
rect 9318 5414 9330 5466
rect 9382 5414 9394 5466
rect 9446 5414 17326 5466
rect 17378 5414 17390 5466
rect 17442 5414 17454 5466
rect 17506 5414 17518 5466
rect 17570 5414 17582 5466
rect 17634 5414 25514 5466
rect 25566 5414 25578 5466
rect 25630 5414 25642 5466
rect 25694 5414 25706 5466
rect 25758 5414 25770 5466
rect 25822 5414 33702 5466
rect 33754 5414 33766 5466
rect 33818 5414 33830 5466
rect 33882 5414 33894 5466
rect 33946 5414 33958 5466
rect 34010 5414 34016 5466
rect 1104 5392 34016 5414
rect 3510 5312 3516 5364
rect 3568 5312 3574 5364
rect 3602 5312 3608 5364
rect 3660 5312 3666 5364
rect 10042 5312 10048 5364
rect 10100 5312 10106 5364
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 12342 5352 12348 5364
rect 11756 5324 12348 5352
rect 11756 5312 11762 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 26050 5312 26056 5364
rect 26108 5312 26114 5364
rect 30098 5312 30104 5364
rect 30156 5312 30162 5364
rect 33502 5312 33508 5364
rect 33560 5312 33566 5364
rect 2317 5287 2375 5293
rect 2317 5253 2329 5287
rect 2363 5284 2375 5287
rect 2590 5284 2596 5296
rect 2363 5256 2596 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 2590 5244 2596 5256
rect 2648 5244 2654 5296
rect 8113 5287 8171 5293
rect 8113 5253 8125 5287
rect 8159 5284 8171 5287
rect 8386 5284 8392 5296
rect 8159 5256 8392 5284
rect 8159 5253 8171 5256
rect 8113 5247 8171 5253
rect 8386 5244 8392 5256
rect 8444 5284 8450 5296
rect 8754 5284 8760 5296
rect 8444 5256 8760 5284
rect 8444 5244 8450 5256
rect 8754 5244 8760 5256
rect 8812 5244 8818 5296
rect 13541 5287 13599 5293
rect 13541 5253 13553 5287
rect 13587 5284 13599 5287
rect 13630 5284 13636 5296
rect 13587 5256 13636 5284
rect 13587 5253 13599 5256
rect 13541 5247 13599 5253
rect 13630 5244 13636 5256
rect 13688 5284 13694 5296
rect 14185 5287 14243 5293
rect 14185 5284 14197 5287
rect 13688 5256 14197 5284
rect 13688 5244 13694 5256
rect 14185 5253 14197 5256
rect 14231 5284 14243 5287
rect 15197 5287 15255 5293
rect 15197 5284 15209 5287
rect 14231 5256 15209 5284
rect 14231 5253 14243 5256
rect 14185 5247 14243 5253
rect 15197 5253 15209 5256
rect 15243 5284 15255 5287
rect 15930 5284 15936 5296
rect 15243 5256 15936 5284
rect 15243 5253 15255 5256
rect 15197 5247 15255 5253
rect 15930 5244 15936 5256
rect 15988 5284 15994 5296
rect 16301 5287 16359 5293
rect 16301 5284 16313 5287
rect 15988 5256 16313 5284
rect 15988 5244 15994 5256
rect 16301 5253 16313 5256
rect 16347 5253 16359 5287
rect 16301 5247 16359 5253
rect 23382 5244 23388 5296
rect 23440 5284 23446 5296
rect 25222 5284 25228 5296
rect 23440 5256 25228 5284
rect 23440 5244 23446 5256
rect 25222 5244 25228 5256
rect 25280 5284 25286 5296
rect 25593 5287 25651 5293
rect 25593 5284 25605 5287
rect 25280 5256 25605 5284
rect 25280 5244 25286 5256
rect 25593 5253 25605 5256
rect 25639 5284 25651 5287
rect 27062 5284 27068 5296
rect 25639 5256 27068 5284
rect 25639 5253 25651 5256
rect 25593 5247 25651 5253
rect 27062 5244 27068 5256
rect 27120 5244 27126 5296
rect 29086 5244 29092 5296
rect 29144 5244 29150 5296
rect 29178 5244 29184 5296
rect 29236 5284 29242 5296
rect 32370 5287 32428 5293
rect 32370 5284 32382 5287
rect 29236 5256 32382 5284
rect 29236 5244 29242 5256
rect 32370 5253 32382 5256
rect 32416 5253 32428 5287
rect 32370 5247 32428 5253
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 2774 5216 2780 5228
rect 2731 5188 2780 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 2774 5176 2780 5188
rect 2832 5176 2838 5228
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 3142 5216 3148 5228
rect 3007 5188 3148 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4430 5216 4436 5228
rect 4111 5188 4436 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 9766 5216 9772 5228
rect 8220 5188 9772 5216
rect 3789 5083 3847 5089
rect 3789 5049 3801 5083
rect 3835 5080 3847 5083
rect 4522 5080 4528 5092
rect 3835 5052 4528 5080
rect 3835 5049 3847 5052
rect 3789 5043 3847 5049
rect 4522 5040 4528 5052
rect 4580 5040 4586 5092
rect 8220 5080 8248 5188
rect 9766 5176 9772 5188
rect 9824 5216 9830 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 9824 5188 11529 5216
rect 9824 5176 9830 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 13909 5219 13967 5225
rect 13909 5216 13921 5219
rect 13780 5188 13921 5216
rect 13780 5176 13786 5188
rect 13909 5185 13921 5188
rect 13955 5216 13967 5219
rect 14553 5219 14611 5225
rect 14553 5216 14565 5219
rect 13955 5188 14565 5216
rect 13955 5185 13967 5188
rect 13909 5179 13967 5185
rect 14553 5185 14565 5188
rect 14599 5185 14611 5219
rect 14553 5179 14611 5185
rect 16758 5176 16764 5228
rect 16816 5176 16822 5228
rect 24302 5176 24308 5228
rect 24360 5216 24366 5228
rect 24765 5219 24823 5225
rect 24765 5216 24777 5219
rect 24360 5188 24777 5216
rect 24360 5176 24366 5188
rect 24765 5185 24777 5188
rect 24811 5185 24823 5219
rect 24765 5179 24823 5185
rect 26234 5176 26240 5228
rect 26292 5176 26298 5228
rect 26789 5219 26847 5225
rect 26789 5185 26801 5219
rect 26835 5216 26847 5219
rect 28810 5216 28816 5228
rect 26835 5188 28816 5216
rect 26835 5185 26847 5188
rect 26789 5179 26847 5185
rect 28810 5176 28816 5188
rect 28868 5176 28874 5228
rect 28977 5219 29035 5225
rect 28977 5185 28989 5219
rect 29023 5216 29035 5219
rect 29104 5216 29132 5244
rect 29023 5188 29132 5216
rect 31573 5219 31631 5225
rect 29023 5185 29035 5188
rect 28977 5179 29035 5185
rect 31573 5185 31585 5219
rect 31619 5216 31631 5219
rect 31938 5216 31944 5228
rect 31619 5188 31944 5216
rect 31619 5185 31631 5188
rect 31573 5179 31631 5185
rect 31938 5176 31944 5188
rect 31996 5176 32002 5228
rect 32122 5176 32128 5228
rect 32180 5176 32186 5228
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 9030 5148 9036 5160
rect 8352 5120 9036 5148
rect 8352 5108 8358 5120
rect 9030 5108 9036 5120
rect 9088 5148 9094 5160
rect 9217 5151 9275 5157
rect 9217 5148 9229 5151
rect 9088 5120 9229 5148
rect 9088 5108 9094 5120
rect 9217 5117 9229 5120
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 10502 5148 10508 5160
rect 9539 5120 10508 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 10778 5108 10784 5160
rect 10836 5108 10842 5160
rect 12066 5108 12072 5160
rect 12124 5108 12130 5160
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12492 5120 12909 5148
rect 12492 5108 12498 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5148 15715 5151
rect 16574 5148 16580 5160
rect 15703 5120 16580 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 16574 5108 16580 5120
rect 16632 5108 16638 5160
rect 8389 5083 8447 5089
rect 8389 5080 8401 5083
rect 8220 5052 8401 5080
rect 8389 5049 8401 5052
rect 8435 5049 8447 5083
rect 8389 5043 8447 5049
rect 8478 5040 8484 5092
rect 8536 5080 8542 5092
rect 10229 5083 10287 5089
rect 10229 5080 10241 5083
rect 8536 5052 10241 5080
rect 8536 5040 8542 5052
rect 10229 5049 10241 5052
rect 10275 5049 10287 5083
rect 10229 5043 10287 5049
rect 15565 5083 15623 5089
rect 15565 5049 15577 5083
rect 15611 5080 15623 5083
rect 16776 5080 16804 5176
rect 24578 5108 24584 5160
rect 24636 5108 24642 5160
rect 26970 5108 26976 5160
rect 27028 5108 27034 5160
rect 27617 5151 27675 5157
rect 27617 5117 27629 5151
rect 27663 5148 27675 5151
rect 28261 5151 28319 5157
rect 28261 5148 28273 5151
rect 27663 5120 28273 5148
rect 27663 5117 27675 5120
rect 27617 5111 27675 5117
rect 28261 5117 28273 5120
rect 28307 5117 28319 5151
rect 28261 5111 28319 5117
rect 28718 5108 28724 5160
rect 28776 5108 28782 5160
rect 30098 5108 30104 5160
rect 30156 5148 30162 5160
rect 30377 5151 30435 5157
rect 30377 5148 30389 5151
rect 30156 5120 30389 5148
rect 30156 5108 30162 5120
rect 30377 5117 30389 5120
rect 30423 5117 30435 5151
rect 30377 5111 30435 5117
rect 15611 5052 16804 5080
rect 25961 5083 26019 5089
rect 15611 5049 15623 5052
rect 15565 5043 15623 5049
rect 25961 5049 25973 5083
rect 26007 5080 26019 5083
rect 26007 5052 28764 5080
rect 26007 5049 26019 5052
rect 25961 5043 26019 5049
rect 4430 4972 4436 5024
rect 4488 4972 4494 5024
rect 8570 4972 8576 5024
rect 8628 4972 8634 5024
rect 8662 4972 8668 5024
rect 8720 4972 8726 5024
rect 8754 4972 8760 5024
rect 8812 5012 8818 5024
rect 9858 5012 9864 5024
rect 8812 4984 9864 5012
rect 8812 4972 8818 4984
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 17313 5015 17371 5021
rect 17313 4981 17325 5015
rect 17359 5012 17371 5015
rect 19334 5012 19340 5024
rect 17359 4984 19340 5012
rect 17359 4981 17371 4984
rect 17313 4975 17371 4981
rect 19334 4972 19340 4984
rect 19392 4972 19398 5024
rect 24026 4972 24032 5024
rect 24084 4972 24090 5024
rect 25409 5015 25467 5021
rect 25409 4981 25421 5015
rect 25455 5012 25467 5015
rect 26602 5012 26608 5024
rect 25455 4984 26608 5012
rect 25455 4981 25467 4984
rect 25409 4975 25467 4981
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 27706 4972 27712 5024
rect 27764 4972 27770 5024
rect 28736 5012 28764 5052
rect 30006 5040 30012 5092
rect 30064 5040 30070 5092
rect 30024 5012 30052 5040
rect 28736 4984 30052 5012
rect 1104 4922 33856 4944
rect 1104 4870 5044 4922
rect 5096 4870 5108 4922
rect 5160 4870 5172 4922
rect 5224 4870 5236 4922
rect 5288 4870 5300 4922
rect 5352 4870 13232 4922
rect 13284 4870 13296 4922
rect 13348 4870 13360 4922
rect 13412 4870 13424 4922
rect 13476 4870 13488 4922
rect 13540 4870 21420 4922
rect 21472 4870 21484 4922
rect 21536 4870 21548 4922
rect 21600 4870 21612 4922
rect 21664 4870 21676 4922
rect 21728 4870 29608 4922
rect 29660 4870 29672 4922
rect 29724 4870 29736 4922
rect 29788 4870 29800 4922
rect 29852 4870 29864 4922
rect 29916 4870 33856 4922
rect 1104 4848 33856 4870
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 4488 4780 6914 4808
rect 4488 4768 4494 4780
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4672 2467 4675
rect 3234 4672 3240 4684
rect 2455 4644 3240 4672
rect 2455 4641 2467 4644
rect 2409 4635 2467 4641
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 4246 4604 4252 4616
rect 2731 4576 4252 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 6886 4604 6914 4780
rect 8478 4768 8484 4820
rect 8536 4768 8542 4820
rect 8570 4768 8576 4820
rect 8628 4768 8634 4820
rect 8754 4768 8760 4820
rect 8812 4768 8818 4820
rect 9490 4808 9496 4820
rect 9140 4780 9496 4808
rect 7929 4743 7987 4749
rect 7929 4709 7941 4743
rect 7975 4740 7987 4743
rect 8294 4740 8300 4752
rect 7975 4712 8300 4740
rect 7975 4709 7987 4712
rect 7929 4703 7987 4709
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4672 8263 4675
rect 8496 4672 8524 4768
rect 8251 4644 8524 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 6886 4576 7481 4604
rect 7469 4573 7481 4576
rect 7515 4604 7527 4607
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7515 4576 7573 4604
rect 7515 4573 7527 4576
rect 7469 4567 7527 4573
rect 7561 4573 7573 4576
rect 7607 4604 7619 4607
rect 8386 4604 8392 4616
rect 7607 4576 8392 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8588 4604 8616 4768
rect 9140 4681 9168 4780
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 10502 4768 10508 4820
rect 10560 4768 10566 4820
rect 10686 4768 10692 4820
rect 10744 4768 10750 4820
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 13722 4768 13728 4820
rect 13780 4768 13786 4820
rect 24026 4768 24032 4820
rect 24084 4768 24090 4820
rect 24397 4811 24455 4817
rect 24397 4777 24409 4811
rect 24443 4808 24455 4811
rect 24578 4808 24584 4820
rect 24443 4780 24584 4808
rect 24443 4777 24455 4780
rect 24397 4771 24455 4777
rect 24578 4768 24584 4780
rect 24636 4768 24642 4820
rect 26418 4808 26424 4820
rect 24826 4780 26424 4808
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 11333 4675 11391 4681
rect 11333 4641 11345 4675
rect 11379 4672 11391 4675
rect 11514 4672 11520 4684
rect 11379 4644 11520 4672
rect 11379 4641 11391 4644
rect 11333 4635 11391 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 12342 4632 12348 4684
rect 12400 4632 12406 4684
rect 13740 4672 13768 4768
rect 14366 4700 14372 4752
rect 14424 4740 14430 4752
rect 15657 4743 15715 4749
rect 14424 4712 14780 4740
rect 14424 4700 14430 4712
rect 14752 4681 14780 4712
rect 15657 4709 15669 4743
rect 15703 4709 15715 4743
rect 15657 4703 15715 4709
rect 17037 4743 17095 4749
rect 17037 4709 17049 4743
rect 17083 4740 17095 4743
rect 18690 4740 18696 4752
rect 17083 4712 18696 4740
rect 17083 4709 17095 4712
rect 17037 4703 17095 4709
rect 14093 4675 14151 4681
rect 14093 4672 14105 4675
rect 13740 4644 14105 4672
rect 14093 4641 14105 4644
rect 14139 4641 14151 4675
rect 14093 4635 14151 4641
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4641 14795 4675
rect 15672 4672 15700 4703
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 22925 4743 22983 4749
rect 22925 4709 22937 4743
rect 22971 4740 22983 4743
rect 22971 4712 23704 4740
rect 22971 4709 22983 4712
rect 22925 4703 22983 4709
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 15672 4644 16129 4672
rect 14737 4635 14795 4641
rect 16117 4641 16129 4644
rect 16163 4672 16175 4675
rect 23201 4675 23259 4681
rect 16163 4644 16574 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 9381 4607 9439 4613
rect 9381 4604 9393 4607
rect 8588 4576 9393 4604
rect 9381 4573 9393 4576
rect 9427 4573 9439 4607
rect 9381 4567 9439 4573
rect 11422 4564 11428 4616
rect 11480 4564 11486 4616
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 13814 4604 13820 4616
rect 13771 4576 13820 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 15930 4564 15936 4616
rect 15988 4564 15994 4616
rect 16546 4604 16574 4644
rect 23201 4641 23213 4675
rect 23247 4672 23259 4675
rect 23382 4672 23388 4684
rect 23247 4644 23388 4672
rect 23247 4641 23259 4644
rect 23201 4635 23259 4641
rect 23382 4632 23388 4644
rect 23440 4632 23446 4684
rect 23676 4681 23704 4712
rect 23661 4675 23719 4681
rect 23661 4641 23673 4675
rect 23707 4672 23719 4675
rect 24044 4672 24072 4768
rect 23707 4644 24072 4672
rect 23707 4641 23719 4644
rect 23661 4635 23719 4641
rect 16666 4604 16672 4616
rect 16546 4576 16672 4604
rect 16666 4564 16672 4576
rect 16724 4564 16730 4616
rect 17313 4607 17371 4613
rect 17313 4573 17325 4607
rect 17359 4604 17371 4607
rect 17681 4607 17739 4613
rect 17681 4604 17693 4607
rect 17359 4576 17693 4604
rect 17359 4573 17371 4576
rect 17313 4567 17371 4573
rect 17681 4573 17693 4576
rect 17727 4604 17739 4607
rect 24826 4604 24854 4780
rect 26418 4768 26424 4780
rect 26476 4768 26482 4820
rect 26786 4768 26792 4820
rect 26844 4808 26850 4820
rect 29086 4808 29092 4820
rect 26844 4780 29092 4808
rect 26844 4768 26850 4780
rect 29086 4768 29092 4780
rect 29144 4768 29150 4820
rect 30742 4768 30748 4820
rect 30800 4808 30806 4820
rect 31573 4811 31631 4817
rect 31573 4808 31585 4811
rect 30800 4780 31585 4808
rect 30800 4768 30806 4780
rect 31573 4777 31585 4780
rect 31619 4777 31631 4811
rect 31573 4771 31631 4777
rect 27617 4743 27675 4749
rect 27617 4709 27629 4743
rect 27663 4740 27675 4743
rect 27663 4712 29592 4740
rect 27663 4709 27675 4712
rect 27617 4703 27675 4709
rect 26510 4632 26516 4684
rect 26568 4672 26574 4684
rect 26789 4675 26847 4681
rect 26789 4672 26801 4675
rect 26568 4644 26801 4672
rect 26568 4632 26574 4644
rect 26789 4641 26801 4644
rect 26835 4672 26847 4675
rect 27706 4672 27712 4684
rect 26835 4644 27712 4672
rect 26835 4641 26847 4644
rect 26789 4635 26847 4641
rect 27706 4632 27712 4644
rect 27764 4632 27770 4684
rect 28902 4632 28908 4684
rect 28960 4632 28966 4684
rect 29564 4616 29592 4712
rect 30926 4632 30932 4684
rect 30984 4632 30990 4684
rect 32030 4632 32036 4684
rect 32088 4672 32094 4684
rect 32493 4675 32551 4681
rect 32493 4672 32505 4675
rect 32088 4644 32505 4672
rect 32088 4632 32094 4644
rect 32493 4641 32505 4644
rect 32539 4641 32551 4675
rect 32493 4635 32551 4641
rect 17727 4576 24854 4604
rect 17727 4573 17739 4576
rect 17681 4567 17739 4573
rect 15948 4536 15976 4564
rect 17328 4536 17356 4567
rect 24946 4564 24952 4616
rect 25004 4564 25010 4616
rect 25133 4607 25191 4613
rect 25133 4573 25145 4607
rect 25179 4573 25191 4607
rect 25133 4567 25191 4573
rect 15948 4508 17356 4536
rect 24854 4496 24860 4548
rect 24912 4536 24918 4548
rect 25148 4536 25176 4567
rect 25406 4564 25412 4616
rect 25464 4604 25470 4616
rect 25869 4607 25927 4613
rect 25869 4604 25881 4607
rect 25464 4576 25881 4604
rect 25464 4564 25470 4576
rect 25869 4573 25881 4576
rect 25915 4573 25927 4607
rect 25869 4567 25927 4573
rect 29273 4607 29331 4613
rect 29273 4573 29285 4607
rect 29319 4573 29331 4607
rect 29273 4567 29331 4573
rect 24912 4508 25176 4536
rect 26513 4539 26571 4545
rect 24912 4496 24918 4508
rect 26513 4505 26525 4539
rect 26559 4536 26571 4539
rect 27522 4536 27528 4548
rect 26559 4508 27528 4536
rect 26559 4505 26571 4508
rect 26513 4499 26571 4505
rect 27522 4496 27528 4508
rect 27580 4496 27586 4548
rect 27890 4496 27896 4548
rect 27948 4496 27954 4548
rect 29288 4536 29316 4567
rect 29546 4564 29552 4616
rect 29604 4564 29610 4616
rect 29730 4564 29736 4616
rect 29788 4604 29794 4616
rect 30653 4607 30711 4613
rect 30653 4604 30665 4607
rect 29788 4576 30665 4604
rect 29788 4564 29794 4576
rect 30653 4573 30665 4576
rect 30699 4573 30711 4607
rect 30653 4567 30711 4573
rect 32214 4564 32220 4616
rect 32272 4564 32278 4616
rect 31662 4536 31668 4548
rect 29288 4508 31668 4536
rect 31662 4496 31668 4508
rect 31720 4496 31726 4548
rect 31846 4496 31852 4548
rect 31904 4496 31910 4548
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 9582 4468 9588 4480
rect 8067 4440 9588 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 12986 4428 12992 4480
rect 13044 4428 13050 4480
rect 13081 4471 13139 4477
rect 13081 4437 13093 4471
rect 13127 4468 13139 4471
rect 13630 4468 13636 4480
rect 13127 4440 13636 4468
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 14458 4428 14464 4480
rect 14516 4468 14522 4480
rect 14553 4471 14611 4477
rect 14553 4468 14565 4471
rect 14516 4440 14565 4468
rect 14516 4428 14522 4440
rect 14553 4437 14565 4440
rect 14599 4437 14611 4471
rect 14553 4431 14611 4437
rect 15378 4428 15384 4480
rect 15436 4428 15442 4480
rect 15470 4428 15476 4480
rect 15528 4428 15534 4480
rect 16758 4428 16764 4480
rect 16816 4428 16822 4480
rect 16850 4428 16856 4480
rect 16908 4428 16914 4480
rect 22738 4428 22744 4480
rect 22796 4428 22802 4480
rect 24210 4428 24216 4480
rect 24268 4428 24274 4480
rect 25777 4471 25835 4477
rect 25777 4437 25789 4471
rect 25823 4468 25835 4471
rect 26050 4468 26056 4480
rect 25823 4440 26056 4468
rect 25823 4437 25835 4440
rect 25777 4431 25835 4437
rect 26050 4428 26056 4440
rect 26108 4428 26114 4480
rect 27338 4428 27344 4480
rect 27396 4428 27402 4480
rect 27433 4471 27491 4477
rect 27433 4437 27445 4471
rect 27479 4468 27491 4471
rect 27798 4468 27804 4480
rect 27479 4440 27804 4468
rect 27479 4437 27491 4440
rect 27433 4431 27491 4437
rect 27798 4428 27804 4440
rect 27856 4428 27862 4480
rect 30190 4428 30196 4480
rect 30248 4428 30254 4480
rect 1104 4378 34016 4400
rect 1104 4326 9138 4378
rect 9190 4326 9202 4378
rect 9254 4326 9266 4378
rect 9318 4326 9330 4378
rect 9382 4326 9394 4378
rect 9446 4326 17326 4378
rect 17378 4326 17390 4378
rect 17442 4326 17454 4378
rect 17506 4326 17518 4378
rect 17570 4326 17582 4378
rect 17634 4326 25514 4378
rect 25566 4326 25578 4378
rect 25630 4326 25642 4378
rect 25694 4326 25706 4378
rect 25758 4326 25770 4378
rect 25822 4326 33702 4378
rect 33754 4326 33766 4378
rect 33818 4326 33830 4378
rect 33882 4326 33894 4378
rect 33946 4326 33958 4378
rect 34010 4326 34016 4378
rect 1104 4304 34016 4326
rect 9490 4224 9496 4276
rect 9548 4224 9554 4276
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 10778 4264 10784 4276
rect 10735 4236 10784 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 10778 4224 10784 4236
rect 10836 4224 10842 4276
rect 12526 4224 12532 4276
rect 12584 4224 12590 4276
rect 13814 4224 13820 4276
rect 13872 4224 13878 4276
rect 24765 4267 24823 4273
rect 24765 4233 24777 4267
rect 24811 4264 24823 4267
rect 24946 4264 24952 4276
rect 24811 4236 24952 4264
rect 24811 4233 24823 4236
rect 24765 4227 24823 4233
rect 24946 4224 24952 4236
rect 25004 4224 25010 4276
rect 27893 4267 27951 4273
rect 27893 4233 27905 4267
rect 27939 4264 27951 4267
rect 28166 4264 28172 4276
rect 27939 4236 28172 4264
rect 27939 4233 27951 4236
rect 27893 4227 27951 4233
rect 28166 4224 28172 4236
rect 28224 4224 28230 4276
rect 29270 4224 29276 4276
rect 29328 4264 29334 4276
rect 29549 4267 29607 4273
rect 29549 4264 29561 4267
rect 29328 4236 29561 4264
rect 29328 4224 29334 4236
rect 29549 4233 29561 4236
rect 29595 4233 29607 4267
rect 29549 4227 29607 4233
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2958 4128 2964 4140
rect 2731 4100 2964 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6595 4100 6684 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4029 2467 4063
rect 2409 4023 2467 4029
rect 2424 3924 2452 4023
rect 6656 3936 6684 4100
rect 7834 4088 7840 4140
rect 7892 4088 7898 4140
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4128 9367 4131
rect 9508 4128 9536 4224
rect 12544 4196 12572 4224
rect 12452 4168 12572 4196
rect 24826 4168 27108 4196
rect 9582 4137 9588 4140
rect 9355 4100 9536 4128
rect 9355 4097 9367 4100
rect 9309 4091 9367 4097
rect 9576 4091 9588 4137
rect 9640 4128 9646 4140
rect 10873 4131 10931 4137
rect 9640 4100 9676 4128
rect 9582 4088 9588 4091
rect 9640 4088 9646 4100
rect 10873 4097 10885 4131
rect 10919 4128 10931 4131
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 10919 4100 11805 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 11793 4097 11805 4100
rect 11839 4128 11851 4131
rect 12452 4128 12480 4168
rect 11839 4100 12480 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 15378 4088 15384 4140
rect 15436 4128 15442 4140
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 15436 4100 15485 4128
rect 15436 4088 15442 4100
rect 15473 4097 15485 4100
rect 15519 4097 15531 4131
rect 15473 4091 15531 4097
rect 16758 4088 16764 4140
rect 16816 4088 16822 4140
rect 18690 4088 18696 4140
rect 18748 4128 18754 4140
rect 18877 4131 18935 4137
rect 18877 4128 18889 4131
rect 18748 4100 18889 4128
rect 18748 4088 18754 4100
rect 18877 4097 18889 4100
rect 18923 4097 18935 4131
rect 18877 4091 18935 4097
rect 23652 4131 23710 4137
rect 23652 4097 23664 4131
rect 23698 4128 23710 4131
rect 24394 4128 24400 4140
rect 23698 4100 24400 4128
rect 23698 4097 23710 4100
rect 23652 4091 23710 4097
rect 24394 4088 24400 4100
rect 24452 4088 24458 4140
rect 24578 4088 24584 4140
rect 24636 4128 24642 4140
rect 24826 4128 24854 4168
rect 24636 4100 24854 4128
rect 26237 4131 26295 4137
rect 24636 4088 24642 4100
rect 26237 4097 26249 4131
rect 26283 4128 26295 4131
rect 26878 4128 26884 4140
rect 26283 4100 26884 4128
rect 26283 4097 26295 4100
rect 26237 4091 26295 4097
rect 26878 4088 26884 4100
rect 26936 4088 26942 4140
rect 6730 4020 6736 4072
rect 6788 4060 6794 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6788 4032 6837 4060
rect 6788 4020 6794 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 7800 4032 8309 4060
rect 7800 4020 7806 4032
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 8297 4023 8355 4029
rect 12618 4020 12624 4072
rect 12676 4020 12682 4072
rect 13078 4020 13084 4072
rect 13136 4060 13142 4072
rect 13173 4063 13231 4069
rect 13173 4060 13185 4063
rect 13136 4032 13185 4060
rect 13136 4020 13142 4032
rect 13173 4029 13185 4032
rect 13219 4029 13231 4063
rect 13173 4023 13231 4029
rect 14090 4020 14096 4072
rect 14148 4020 14154 4072
rect 16022 4020 16028 4072
rect 16080 4020 16086 4072
rect 17034 4020 17040 4072
rect 17092 4020 17098 4072
rect 19518 4020 19524 4072
rect 19576 4020 19582 4072
rect 22741 4063 22799 4069
rect 22741 4029 22753 4063
rect 22787 4060 22799 4063
rect 23198 4060 23204 4072
rect 22787 4032 23204 4060
rect 22787 4029 22799 4032
rect 22741 4023 22799 4029
rect 23198 4020 23204 4032
rect 23256 4020 23262 4072
rect 23385 4063 23443 4069
rect 23385 4029 23397 4063
rect 23431 4029 23443 4063
rect 23385 4023 23443 4029
rect 11241 3995 11299 4001
rect 11241 3961 11253 3995
rect 11287 3992 11299 3995
rect 13630 3992 13636 4004
rect 11287 3964 13636 3992
rect 11287 3961 11299 3964
rect 11241 3955 11299 3961
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 23400 3936 23428 4023
rect 24762 4020 24768 4072
rect 24820 4060 24826 4072
rect 25041 4063 25099 4069
rect 25041 4060 25053 4063
rect 24820 4032 25053 4060
rect 24820 4020 24826 4032
rect 25041 4029 25053 4032
rect 25087 4029 25099 4063
rect 25041 4023 25099 4029
rect 26326 4020 26332 4072
rect 26384 4020 26390 4072
rect 27080 4069 27108 4168
rect 28736 4168 30972 4196
rect 28736 4140 28764 4168
rect 28718 4088 28724 4140
rect 28776 4088 28782 4140
rect 28994 4088 29000 4140
rect 29052 4137 29058 4140
rect 29288 4137 29316 4168
rect 29052 4128 29064 4137
rect 29273 4131 29331 4137
rect 29052 4100 29097 4128
rect 29052 4091 29064 4100
rect 29273 4097 29285 4131
rect 29319 4097 29331 4131
rect 29273 4091 29331 4097
rect 30673 4131 30731 4137
rect 30673 4097 30685 4131
rect 30719 4128 30731 4131
rect 30834 4128 30840 4140
rect 30719 4100 30840 4128
rect 30719 4097 30731 4100
rect 30673 4091 30731 4097
rect 29052 4088 29058 4091
rect 30834 4088 30840 4100
rect 30892 4088 30898 4140
rect 30944 4137 30972 4168
rect 31754 4156 31760 4208
rect 31812 4196 31818 4208
rect 31812 4168 32260 4196
rect 31812 4156 31818 4168
rect 30929 4131 30987 4137
rect 30929 4097 30941 4131
rect 30975 4128 30987 4131
rect 32122 4128 32128 4140
rect 30975 4100 32128 4128
rect 30975 4097 30987 4100
rect 30929 4091 30987 4097
rect 32122 4088 32128 4100
rect 32180 4088 32186 4140
rect 32232 4137 32260 4168
rect 32217 4131 32275 4137
rect 32217 4097 32229 4131
rect 32263 4097 32275 4131
rect 32217 4091 32275 4097
rect 26789 4063 26847 4069
rect 26789 4029 26801 4063
rect 26835 4029 26847 4063
rect 26789 4023 26847 4029
rect 27065 4063 27123 4069
rect 27065 4029 27077 4063
rect 27111 4060 27123 4063
rect 27154 4060 27160 4072
rect 27111 4032 27160 4060
rect 27111 4029 27123 4032
rect 27065 4023 27123 4029
rect 26344 3992 26372 4020
rect 24320 3964 26372 3992
rect 2590 3924 2596 3936
rect 2424 3896 2596 3924
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 6638 3884 6644 3936
rect 6696 3884 6702 3936
rect 11330 3884 11336 3936
rect 11388 3884 11394 3936
rect 14642 3884 14648 3936
rect 14700 3884 14706 3936
rect 18138 3884 18144 3936
rect 18196 3884 18202 3936
rect 23290 3884 23296 3936
rect 23348 3884 23354 3936
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 24320 3924 24348 3964
rect 26510 3952 26516 4004
rect 26568 3952 26574 4004
rect 26804 3992 26832 4023
rect 27154 4020 27160 4032
rect 27212 4020 27218 4072
rect 27890 4020 27896 4072
rect 27948 4020 27954 4072
rect 31110 4020 31116 4072
rect 31168 4060 31174 4072
rect 31573 4063 31631 4069
rect 31573 4060 31585 4063
rect 31168 4032 31585 4060
rect 31168 4020 31174 4032
rect 31573 4029 31585 4032
rect 31619 4029 31631 4063
rect 31573 4023 31631 4029
rect 31662 4020 31668 4072
rect 31720 4060 31726 4072
rect 32493 4063 32551 4069
rect 32493 4060 32505 4063
rect 31720 4032 32505 4060
rect 31720 4020 31726 4032
rect 32493 4029 32505 4032
rect 32539 4029 32551 4063
rect 32493 4023 32551 4029
rect 27908 3992 27936 4020
rect 26804 3964 27936 3992
rect 27080 3936 27108 3964
rect 23440 3896 24348 3924
rect 23440 3884 23446 3896
rect 26234 3884 26240 3936
rect 26292 3924 26298 3936
rect 26329 3927 26387 3933
rect 26329 3924 26341 3927
rect 26292 3896 26341 3924
rect 26292 3884 26298 3896
rect 26329 3893 26341 3896
rect 26375 3893 26387 3927
rect 26329 3887 26387 3893
rect 27062 3884 27068 3936
rect 27120 3884 27126 3936
rect 27614 3884 27620 3936
rect 27672 3884 27678 3936
rect 29546 3884 29552 3936
rect 29604 3924 29610 3936
rect 31021 3927 31079 3933
rect 31021 3924 31033 3927
rect 29604 3896 31033 3924
rect 29604 3884 29610 3896
rect 31021 3893 31033 3896
rect 31067 3893 31079 3927
rect 31021 3887 31079 3893
rect 1104 3834 33856 3856
rect 1104 3782 5044 3834
rect 5096 3782 5108 3834
rect 5160 3782 5172 3834
rect 5224 3782 5236 3834
rect 5288 3782 5300 3834
rect 5352 3782 13232 3834
rect 13284 3782 13296 3834
rect 13348 3782 13360 3834
rect 13412 3782 13424 3834
rect 13476 3782 13488 3834
rect 13540 3782 21420 3834
rect 21472 3782 21484 3834
rect 21536 3782 21548 3834
rect 21600 3782 21612 3834
rect 21664 3782 21676 3834
rect 21728 3782 29608 3834
rect 29660 3782 29672 3834
rect 29724 3782 29736 3834
rect 29788 3782 29800 3834
rect 29852 3782 29864 3834
rect 29916 3782 33856 3834
rect 1104 3760 33856 3782
rect 8938 3720 8944 3732
rect 6886 3692 8944 3720
rect 1578 3544 1584 3596
rect 1636 3544 1642 3596
rect 6638 3544 6644 3596
rect 6696 3544 6702 3596
rect 2590 3476 2596 3528
rect 2648 3476 2654 3528
rect 5721 3519 5779 3525
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 6886 3516 6914 3692
rect 8938 3680 8944 3692
rect 8996 3680 9002 3732
rect 10152 3692 11468 3720
rect 10152 3652 10180 3692
rect 7208 3624 10180 3652
rect 11440 3652 11468 3692
rect 11514 3680 11520 3732
rect 11572 3680 11578 3732
rect 13906 3720 13912 3732
rect 12084 3692 13912 3720
rect 12084 3652 12112 3692
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 14090 3680 14096 3732
rect 14148 3680 14154 3732
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 19889 3723 19947 3729
rect 19889 3720 19901 3723
rect 19576 3692 19901 3720
rect 19576 3680 19582 3692
rect 19889 3689 19901 3692
rect 19935 3689 19947 3723
rect 19889 3683 19947 3689
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 23382 3720 23388 3732
rect 22143 3692 23388 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 11440 3624 12112 3652
rect 18417 3655 18475 3661
rect 7208 3525 7236 3624
rect 18417 3621 18429 3655
rect 18463 3652 18475 3655
rect 18463 3624 19288 3652
rect 18463 3621 18475 3624
rect 18417 3615 18475 3621
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 9548 3556 10149 3584
rect 9548 3544 9554 3556
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 5767 3488 6914 3516
rect 7193 3519 7251 3525
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 7193 3485 7205 3519
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 8662 3476 8668 3528
rect 8720 3476 8726 3528
rect 9858 3476 9864 3528
rect 9916 3516 9922 3528
rect 9953 3519 10011 3525
rect 9953 3516 9965 3519
rect 9916 3488 9965 3516
rect 9916 3476 9922 3488
rect 9953 3485 9965 3488
rect 9999 3485 10011 3519
rect 10152 3516 10180 3547
rect 13630 3544 13636 3596
rect 13688 3544 13694 3596
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 19260 3593 19288 3624
rect 22204 3596 22232 3692
rect 23382 3680 23388 3692
rect 23440 3680 23446 3732
rect 24302 3720 24308 3732
rect 24044 3692 24308 3720
rect 24044 3661 24072 3692
rect 24302 3680 24308 3692
rect 24360 3680 24366 3732
rect 24394 3680 24400 3732
rect 24452 3680 24458 3732
rect 24578 3720 24584 3732
rect 24504 3692 24584 3720
rect 24504 3661 24532 3692
rect 24578 3680 24584 3692
rect 24636 3680 24642 3732
rect 24854 3720 24860 3732
rect 24826 3680 24860 3720
rect 24912 3680 24918 3732
rect 24949 3723 25007 3729
rect 24949 3689 24961 3723
rect 24995 3720 25007 3723
rect 25406 3720 25412 3732
rect 24995 3692 25412 3720
rect 24995 3689 25007 3692
rect 24949 3683 25007 3689
rect 25406 3680 25412 3692
rect 25464 3680 25470 3732
rect 27338 3680 27344 3732
rect 27396 3680 27402 3732
rect 31846 3680 31852 3732
rect 31904 3720 31910 3732
rect 32585 3723 32643 3729
rect 32585 3720 32597 3723
rect 31904 3692 32597 3720
rect 31904 3680 31910 3692
rect 32585 3689 32597 3692
rect 32631 3689 32643 3723
rect 32585 3683 32643 3689
rect 32858 3680 32864 3732
rect 32916 3680 32922 3732
rect 23569 3655 23627 3661
rect 23569 3621 23581 3655
rect 23615 3621 23627 3655
rect 23569 3615 23627 3621
rect 24029 3655 24087 3661
rect 24029 3621 24041 3655
rect 24075 3621 24087 3655
rect 24029 3615 24087 3621
rect 24489 3655 24547 3661
rect 24489 3621 24501 3655
rect 24535 3621 24547 3655
rect 24489 3615 24547 3621
rect 19245 3587 19303 3593
rect 16632 3556 17172 3584
rect 16632 3544 16638 3556
rect 12986 3516 12992 3528
rect 10152 3488 12992 3516
rect 9953 3479 10011 3485
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 15473 3519 15531 3525
rect 15473 3516 15485 3519
rect 13740 3488 15485 3516
rect 5353 3451 5411 3457
rect 5353 3417 5365 3451
rect 5399 3448 5411 3451
rect 5399 3420 6040 3448
rect 5399 3417 5411 3420
rect 5353 3411 5411 3417
rect 6012 3392 6040 3420
rect 8294 3408 8300 3460
rect 8352 3408 8358 3460
rect 10226 3408 10232 3460
rect 10284 3448 10290 3460
rect 10382 3451 10440 3457
rect 10382 3448 10394 3451
rect 10284 3420 10394 3448
rect 10284 3408 10290 3420
rect 10382 3417 10394 3420
rect 10428 3417 10440 3451
rect 10382 3411 10440 3417
rect 11330 3408 11336 3460
rect 11388 3448 11394 3460
rect 12722 3451 12780 3457
rect 12722 3448 12734 3451
rect 11388 3420 12734 3448
rect 11388 3408 11394 3420
rect 12722 3417 12734 3420
rect 12768 3417 12780 3451
rect 13004 3448 13032 3476
rect 13740 3448 13768 3488
rect 15473 3485 15485 3488
rect 15519 3516 15531 3519
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 15519 3488 15577 3516
rect 15519 3485 15531 3488
rect 15473 3479 15531 3485
rect 15565 3485 15577 3488
rect 15611 3516 15623 3519
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 15611 3488 17049 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 17037 3485 17049 3488
rect 17083 3485 17095 3519
rect 17144 3516 17172 3556
rect 19245 3553 19257 3587
rect 19291 3553 19303 3587
rect 19245 3547 19303 3553
rect 22186 3544 22192 3596
rect 22244 3544 22250 3596
rect 23584 3584 23612 3615
rect 24826 3584 24854 3680
rect 23584 3556 24854 3584
rect 26881 3587 26939 3593
rect 26881 3553 26893 3587
rect 26927 3553 26939 3587
rect 26881 3547 26939 3553
rect 17293 3519 17351 3525
rect 17293 3516 17305 3519
rect 17144 3488 17305 3516
rect 17037 3479 17095 3485
rect 17293 3485 17305 3488
rect 17339 3485 17351 3519
rect 17293 3479 17351 3485
rect 20346 3476 20352 3528
rect 20404 3476 20410 3528
rect 22456 3519 22514 3525
rect 22456 3485 22468 3519
rect 22502 3516 22514 3519
rect 22738 3516 22744 3528
rect 22502 3488 22744 3516
rect 22502 3485 22514 3488
rect 22456 3479 22514 3485
rect 22738 3476 22744 3488
rect 22796 3476 22802 3528
rect 22922 3476 22928 3528
rect 22980 3516 22986 3528
rect 24762 3516 24768 3528
rect 22980 3488 24768 3516
rect 22980 3476 22986 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 24857 3519 24915 3525
rect 24857 3485 24869 3519
rect 24903 3512 24915 3519
rect 25314 3516 25320 3528
rect 24964 3512 25320 3516
rect 24903 3488 25320 3512
rect 24903 3485 24992 3488
rect 24857 3484 24992 3485
rect 24857 3479 24915 3484
rect 13004 3420 13768 3448
rect 15228 3451 15286 3457
rect 12722 3411 12780 3417
rect 15228 3417 15240 3451
rect 15274 3448 15286 3451
rect 15832 3451 15890 3457
rect 15274 3420 15516 3448
rect 15274 3417 15286 3420
rect 15228 3411 15286 3417
rect 15488 3392 15516 3420
rect 15832 3417 15844 3451
rect 15878 3448 15890 3451
rect 16850 3448 16856 3460
rect 15878 3420 16856 3448
rect 15878 3417 15890 3420
rect 15832 3411 15890 3417
rect 16850 3408 16856 3420
rect 16908 3408 16914 3460
rect 20901 3451 20959 3457
rect 20901 3417 20913 3451
rect 20947 3448 20959 3451
rect 21910 3448 21916 3460
rect 20947 3420 21916 3448
rect 20947 3417 20959 3420
rect 20901 3411 20959 3417
rect 21910 3408 21916 3420
rect 21968 3408 21974 3460
rect 23382 3408 23388 3460
rect 23440 3448 23446 3460
rect 23661 3451 23719 3457
rect 23661 3448 23673 3451
rect 23440 3420 23673 3448
rect 23440 3408 23446 3420
rect 23661 3417 23673 3420
rect 23707 3448 23719 3451
rect 24872 3448 24900 3479
rect 25314 3476 25320 3488
rect 25372 3476 25378 3528
rect 26073 3519 26131 3525
rect 26073 3485 26085 3519
rect 26119 3516 26131 3519
rect 26234 3516 26240 3528
rect 26119 3488 26240 3516
rect 26119 3485 26131 3488
rect 26073 3479 26131 3485
rect 26234 3476 26240 3488
rect 26292 3476 26298 3528
rect 26326 3476 26332 3528
rect 26384 3476 26390 3528
rect 26418 3476 26424 3528
rect 26476 3476 26482 3528
rect 23707 3420 24900 3448
rect 23707 3417 23719 3420
rect 23661 3411 23719 3417
rect 5994 3340 6000 3392
rect 6052 3340 6058 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 9401 3383 9459 3389
rect 9401 3380 9413 3383
rect 8168 3352 9413 3380
rect 8168 3340 8174 3352
rect 9401 3349 9413 3352
rect 9447 3349 9459 3383
rect 9401 3343 9459 3349
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 12894 3340 12900 3392
rect 12952 3380 12958 3392
rect 13081 3383 13139 3389
rect 13081 3380 13093 3383
rect 12952 3352 13093 3380
rect 12952 3340 12958 3352
rect 13081 3349 13093 3352
rect 13127 3349 13139 3383
rect 13081 3343 13139 3349
rect 15470 3340 15476 3392
rect 15528 3340 15534 3392
rect 16942 3340 16948 3392
rect 17000 3340 17006 3392
rect 24118 3340 24124 3392
rect 24176 3340 24182 3392
rect 24486 3340 24492 3392
rect 24544 3380 24550 3392
rect 26896 3380 26924 3547
rect 27356 3516 27384 3680
rect 30006 3612 30012 3664
rect 30064 3652 30070 3664
rect 30064 3624 30374 3652
rect 30064 3612 30070 3624
rect 30346 3584 30374 3624
rect 33413 3587 33471 3593
rect 33413 3584 33425 3587
rect 30346 3556 33425 3584
rect 33413 3553 33425 3556
rect 33459 3553 33471 3587
rect 33413 3547 33471 3553
rect 27985 3519 28043 3525
rect 27985 3516 27997 3519
rect 27356 3488 27997 3516
rect 27985 3485 27997 3488
rect 28031 3485 28043 3519
rect 27985 3479 28043 3485
rect 28537 3519 28595 3525
rect 28537 3485 28549 3519
rect 28583 3516 28595 3519
rect 29914 3516 29920 3528
rect 28583 3488 29920 3516
rect 28583 3485 28595 3488
rect 28537 3479 28595 3485
rect 29914 3476 29920 3488
rect 29972 3476 29978 3528
rect 30190 3476 30196 3528
rect 30248 3476 30254 3528
rect 31754 3476 31760 3528
rect 31812 3476 31818 3528
rect 31938 3476 31944 3528
rect 31996 3516 32002 3528
rect 32125 3519 32183 3525
rect 32125 3516 32137 3519
rect 31996 3488 32137 3516
rect 31996 3476 32002 3488
rect 32125 3485 32137 3488
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 32769 3519 32827 3525
rect 32769 3485 32781 3519
rect 32815 3516 32827 3519
rect 32815 3488 33548 3516
rect 32815 3485 32827 3488
rect 32769 3479 32827 3485
rect 29825 3451 29883 3457
rect 29825 3417 29837 3451
rect 29871 3448 29883 3451
rect 31110 3448 31116 3460
rect 29871 3420 31116 3448
rect 29871 3417 29883 3420
rect 29825 3411 29883 3417
rect 31110 3408 31116 3420
rect 31168 3408 31174 3460
rect 33520 3392 33548 3488
rect 24544 3352 26924 3380
rect 24544 3340 24550 3352
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28997 3383 29055 3389
rect 28997 3380 29009 3383
rect 27948 3352 29009 3380
rect 27948 3340 27954 3352
rect 28997 3349 29009 3352
rect 29043 3380 29055 3383
rect 29365 3383 29423 3389
rect 29365 3380 29377 3383
rect 29043 3352 29377 3380
rect 29043 3349 29055 3352
rect 28997 3343 29055 3349
rect 29365 3349 29377 3352
rect 29411 3380 29423 3383
rect 30653 3383 30711 3389
rect 30653 3380 30665 3383
rect 29411 3352 30665 3380
rect 29411 3349 29423 3352
rect 29365 3343 29423 3349
rect 30653 3349 30665 3352
rect 30699 3380 30711 3383
rect 31297 3383 31355 3389
rect 31297 3380 31309 3383
rect 30699 3352 31309 3380
rect 30699 3349 30711 3352
rect 30653 3343 30711 3349
rect 31297 3349 31309 3352
rect 31343 3380 31355 3383
rect 31846 3380 31852 3392
rect 31343 3352 31852 3380
rect 31343 3349 31355 3352
rect 31297 3343 31355 3349
rect 31846 3340 31852 3352
rect 31904 3340 31910 3392
rect 33502 3340 33508 3392
rect 33560 3340 33566 3392
rect 1104 3290 34016 3312
rect 1104 3238 9138 3290
rect 9190 3238 9202 3290
rect 9254 3238 9266 3290
rect 9318 3238 9330 3290
rect 9382 3238 9394 3290
rect 9446 3238 17326 3290
rect 17378 3238 17390 3290
rect 17442 3238 17454 3290
rect 17506 3238 17518 3290
rect 17570 3238 17582 3290
rect 17634 3238 25514 3290
rect 25566 3238 25578 3290
rect 25630 3238 25642 3290
rect 25694 3238 25706 3290
rect 25758 3238 25770 3290
rect 25822 3238 33702 3290
rect 33754 3238 33766 3290
rect 33818 3238 33830 3290
rect 33882 3238 33894 3290
rect 33946 3238 33958 3290
rect 34010 3238 34016 3290
rect 1104 3216 34016 3238
rect 8294 3136 8300 3188
rect 8352 3136 8358 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3176 9919 3179
rect 11422 3176 11428 3188
rect 9907 3148 11428 3176
rect 9907 3145 9919 3148
rect 9861 3139 9919 3145
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 12894 3136 12900 3188
rect 12952 3136 12958 3188
rect 12986 3136 12992 3188
rect 13044 3136 13050 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 13173 3179 13231 3185
rect 13173 3176 13185 3179
rect 13136 3148 13185 3176
rect 13136 3136 13142 3148
rect 13173 3145 13185 3148
rect 13219 3145 13231 3179
rect 13173 3139 13231 3145
rect 16022 3136 16028 3188
rect 16080 3136 16086 3188
rect 16666 3136 16672 3188
rect 16724 3136 16730 3188
rect 18138 3136 18144 3188
rect 18196 3136 18202 3188
rect 22186 3136 22192 3188
rect 22244 3176 22250 3188
rect 22281 3179 22339 3185
rect 22281 3176 22293 3179
rect 22244 3148 22293 3176
rect 22244 3136 22250 3148
rect 22281 3145 22293 3148
rect 22327 3145 22339 3179
rect 22281 3139 22339 3145
rect 23198 3136 23204 3188
rect 23256 3176 23262 3188
rect 23256 3148 24072 3176
rect 23256 3136 23262 3148
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3040 2743 3043
rect 3418 3040 3424 3052
rect 2731 3012 3424 3040
rect 2731 3009 2743 3012
rect 2685 3003 2743 3009
rect 3418 3000 3424 3012
rect 3476 3000 3482 3052
rect 5994 3000 6000 3052
rect 6052 3000 6058 3052
rect 8312 3049 8340 3136
rect 8496 3080 9536 3108
rect 8496 3049 8524 3080
rect 9508 3052 9536 3080
rect 8754 3049 8760 3052
rect 8297 3043 8355 3049
rect 8297 3009 8309 3043
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3009 8539 3043
rect 8748 3040 8760 3049
rect 8715 3012 8760 3040
rect 8481 3003 8539 3009
rect 8748 3003 8760 3012
rect 8754 3000 8760 3003
rect 8812 3000 8818 3052
rect 9490 3000 9496 3052
rect 9548 3000 9554 3052
rect 9950 3000 9956 3052
rect 10008 3000 10014 3052
rect 12912 3040 12940 3136
rect 13004 3108 13032 3136
rect 13004 3080 14596 3108
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12912 3012 13001 3040
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 12989 3003 13047 3009
rect 14297 3043 14355 3049
rect 14297 3009 14309 3043
rect 14343 3040 14355 3043
rect 14458 3040 14464 3052
rect 14343 3012 14464 3040
rect 14343 3009 14355 3012
rect 14297 3003 14355 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14568 3049 14596 3080
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 16040 3040 16068 3136
rect 18156 3049 18184 3136
rect 23124 3080 23704 3108
rect 16301 3043 16359 3049
rect 16301 3040 16313 3043
rect 16040 3012 16313 3040
rect 14553 3003 14611 3009
rect 16301 3009 16313 3012
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3009 18199 3043
rect 18141 3003 18199 3009
rect 19702 3000 19708 3052
rect 19760 3000 19766 3052
rect 23124 3049 23152 3080
rect 23676 3052 23704 3080
rect 23109 3043 23167 3049
rect 23109 3009 23121 3043
rect 23155 3009 23167 3043
rect 23109 3003 23167 3009
rect 23293 3043 23351 3049
rect 23293 3009 23305 3043
rect 23339 3009 23351 3043
rect 23293 3003 23351 3009
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 2590 2972 2596 2984
rect 2455 2944 2596 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 2590 2932 2596 2944
rect 2648 2932 2654 2984
rect 4982 2932 4988 2984
rect 5040 2932 5046 2984
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 7944 2836 7972 2935
rect 10502 2932 10508 2984
rect 10560 2932 10566 2984
rect 12526 2932 12532 2984
rect 12584 2932 12590 2984
rect 14826 2932 14832 2984
rect 14884 2972 14890 2984
rect 15289 2975 15347 2981
rect 15289 2972 15301 2975
rect 14884 2944 15301 2972
rect 14884 2932 14890 2944
rect 15289 2941 15301 2944
rect 15335 2941 15347 2975
rect 15289 2935 15347 2941
rect 17310 2932 17316 2984
rect 17368 2932 17374 2984
rect 17678 2932 17684 2984
rect 17736 2932 17742 2984
rect 18782 2932 18788 2984
rect 18840 2972 18846 2984
rect 19981 2975 20039 2981
rect 19981 2972 19993 2975
rect 18840 2944 19993 2972
rect 18840 2932 18846 2944
rect 19981 2941 19993 2944
rect 20027 2941 20039 2975
rect 19981 2935 20039 2941
rect 22833 2975 22891 2981
rect 22833 2941 22845 2975
rect 22879 2972 22891 2975
rect 23308 2972 23336 3003
rect 23658 3000 23664 3052
rect 23716 3000 23722 3052
rect 22879 2944 23336 2972
rect 23753 2975 23811 2981
rect 22879 2941 22891 2944
rect 22833 2935 22891 2941
rect 23753 2941 23765 2975
rect 23799 2941 23811 2975
rect 23753 2935 23811 2941
rect 21818 2864 21824 2916
rect 21876 2904 21882 2916
rect 23768 2904 23796 2935
rect 21876 2876 23796 2904
rect 24044 2904 24072 3148
rect 24118 3136 24124 3188
rect 24176 3136 24182 3188
rect 26970 3136 26976 3188
rect 27028 3136 27034 3188
rect 30834 3136 30840 3188
rect 30892 3176 30898 3188
rect 31389 3179 31447 3185
rect 31389 3176 31401 3179
rect 30892 3148 31401 3176
rect 30892 3136 30898 3148
rect 31389 3145 31401 3148
rect 31435 3145 31447 3179
rect 31389 3139 31447 3145
rect 32582 3136 32588 3188
rect 32640 3176 32646 3188
rect 33505 3179 33563 3185
rect 33505 3176 33517 3179
rect 32640 3148 33517 3176
rect 32640 3136 32646 3148
rect 33505 3145 33517 3148
rect 33551 3145 33563 3179
rect 33505 3139 33563 3145
rect 24136 3108 24164 3136
rect 25878 3111 25936 3117
rect 25878 3108 25890 3111
rect 24136 3080 25890 3108
rect 25878 3077 25890 3080
rect 25924 3077 25936 3111
rect 26326 3108 26332 3120
rect 25878 3071 25936 3077
rect 26160 3080 26332 3108
rect 26160 3049 26188 3080
rect 26326 3068 26332 3080
rect 26384 3108 26390 3120
rect 26384 3080 28396 3108
rect 26384 3068 26390 3080
rect 26145 3043 26203 3049
rect 26145 3009 26157 3043
rect 26191 3009 26203 3043
rect 26145 3003 26203 3009
rect 27062 3000 27068 3052
rect 27120 3000 27126 3052
rect 27798 3000 27804 3052
rect 27856 3040 27862 3052
rect 28086 3043 28144 3049
rect 28086 3040 28098 3043
rect 27856 3012 28098 3040
rect 27856 3000 27862 3012
rect 28086 3009 28098 3012
rect 28132 3009 28144 3043
rect 28086 3003 28144 3009
rect 26326 2932 26332 2984
rect 26384 2972 26390 2984
rect 27080 2972 27108 3000
rect 28368 2984 28396 3080
rect 31846 3068 31852 3120
rect 31904 3068 31910 3120
rect 29825 3043 29883 3049
rect 29825 3009 29837 3043
rect 29871 3009 29883 3043
rect 29825 3003 29883 3009
rect 26384 2944 27108 2972
rect 26384 2932 26390 2944
rect 28350 2932 28356 2984
rect 28408 2932 28414 2984
rect 28626 2932 28632 2984
rect 28684 2932 28690 2984
rect 29840 2972 29868 3003
rect 29914 3000 29920 3052
rect 29972 3000 29978 3052
rect 32122 3000 32128 3052
rect 32180 3000 32186 3052
rect 32381 3043 32439 3049
rect 32381 3040 32393 3043
rect 32232 3012 32393 3040
rect 30006 2972 30012 2984
rect 29840 2944 30012 2972
rect 30006 2932 30012 2944
rect 30064 2932 30070 2984
rect 30190 2932 30196 2984
rect 30248 2972 30254 2984
rect 30377 2975 30435 2981
rect 30377 2972 30389 2975
rect 30248 2944 30389 2972
rect 30248 2932 30254 2944
rect 30377 2941 30389 2944
rect 30423 2941 30435 2975
rect 32232 2972 32260 3012
rect 32381 3009 32393 3012
rect 32427 3009 32439 3043
rect 32381 3003 32439 3009
rect 30377 2935 30435 2941
rect 31588 2944 32260 2972
rect 24765 2907 24823 2913
rect 24765 2904 24777 2907
rect 24044 2876 24777 2904
rect 21876 2864 21882 2876
rect 24765 2873 24777 2876
rect 24811 2873 24823 2907
rect 24765 2867 24823 2873
rect 26694 2864 26700 2916
rect 26752 2864 26758 2916
rect 28810 2864 28816 2916
rect 28868 2904 28874 2916
rect 31481 2907 31539 2913
rect 31481 2904 31493 2907
rect 28868 2876 31493 2904
rect 28868 2864 28874 2876
rect 31481 2873 31493 2876
rect 31527 2873 31539 2907
rect 31481 2867 31539 2873
rect 9122 2836 9128 2848
rect 7944 2808 9128 2836
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 26789 2839 26847 2845
rect 26789 2805 26801 2839
rect 26835 2836 26847 2839
rect 31588 2836 31616 2944
rect 26835 2808 31616 2836
rect 26835 2805 26847 2808
rect 26789 2799 26847 2805
rect 1104 2746 33856 2768
rect 1104 2694 5044 2746
rect 5096 2694 5108 2746
rect 5160 2694 5172 2746
rect 5224 2694 5236 2746
rect 5288 2694 5300 2746
rect 5352 2694 13232 2746
rect 13284 2694 13296 2746
rect 13348 2694 13360 2746
rect 13412 2694 13424 2746
rect 13476 2694 13488 2746
rect 13540 2694 21420 2746
rect 21472 2694 21484 2746
rect 21536 2694 21548 2746
rect 21600 2694 21612 2746
rect 21664 2694 21676 2746
rect 21728 2694 29608 2746
rect 29660 2694 29672 2746
rect 29724 2694 29736 2746
rect 29788 2694 29800 2746
rect 29852 2694 29864 2746
rect 29916 2694 33856 2746
rect 1104 2672 33856 2694
rect 12434 2592 12440 2644
rect 12492 2592 12498 2644
rect 14366 2592 14372 2644
rect 14424 2592 14430 2644
rect 17310 2592 17316 2644
rect 17368 2592 17374 2644
rect 19058 2592 19064 2644
rect 19116 2632 19122 2644
rect 29546 2632 29552 2644
rect 19116 2604 29552 2632
rect 19116 2592 19122 2604
rect 29546 2592 29552 2604
rect 29604 2592 29610 2644
rect 31665 2635 31723 2641
rect 31665 2601 31677 2635
rect 31711 2632 31723 2635
rect 31754 2632 31760 2644
rect 31711 2604 31760 2632
rect 31711 2601 31723 2604
rect 31665 2595 31723 2601
rect 31754 2592 31760 2604
rect 31812 2592 31818 2644
rect 2498 2524 2504 2576
rect 2556 2564 2562 2576
rect 2869 2567 2927 2573
rect 2869 2564 2881 2567
rect 2556 2536 2881 2564
rect 2556 2524 2562 2536
rect 2869 2533 2881 2536
rect 2915 2533 2927 2567
rect 2869 2527 2927 2533
rect 21545 2567 21603 2573
rect 21545 2533 21557 2567
rect 21591 2564 21603 2567
rect 23937 2567 23995 2573
rect 21591 2536 23888 2564
rect 21591 2533 21603 2536
rect 21545 2527 21603 2533
rect 1578 2456 1584 2508
rect 1636 2456 1642 2508
rect 5813 2499 5871 2505
rect 5813 2465 5825 2499
rect 5859 2496 5871 2499
rect 7834 2496 7840 2508
rect 5859 2468 7840 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 7834 2456 7840 2468
rect 7892 2456 7898 2508
rect 8389 2499 8447 2505
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 9950 2496 9956 2508
rect 8435 2468 9956 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 10873 2499 10931 2505
rect 10873 2465 10885 2499
rect 10919 2496 10931 2499
rect 10919 2468 11560 2496
rect 10919 2465 10931 2468
rect 10873 2459 10931 2465
rect 2590 2388 2596 2440
rect 2648 2388 2654 2440
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 842 2320 848 2372
rect 900 2360 906 2372
rect 3160 2360 3188 2391
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 6089 2431 6147 2437
rect 6089 2397 6101 2431
rect 6135 2428 6147 2431
rect 8110 2428 8116 2440
rect 6135 2400 8116 2428
rect 6135 2397 6147 2400
rect 6089 2391 6147 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 8711 2400 9229 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 9766 2388 9772 2440
rect 9824 2388 9830 2440
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2397 11391 2431
rect 11532 2428 11560 2468
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11664 2468 11805 2496
rect 11664 2456 11670 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 13262 2456 13268 2508
rect 13320 2456 13326 2508
rect 14642 2456 14648 2508
rect 14700 2496 14706 2508
rect 14921 2499 14979 2505
rect 14921 2496 14933 2499
rect 14700 2468 14933 2496
rect 14700 2456 14706 2468
rect 14921 2465 14933 2468
rect 14967 2465 14979 2499
rect 14921 2459 14979 2465
rect 16022 2456 16028 2508
rect 16080 2456 16086 2508
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2496 16819 2499
rect 16942 2496 16948 2508
rect 16807 2468 16948 2496
rect 16807 2465 16819 2468
rect 16761 2459 16819 2465
rect 16942 2456 16948 2468
rect 17000 2456 17006 2508
rect 17954 2456 17960 2508
rect 18012 2496 18018 2508
rect 18141 2499 18199 2505
rect 18141 2496 18153 2499
rect 18012 2468 18153 2496
rect 18012 2456 18018 2468
rect 18141 2465 18153 2468
rect 18187 2465 18199 2499
rect 18141 2459 18199 2465
rect 19702 2456 19708 2508
rect 19760 2456 19766 2508
rect 21637 2499 21695 2505
rect 21637 2465 21649 2499
rect 21683 2465 21695 2499
rect 21637 2459 21695 2465
rect 11882 2428 11888 2440
rect 11532 2400 11888 2428
rect 11333 2391 11391 2397
rect 900 2332 3188 2360
rect 11348 2360 11376 2391
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2428 16543 2431
rect 17034 2428 17040 2440
rect 16531 2400 17040 2428
rect 16531 2397 16543 2400
rect 16485 2391 16543 2397
rect 17034 2388 17040 2400
rect 17092 2388 17098 2440
rect 17678 2388 17684 2440
rect 17736 2388 17742 2440
rect 19334 2388 19340 2440
rect 19392 2388 19398 2440
rect 12636 2360 12664 2388
rect 11348 2332 12664 2360
rect 21085 2363 21143 2369
rect 900 2320 906 2332
rect 21085 2329 21097 2363
rect 21131 2360 21143 2363
rect 21177 2363 21235 2369
rect 21177 2360 21189 2363
rect 21131 2332 21189 2360
rect 21131 2329 21143 2332
rect 21085 2323 21143 2329
rect 21177 2329 21189 2332
rect 21223 2329 21235 2363
rect 21652 2360 21680 2459
rect 22002 2456 22008 2508
rect 22060 2496 22066 2508
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 22060 2468 22293 2496
rect 22060 2456 22066 2468
rect 22281 2465 22293 2468
rect 22327 2465 22339 2499
rect 22281 2459 22339 2465
rect 23290 2456 23296 2508
rect 23348 2456 23354 2508
rect 23860 2440 23888 2536
rect 23937 2533 23949 2567
rect 23983 2564 23995 2567
rect 24946 2564 24952 2576
rect 23983 2536 24952 2564
rect 23983 2533 23995 2536
rect 23937 2527 23995 2533
rect 24946 2524 24952 2536
rect 25004 2524 25010 2576
rect 25314 2524 25320 2576
rect 25372 2564 25378 2576
rect 25501 2567 25559 2573
rect 25501 2564 25513 2567
rect 25372 2536 25513 2564
rect 25372 2524 25378 2536
rect 25501 2533 25513 2536
rect 25547 2564 25559 2567
rect 26326 2564 26332 2576
rect 25547 2536 26332 2564
rect 25547 2533 25559 2536
rect 25501 2527 25559 2533
rect 26326 2524 26332 2536
rect 26384 2524 26390 2576
rect 26418 2524 26424 2576
rect 26476 2524 26482 2576
rect 27614 2524 27620 2576
rect 27672 2524 27678 2576
rect 28077 2567 28135 2573
rect 28077 2533 28089 2567
rect 28123 2564 28135 2567
rect 28350 2564 28356 2576
rect 28123 2536 28356 2564
rect 28123 2533 28135 2536
rect 28077 2527 28135 2533
rect 28350 2524 28356 2536
rect 28408 2564 28414 2576
rect 30561 2567 30619 2573
rect 30561 2564 30573 2567
rect 28408 2536 30573 2564
rect 28408 2524 28414 2536
rect 30561 2533 30573 2536
rect 30607 2533 30619 2567
rect 30561 2527 30619 2533
rect 25041 2499 25099 2505
rect 25041 2465 25053 2499
rect 25087 2496 25099 2499
rect 26436 2496 26464 2524
rect 25087 2468 26464 2496
rect 25087 2465 25099 2468
rect 25041 2459 25099 2465
rect 26878 2456 26884 2508
rect 26936 2496 26942 2508
rect 27341 2499 27399 2505
rect 27341 2496 27353 2499
rect 26936 2468 27353 2496
rect 26936 2456 26942 2468
rect 27341 2465 27353 2468
rect 27387 2465 27399 2499
rect 27341 2459 27399 2465
rect 27522 2456 27528 2508
rect 27580 2456 27586 2508
rect 27632 2496 27660 2524
rect 27632 2468 29684 2496
rect 21910 2388 21916 2440
rect 21968 2388 21974 2440
rect 23842 2388 23848 2440
rect 23900 2388 23906 2440
rect 24210 2388 24216 2440
rect 24268 2428 24274 2440
rect 24489 2431 24547 2437
rect 24489 2428 24501 2431
rect 24268 2400 24501 2428
rect 24268 2388 24274 2400
rect 24489 2397 24501 2400
rect 24535 2397 24547 2431
rect 24489 2391 24547 2397
rect 24670 2388 24676 2440
rect 24728 2428 24734 2440
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 24728 2400 25881 2428
rect 24728 2388 24734 2400
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26050 2388 26056 2440
rect 26108 2428 26114 2440
rect 26421 2431 26479 2437
rect 26421 2428 26433 2431
rect 26108 2400 26433 2428
rect 26108 2388 26114 2400
rect 26421 2397 26433 2400
rect 26467 2397 26479 2431
rect 26421 2391 26479 2397
rect 26602 2388 26608 2440
rect 26660 2428 26666 2440
rect 27065 2431 27123 2437
rect 27065 2428 27077 2431
rect 26660 2400 27077 2428
rect 26660 2388 26666 2400
rect 27065 2397 27077 2400
rect 27111 2397 27123 2431
rect 27540 2428 27568 2456
rect 29656 2437 29684 2468
rect 30006 2456 30012 2508
rect 30064 2456 30070 2508
rect 32585 2499 32643 2505
rect 32585 2496 32597 2499
rect 30346 2468 32597 2496
rect 28997 2431 29055 2437
rect 28997 2428 29009 2431
rect 27540 2400 29009 2428
rect 27065 2391 27123 2397
rect 28997 2397 29009 2400
rect 29043 2397 29055 2431
rect 28997 2391 29055 2397
rect 29641 2431 29699 2437
rect 29641 2397 29653 2431
rect 29687 2397 29699 2431
rect 29641 2391 29699 2397
rect 26786 2360 26792 2372
rect 21652 2332 26792 2360
rect 21177 2323 21235 2329
rect 21192 2292 21220 2323
rect 26786 2320 26792 2332
rect 26844 2320 26850 2372
rect 27154 2320 27160 2372
rect 27212 2360 27218 2372
rect 28445 2363 28503 2369
rect 28445 2360 28457 2363
rect 27212 2332 28457 2360
rect 27212 2320 27218 2332
rect 28445 2329 28457 2332
rect 28491 2329 28503 2363
rect 28445 2323 28503 2329
rect 28534 2320 28540 2372
rect 28592 2360 28598 2372
rect 30346 2360 30374 2468
rect 32585 2465 32597 2468
rect 32631 2465 32643 2499
rect 32585 2459 32643 2465
rect 30466 2388 30472 2440
rect 30524 2428 30530 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30524 2400 31033 2428
rect 30524 2388 30530 2400
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 31110 2388 31116 2440
rect 31168 2428 31174 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31168 2400 32137 2428
rect 31168 2388 31174 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 28592 2332 30374 2360
rect 28592 2320 28598 2332
rect 23382 2292 23388 2304
rect 21192 2264 23388 2292
rect 23382 2252 23388 2264
rect 23440 2252 23446 2304
rect 28902 2252 28908 2304
rect 28960 2292 28966 2304
rect 32582 2292 32588 2304
rect 28960 2264 32588 2292
rect 28960 2252 28966 2264
rect 32582 2252 32588 2264
rect 32640 2252 32646 2304
rect 1104 2202 34016 2224
rect 1104 2150 9138 2202
rect 9190 2150 9202 2202
rect 9254 2150 9266 2202
rect 9318 2150 9330 2202
rect 9382 2150 9394 2202
rect 9446 2150 17326 2202
rect 17378 2150 17390 2202
rect 17442 2150 17454 2202
rect 17506 2150 17518 2202
rect 17570 2150 17582 2202
rect 17634 2150 25514 2202
rect 25566 2150 25578 2202
rect 25630 2150 25642 2202
rect 25694 2150 25706 2202
rect 25758 2150 25770 2202
rect 25822 2150 33702 2202
rect 33754 2150 33766 2202
rect 33818 2150 33830 2202
rect 33882 2150 33894 2202
rect 33946 2150 33958 2202
rect 34010 2150 34016 2202
rect 1104 2128 34016 2150
rect 23842 2048 23848 2100
rect 23900 2088 23906 2100
rect 28074 2088 28080 2100
rect 23900 2060 28080 2088
rect 23900 2048 23906 2060
rect 28074 2048 28080 2060
rect 28132 2048 28138 2100
rect 27062 1504 27068 1556
rect 27120 1544 27126 1556
rect 30190 1544 30196 1556
rect 27120 1516 30196 1544
rect 27120 1504 27126 1516
rect 30190 1504 30196 1516
rect 30248 1504 30254 1556
rect 25682 1436 25688 1488
rect 25740 1476 25746 1488
rect 28626 1476 28632 1488
rect 25740 1448 28632 1476
rect 25740 1436 25746 1448
rect 28626 1436 28632 1448
rect 28684 1436 28690 1488
rect 20346 1368 20352 1420
rect 20404 1408 20410 1420
rect 22002 1408 22008 1420
rect 20404 1380 22008 1408
rect 20404 1368 20410 1380
rect 22002 1368 22008 1380
rect 22060 1368 22066 1420
<< via1 >>
rect 9138 32614 9190 32666
rect 9202 32614 9254 32666
rect 9266 32614 9318 32666
rect 9330 32614 9382 32666
rect 9394 32614 9446 32666
rect 17326 32614 17378 32666
rect 17390 32614 17442 32666
rect 17454 32614 17506 32666
rect 17518 32614 17570 32666
rect 17582 32614 17634 32666
rect 25514 32614 25566 32666
rect 25578 32614 25630 32666
rect 25642 32614 25694 32666
rect 25706 32614 25758 32666
rect 25770 32614 25822 32666
rect 33702 32614 33754 32666
rect 33766 32614 33818 32666
rect 33830 32614 33882 32666
rect 33894 32614 33946 32666
rect 33958 32614 34010 32666
rect 5724 32444 5776 32496
rect 2872 32419 2924 32428
rect 2872 32385 2881 32419
rect 2881 32385 2915 32419
rect 2915 32385 2924 32419
rect 2872 32376 2924 32385
rect 7012 32444 7064 32496
rect 10416 32487 10468 32496
rect 10416 32453 10425 32487
rect 10425 32453 10459 32487
rect 10459 32453 10468 32487
rect 10416 32444 10468 32453
rect 15200 32444 15252 32496
rect 21364 32444 21416 32496
rect 1584 32351 1636 32360
rect 1584 32317 1593 32351
rect 1593 32317 1627 32351
rect 1627 32317 1636 32351
rect 1584 32308 1636 32317
rect 8668 32419 8720 32428
rect 8668 32385 8677 32419
rect 8677 32385 8711 32419
rect 8711 32385 8720 32419
rect 8668 32376 8720 32385
rect 11152 32419 11204 32428
rect 11152 32385 11161 32419
rect 11161 32385 11195 32419
rect 11195 32385 11204 32419
rect 11152 32376 11204 32385
rect 13544 32376 13596 32428
rect 14280 32376 14332 32428
rect 6736 32351 6788 32360
rect 6736 32317 6745 32351
rect 6745 32317 6779 32351
rect 6779 32317 6788 32351
rect 6736 32308 6788 32317
rect 8392 32351 8444 32360
rect 8392 32317 8401 32351
rect 8401 32317 8435 32351
rect 8435 32317 8444 32351
rect 8392 32308 8444 32317
rect 9864 32351 9916 32360
rect 9864 32317 9873 32351
rect 9873 32317 9907 32351
rect 9907 32317 9916 32351
rect 9864 32308 9916 32317
rect 12532 32308 12584 32360
rect 14464 32351 14516 32360
rect 14464 32317 14473 32351
rect 14473 32317 14507 32351
rect 14507 32317 14516 32351
rect 14464 32308 14516 32317
rect 15292 32419 15344 32428
rect 15292 32385 15301 32419
rect 15301 32385 15335 32419
rect 15335 32385 15344 32419
rect 15292 32376 15344 32385
rect 17132 32376 17184 32428
rect 21824 32419 21876 32428
rect 21824 32385 21833 32419
rect 21833 32385 21867 32419
rect 21867 32385 21876 32419
rect 21824 32376 21876 32385
rect 17684 32308 17736 32360
rect 18512 32308 18564 32360
rect 20904 32308 20956 32360
rect 22008 32308 22060 32360
rect 9404 32240 9456 32292
rect 12900 32240 12952 32292
rect 20168 32240 20220 32292
rect 29184 32444 29236 32496
rect 24400 32419 24452 32428
rect 24400 32385 24409 32419
rect 24409 32385 24443 32419
rect 24443 32385 24452 32419
rect 24400 32376 24452 32385
rect 25044 32376 25096 32428
rect 26056 32308 26108 32360
rect 26424 32351 26476 32360
rect 26424 32317 26433 32351
rect 26433 32317 26467 32351
rect 26467 32317 26476 32351
rect 26424 32308 26476 32317
rect 26976 32419 27028 32428
rect 26976 32385 26985 32419
rect 26985 32385 27019 32419
rect 27019 32385 27028 32419
rect 26976 32376 27028 32385
rect 28172 32376 28224 32428
rect 29000 32351 29052 32360
rect 29000 32317 29009 32351
rect 29009 32317 29043 32351
rect 29043 32317 29052 32351
rect 29000 32308 29052 32317
rect 30380 32308 30432 32360
rect 32128 32419 32180 32428
rect 32128 32385 32137 32419
rect 32137 32385 32171 32419
rect 32171 32385 32180 32419
rect 32128 32376 32180 32385
rect 2136 32215 2188 32224
rect 2136 32181 2145 32215
rect 2145 32181 2179 32215
rect 2179 32181 2188 32215
rect 2136 32172 2188 32181
rect 4344 32172 4396 32224
rect 6276 32172 6328 32224
rect 6552 32172 6604 32224
rect 8300 32172 8352 32224
rect 13636 32172 13688 32224
rect 16120 32172 16172 32224
rect 16856 32215 16908 32224
rect 16856 32181 16865 32215
rect 16865 32181 16899 32215
rect 16899 32181 16908 32215
rect 16856 32172 16908 32181
rect 18512 32172 18564 32224
rect 26148 32172 26200 32224
rect 26884 32172 26936 32224
rect 31024 32215 31076 32224
rect 31024 32181 31033 32215
rect 31033 32181 31067 32215
rect 31067 32181 31076 32215
rect 31024 32172 31076 32181
rect 5044 32070 5096 32122
rect 5108 32070 5160 32122
rect 5172 32070 5224 32122
rect 5236 32070 5288 32122
rect 5300 32070 5352 32122
rect 13232 32070 13284 32122
rect 13296 32070 13348 32122
rect 13360 32070 13412 32122
rect 13424 32070 13476 32122
rect 13488 32070 13540 32122
rect 21420 32070 21472 32122
rect 21484 32070 21536 32122
rect 21548 32070 21600 32122
rect 21612 32070 21664 32122
rect 21676 32070 21728 32122
rect 29608 32070 29660 32122
rect 29672 32070 29724 32122
rect 29736 32070 29788 32122
rect 29800 32070 29852 32122
rect 29864 32070 29916 32122
rect 2136 31968 2188 32020
rect 2872 31968 2924 32020
rect 6736 31968 6788 32020
rect 4160 31832 4212 31884
rect 6552 31875 6604 31884
rect 6552 31841 6561 31875
rect 6561 31841 6595 31875
rect 6595 31841 6604 31875
rect 6552 31832 6604 31841
rect 7288 31832 7340 31884
rect 9404 31968 9456 32020
rect 11152 31968 11204 32020
rect 15292 31968 15344 32020
rect 16856 31968 16908 32020
rect 21824 31968 21876 32020
rect 24400 31968 24452 32020
rect 27620 31968 27672 32020
rect 11060 31900 11112 31952
rect 9680 31832 9732 31884
rect 1400 31764 1452 31816
rect 2596 31807 2648 31816
rect 2596 31773 2605 31807
rect 2605 31773 2639 31807
rect 2639 31773 2648 31807
rect 2596 31764 2648 31773
rect 4344 31807 4396 31816
rect 4344 31773 4353 31807
rect 4353 31773 4387 31807
rect 4387 31773 4396 31807
rect 4344 31764 4396 31773
rect 6184 31764 6236 31816
rect 7104 31807 7156 31816
rect 7104 31773 7113 31807
rect 7113 31773 7147 31807
rect 7147 31773 7156 31807
rect 7104 31764 7156 31773
rect 7472 31807 7524 31816
rect 7472 31773 7481 31807
rect 7481 31773 7515 31807
rect 7515 31773 7524 31807
rect 7472 31764 7524 31773
rect 10968 31764 11020 31816
rect 12348 31807 12400 31816
rect 12348 31773 12357 31807
rect 12357 31773 12391 31807
rect 12391 31773 12400 31807
rect 12348 31764 12400 31773
rect 11980 31696 12032 31748
rect 14556 31764 14608 31816
rect 18512 31875 18564 31884
rect 18512 31841 18521 31875
rect 18521 31841 18555 31875
rect 18555 31841 18564 31875
rect 18512 31832 18564 31841
rect 26976 31832 27028 31884
rect 28172 31875 28224 31884
rect 28172 31841 28181 31875
rect 28181 31841 28215 31875
rect 28215 31841 28224 31875
rect 28172 31832 28224 31841
rect 32128 31832 32180 31884
rect 17224 31739 17276 31748
rect 17224 31705 17233 31739
rect 17233 31705 17267 31739
rect 17267 31705 17276 31739
rect 17224 31696 17276 31705
rect 22376 31764 22428 31816
rect 23388 31764 23440 31816
rect 24676 31807 24728 31816
rect 24676 31773 24685 31807
rect 24685 31773 24719 31807
rect 24719 31773 24728 31807
rect 24676 31764 24728 31773
rect 26148 31807 26200 31816
rect 26148 31773 26157 31807
rect 26157 31773 26191 31807
rect 26191 31773 26200 31807
rect 26148 31764 26200 31773
rect 27620 31807 27672 31816
rect 27620 31773 27629 31807
rect 27629 31773 27663 31807
rect 27663 31773 27672 31807
rect 27620 31764 27672 31773
rect 29092 31764 29144 31816
rect 33048 31807 33100 31816
rect 33048 31773 33057 31807
rect 33057 31773 33091 31807
rect 33091 31773 33100 31807
rect 33048 31764 33100 31773
rect 26516 31739 26568 31748
rect 26516 31705 26525 31739
rect 26525 31705 26559 31739
rect 26559 31705 26568 31739
rect 26516 31696 26568 31705
rect 3792 31671 3844 31680
rect 3792 31637 3801 31671
rect 3801 31637 3835 31671
rect 3835 31637 3844 31671
rect 3792 31628 3844 31637
rect 8944 31628 8996 31680
rect 18144 31671 18196 31680
rect 18144 31637 18153 31671
rect 18153 31637 18187 31671
rect 18187 31637 18196 31671
rect 18144 31628 18196 31637
rect 20260 31628 20312 31680
rect 21272 31671 21324 31680
rect 21272 31637 21281 31671
rect 21281 31637 21315 31671
rect 21315 31637 21324 31671
rect 21272 31628 21324 31637
rect 25412 31628 25464 31680
rect 27160 31671 27212 31680
rect 27160 31637 27169 31671
rect 27169 31637 27203 31671
rect 27203 31637 27212 31671
rect 27160 31628 27212 31637
rect 28540 31671 28592 31680
rect 28540 31637 28549 31671
rect 28549 31637 28583 31671
rect 28583 31637 28592 31671
rect 28540 31628 28592 31637
rect 30196 31628 30248 31680
rect 31852 31628 31904 31680
rect 9138 31526 9190 31578
rect 9202 31526 9254 31578
rect 9266 31526 9318 31578
rect 9330 31526 9382 31578
rect 9394 31526 9446 31578
rect 17326 31526 17378 31578
rect 17390 31526 17442 31578
rect 17454 31526 17506 31578
rect 17518 31526 17570 31578
rect 17582 31526 17634 31578
rect 25514 31526 25566 31578
rect 25578 31526 25630 31578
rect 25642 31526 25694 31578
rect 25706 31526 25758 31578
rect 25770 31526 25822 31578
rect 33702 31526 33754 31578
rect 33766 31526 33818 31578
rect 33830 31526 33882 31578
rect 33894 31526 33946 31578
rect 33958 31526 34010 31578
rect 1584 31424 1636 31476
rect 1768 31220 1820 31272
rect 3792 31356 3844 31408
rect 6000 31356 6052 31408
rect 6184 31399 6236 31408
rect 6184 31365 6193 31399
rect 6193 31365 6227 31399
rect 6227 31365 6236 31399
rect 6184 31356 6236 31365
rect 12532 31424 12584 31476
rect 14464 31424 14516 31476
rect 6828 31288 6880 31340
rect 10140 31288 10192 31340
rect 12992 31288 13044 31340
rect 14464 31288 14516 31340
rect 16304 31288 16356 31340
rect 17960 31288 18012 31340
rect 18144 31288 18196 31340
rect 5448 31084 5500 31136
rect 8944 31220 8996 31272
rect 11336 31263 11388 31272
rect 11336 31229 11345 31263
rect 11345 31229 11379 31263
rect 11379 31229 11388 31263
rect 11336 31220 11388 31229
rect 13084 31263 13136 31272
rect 13084 31229 13093 31263
rect 13093 31229 13127 31263
rect 13127 31229 13136 31263
rect 13084 31220 13136 31229
rect 18696 31263 18748 31272
rect 18696 31229 18705 31263
rect 18705 31229 18739 31263
rect 18739 31229 18748 31263
rect 18696 31220 18748 31229
rect 20260 31331 20312 31340
rect 20260 31297 20269 31331
rect 20269 31297 20303 31331
rect 20303 31297 20312 31331
rect 20260 31288 20312 31297
rect 23388 31424 23440 31476
rect 29000 31424 29052 31476
rect 6276 31152 6328 31204
rect 8300 31152 8352 31204
rect 22928 31288 22980 31340
rect 23388 31288 23440 31340
rect 24952 31288 25004 31340
rect 25412 31288 25464 31340
rect 26332 31288 26384 31340
rect 28264 31288 28316 31340
rect 30932 31356 30984 31408
rect 28448 31288 28500 31340
rect 29092 31331 29144 31340
rect 29092 31297 29101 31331
rect 29101 31297 29135 31331
rect 29135 31297 29144 31331
rect 29092 31288 29144 31297
rect 29276 31288 29328 31340
rect 31852 31399 31904 31408
rect 31852 31365 31861 31399
rect 31861 31365 31895 31399
rect 31895 31365 31904 31399
rect 31852 31356 31904 31365
rect 31576 31288 31628 31340
rect 21272 31220 21324 31272
rect 21916 31220 21968 31272
rect 31852 31220 31904 31272
rect 31484 31195 31536 31204
rect 31484 31161 31493 31195
rect 31493 31161 31527 31195
rect 31527 31161 31536 31195
rect 31484 31152 31536 31161
rect 5724 31127 5776 31136
rect 5724 31093 5733 31127
rect 5733 31093 5767 31127
rect 5767 31093 5776 31127
rect 5724 31084 5776 31093
rect 7840 31084 7892 31136
rect 10416 31084 10468 31136
rect 10692 31127 10744 31136
rect 10692 31093 10701 31127
rect 10701 31093 10735 31127
rect 10735 31093 10744 31127
rect 10692 31084 10744 31093
rect 12440 31084 12492 31136
rect 16672 31127 16724 31136
rect 16672 31093 16681 31127
rect 16681 31093 16715 31127
rect 16715 31093 16724 31127
rect 16672 31084 16724 31093
rect 17684 31084 17736 31136
rect 18880 31127 18932 31136
rect 18880 31093 18889 31127
rect 18889 31093 18923 31127
rect 18923 31093 18932 31127
rect 18880 31084 18932 31093
rect 22100 31127 22152 31136
rect 22100 31093 22109 31127
rect 22109 31093 22143 31127
rect 22143 31093 22152 31127
rect 22100 31084 22152 31093
rect 23664 31127 23716 31136
rect 23664 31093 23673 31127
rect 23673 31093 23707 31127
rect 23707 31093 23716 31127
rect 23664 31084 23716 31093
rect 26976 31127 27028 31136
rect 26976 31093 26985 31127
rect 26985 31093 27019 31127
rect 27019 31093 27028 31127
rect 26976 31084 27028 31093
rect 29092 31084 29144 31136
rect 32128 31084 32180 31136
rect 5044 30982 5096 31034
rect 5108 30982 5160 31034
rect 5172 30982 5224 31034
rect 5236 30982 5288 31034
rect 5300 30982 5352 31034
rect 13232 30982 13284 31034
rect 13296 30982 13348 31034
rect 13360 30982 13412 31034
rect 13424 30982 13476 31034
rect 13488 30982 13540 31034
rect 21420 30982 21472 31034
rect 21484 30982 21536 31034
rect 21548 30982 21600 31034
rect 21612 30982 21664 31034
rect 21676 30982 21728 31034
rect 29608 30982 29660 31034
rect 29672 30982 29724 31034
rect 29736 30982 29788 31034
rect 29800 30982 29852 31034
rect 29864 30982 29916 31034
rect 12348 30923 12400 30932
rect 12348 30889 12357 30923
rect 12357 30889 12391 30923
rect 12391 30889 12400 30923
rect 12348 30880 12400 30889
rect 16672 30880 16724 30932
rect 18696 30880 18748 30932
rect 18880 30880 18932 30932
rect 20260 30880 20312 30932
rect 21916 30923 21968 30932
rect 21916 30889 21925 30923
rect 21925 30889 21959 30923
rect 21959 30889 21968 30923
rect 21916 30880 21968 30889
rect 22100 30880 22152 30932
rect 14556 30812 14608 30864
rect 1768 30719 1820 30728
rect 1768 30685 1777 30719
rect 1777 30685 1811 30719
rect 1811 30685 1820 30719
rect 5448 30744 5500 30796
rect 7472 30787 7524 30796
rect 7472 30753 7481 30787
rect 7481 30753 7515 30787
rect 7515 30753 7524 30787
rect 7472 30744 7524 30753
rect 8852 30744 8904 30796
rect 16120 30787 16172 30796
rect 16120 30753 16129 30787
rect 16129 30753 16163 30787
rect 16163 30753 16172 30787
rect 16120 30744 16172 30753
rect 17040 30744 17092 30796
rect 23664 30880 23716 30932
rect 24952 30880 25004 30932
rect 26424 30880 26476 30932
rect 26240 30812 26292 30864
rect 33048 30880 33100 30932
rect 1768 30676 1820 30685
rect 5632 30676 5684 30728
rect 4160 30608 4212 30660
rect 5540 30608 5592 30660
rect 5724 30608 5776 30660
rect 8024 30719 8076 30728
rect 8024 30685 8033 30719
rect 8033 30685 8067 30719
rect 8067 30685 8076 30719
rect 8024 30676 8076 30685
rect 8392 30676 8444 30728
rect 11060 30676 11112 30728
rect 12900 30719 12952 30728
rect 12900 30685 12909 30719
rect 12909 30685 12943 30719
rect 12943 30685 12952 30719
rect 12900 30676 12952 30685
rect 13084 30676 13136 30728
rect 13728 30676 13780 30728
rect 14280 30676 14332 30728
rect 17224 30719 17276 30728
rect 17224 30685 17233 30719
rect 17233 30685 17267 30719
rect 17267 30685 17276 30719
rect 17224 30676 17276 30685
rect 20904 30676 20956 30728
rect 27436 30787 27488 30796
rect 27436 30753 27445 30787
rect 27445 30753 27479 30787
rect 27479 30753 27488 30787
rect 27436 30744 27488 30753
rect 26516 30676 26568 30728
rect 30932 30787 30984 30796
rect 30932 30753 30941 30787
rect 30941 30753 30975 30787
rect 30975 30753 30984 30787
rect 30932 30744 30984 30753
rect 31392 30744 31444 30796
rect 28080 30719 28132 30728
rect 28080 30685 28089 30719
rect 28089 30685 28123 30719
rect 28123 30685 28132 30719
rect 28080 30676 28132 30685
rect 21180 30608 21232 30660
rect 23296 30608 23348 30660
rect 25320 30608 25372 30660
rect 27160 30608 27212 30660
rect 27436 30608 27488 30660
rect 28908 30608 28960 30660
rect 32036 30608 32088 30660
rect 32128 30651 32180 30660
rect 32128 30617 32146 30651
rect 32146 30617 32180 30651
rect 32128 30608 32180 30617
rect 4620 30540 4672 30592
rect 6920 30583 6972 30592
rect 6920 30549 6929 30583
rect 6929 30549 6963 30583
rect 6963 30549 6972 30583
rect 6920 30540 6972 30549
rect 8944 30540 8996 30592
rect 10876 30583 10928 30592
rect 10876 30549 10885 30583
rect 10885 30549 10919 30583
rect 10919 30549 10928 30583
rect 10876 30540 10928 30549
rect 25412 30540 25464 30592
rect 26700 30540 26752 30592
rect 30472 30540 30524 30592
rect 31116 30540 31168 30592
rect 9138 30438 9190 30490
rect 9202 30438 9254 30490
rect 9266 30438 9318 30490
rect 9330 30438 9382 30490
rect 9394 30438 9446 30490
rect 17326 30438 17378 30490
rect 17390 30438 17442 30490
rect 17454 30438 17506 30490
rect 17518 30438 17570 30490
rect 17582 30438 17634 30490
rect 25514 30438 25566 30490
rect 25578 30438 25630 30490
rect 25642 30438 25694 30490
rect 25706 30438 25758 30490
rect 25770 30438 25822 30490
rect 33702 30438 33754 30490
rect 33766 30438 33818 30490
rect 33830 30438 33882 30490
rect 33894 30438 33946 30490
rect 33958 30438 34010 30490
rect 2504 30336 2556 30388
rect 2596 30268 2648 30320
rect 6828 30379 6880 30388
rect 6828 30345 6837 30379
rect 6837 30345 6871 30379
rect 6871 30345 6880 30379
rect 6828 30336 6880 30345
rect 8300 30336 8352 30388
rect 11336 30379 11388 30388
rect 11336 30345 11345 30379
rect 11345 30345 11379 30379
rect 11379 30345 11388 30379
rect 11336 30336 11388 30345
rect 12992 30336 13044 30388
rect 13728 30379 13780 30388
rect 13728 30345 13737 30379
rect 13737 30345 13771 30379
rect 13771 30345 13780 30379
rect 13728 30336 13780 30345
rect 14464 30379 14516 30388
rect 14464 30345 14473 30379
rect 14473 30345 14507 30379
rect 14507 30345 14516 30379
rect 14464 30336 14516 30345
rect 16304 30379 16356 30388
rect 16304 30345 16313 30379
rect 16313 30345 16347 30379
rect 16347 30345 16356 30379
rect 16304 30336 16356 30345
rect 17960 30336 18012 30388
rect 21180 30379 21232 30388
rect 21180 30345 21189 30379
rect 21189 30345 21223 30379
rect 21223 30345 21232 30379
rect 21180 30336 21232 30345
rect 22468 30379 22520 30388
rect 22468 30345 22477 30379
rect 22477 30345 22511 30379
rect 22511 30345 22520 30379
rect 22468 30336 22520 30345
rect 23388 30336 23440 30388
rect 27620 30336 27672 30388
rect 28172 30336 28224 30388
rect 2964 30200 3016 30252
rect 1032 30132 1084 30184
rect 6184 30268 6236 30320
rect 6368 30311 6420 30320
rect 6368 30277 6377 30311
rect 6377 30277 6411 30311
rect 6411 30277 6420 30311
rect 6368 30268 6420 30277
rect 5540 30243 5592 30252
rect 5540 30209 5549 30243
rect 5549 30209 5583 30243
rect 5583 30209 5592 30243
rect 5540 30200 5592 30209
rect 6920 30200 6972 30252
rect 8668 30268 8720 30320
rect 9864 30268 9916 30320
rect 24676 30268 24728 30320
rect 10416 30243 10468 30252
rect 10416 30209 10425 30243
rect 10425 30209 10459 30243
rect 10459 30209 10468 30243
rect 10416 30200 10468 30209
rect 10876 30200 10928 30252
rect 12440 30243 12492 30252
rect 12440 30209 12449 30243
rect 12449 30209 12483 30243
rect 12483 30209 12492 30243
rect 12440 30200 12492 30209
rect 11152 30132 11204 30184
rect 21272 30200 21324 30252
rect 9680 30064 9732 30116
rect 13728 30064 13780 30116
rect 4528 29996 4580 30048
rect 6644 29996 6696 30048
rect 13636 29996 13688 30048
rect 14556 30107 14608 30116
rect 14556 30073 14565 30107
rect 14565 30073 14599 30107
rect 14599 30073 14608 30107
rect 14556 30064 14608 30073
rect 22008 30132 22060 30184
rect 25412 30243 25464 30252
rect 25412 30209 25421 30243
rect 25421 30209 25455 30243
rect 25455 30209 25464 30243
rect 25412 30200 25464 30209
rect 23572 30175 23624 30184
rect 23572 30141 23581 30175
rect 23581 30141 23615 30175
rect 23615 30141 23624 30175
rect 23572 30132 23624 30141
rect 17684 30064 17736 30116
rect 18512 30064 18564 30116
rect 22928 30107 22980 30116
rect 22928 30073 22937 30107
rect 22937 30073 22971 30107
rect 22971 30073 22980 30107
rect 22928 30064 22980 30073
rect 26240 30132 26292 30184
rect 26332 30132 26384 30184
rect 27436 30175 27488 30184
rect 27436 30141 27445 30175
rect 27445 30141 27479 30175
rect 27479 30141 27488 30175
rect 27436 30132 27488 30141
rect 27988 30132 28040 30184
rect 31300 30268 31352 30320
rect 29000 30243 29052 30252
rect 29000 30209 29009 30243
rect 29009 30209 29043 30243
rect 29043 30209 29052 30243
rect 29000 30200 29052 30209
rect 30012 30200 30064 30252
rect 30104 30200 30156 30252
rect 29184 30175 29236 30184
rect 29184 30141 29193 30175
rect 29193 30141 29227 30175
rect 29227 30141 29236 30175
rect 29184 30132 29236 30141
rect 30932 30175 30984 30184
rect 30932 30141 30941 30175
rect 30941 30141 30975 30175
rect 30975 30141 30984 30175
rect 30932 30132 30984 30141
rect 32128 30175 32180 30184
rect 32128 30141 32137 30175
rect 32137 30141 32171 30175
rect 32171 30141 32180 30175
rect 32128 30132 32180 30141
rect 24952 30064 25004 30116
rect 27344 30064 27396 30116
rect 31024 30064 31076 30116
rect 15752 30039 15804 30048
rect 15752 30005 15761 30039
rect 15761 30005 15795 30039
rect 15795 30005 15804 30039
rect 15752 29996 15804 30005
rect 29276 29996 29328 30048
rect 29368 29996 29420 30048
rect 30196 29996 30248 30048
rect 33508 30039 33560 30048
rect 33508 30005 33517 30039
rect 33517 30005 33551 30039
rect 33551 30005 33560 30039
rect 33508 29996 33560 30005
rect 5044 29894 5096 29946
rect 5108 29894 5160 29946
rect 5172 29894 5224 29946
rect 5236 29894 5288 29946
rect 5300 29894 5352 29946
rect 13232 29894 13284 29946
rect 13296 29894 13348 29946
rect 13360 29894 13412 29946
rect 13424 29894 13476 29946
rect 13488 29894 13540 29946
rect 21420 29894 21472 29946
rect 21484 29894 21536 29946
rect 21548 29894 21600 29946
rect 21612 29894 21664 29946
rect 21676 29894 21728 29946
rect 29608 29894 29660 29946
rect 29672 29894 29724 29946
rect 29736 29894 29788 29946
rect 29800 29894 29852 29946
rect 29864 29894 29916 29946
rect 4160 29792 4212 29844
rect 7012 29792 7064 29844
rect 7104 29792 7156 29844
rect 10140 29792 10192 29844
rect 10968 29792 11020 29844
rect 26240 29835 26292 29844
rect 26240 29801 26249 29835
rect 26249 29801 26283 29835
rect 26283 29801 26292 29835
rect 26240 29792 26292 29801
rect 28448 29792 28500 29844
rect 6184 29767 6236 29776
rect 6184 29733 6193 29767
rect 6193 29733 6227 29767
rect 6227 29733 6236 29767
rect 6184 29724 6236 29733
rect 10692 29724 10744 29776
rect 3424 29656 3476 29708
rect 4528 29699 4580 29708
rect 4528 29665 4537 29699
rect 4537 29665 4571 29699
rect 4571 29665 4580 29699
rect 4528 29656 4580 29665
rect 4620 29656 4672 29708
rect 6368 29656 6420 29708
rect 6644 29699 6696 29708
rect 6644 29665 6653 29699
rect 6653 29665 6687 29699
rect 6687 29665 6696 29699
rect 6644 29656 6696 29665
rect 7840 29699 7892 29708
rect 7840 29665 7849 29699
rect 7849 29665 7883 29699
rect 7883 29665 7892 29699
rect 7840 29656 7892 29665
rect 8944 29656 8996 29708
rect 11152 29699 11204 29708
rect 11152 29665 11161 29699
rect 11161 29665 11195 29699
rect 11195 29665 11204 29699
rect 11152 29656 11204 29665
rect 28264 29724 28316 29776
rect 31392 29724 31444 29776
rect 24860 29699 24912 29708
rect 24860 29665 24869 29699
rect 24869 29665 24903 29699
rect 24903 29665 24912 29699
rect 24860 29656 24912 29665
rect 4252 29588 4304 29640
rect 4896 29588 4948 29640
rect 23572 29631 23624 29640
rect 23572 29597 23581 29631
rect 23581 29597 23615 29631
rect 23615 29597 23624 29631
rect 23572 29588 23624 29597
rect 25320 29588 25372 29640
rect 26700 29588 26752 29640
rect 26884 29631 26936 29640
rect 26884 29597 26893 29631
rect 26893 29597 26927 29631
rect 26927 29597 26936 29631
rect 26884 29588 26936 29597
rect 27344 29631 27396 29640
rect 27344 29597 27353 29631
rect 27353 29597 27387 29631
rect 27387 29597 27396 29631
rect 27344 29588 27396 29597
rect 29000 29656 29052 29708
rect 30288 29631 30340 29640
rect 30288 29597 30297 29631
rect 30297 29597 30331 29631
rect 30331 29597 30340 29631
rect 30288 29588 30340 29597
rect 28632 29563 28684 29572
rect 28632 29529 28641 29563
rect 28641 29529 28675 29563
rect 28675 29529 28684 29563
rect 28632 29520 28684 29529
rect 28724 29520 28776 29572
rect 29368 29520 29420 29572
rect 30196 29520 30248 29572
rect 32128 29520 32180 29572
rect 2872 29452 2924 29504
rect 3516 29495 3568 29504
rect 3516 29461 3525 29495
rect 3525 29461 3559 29495
rect 3559 29461 3568 29495
rect 3516 29452 3568 29461
rect 5908 29495 5960 29504
rect 5908 29461 5917 29495
rect 5917 29461 5951 29495
rect 5951 29461 5960 29495
rect 5908 29452 5960 29461
rect 29276 29452 29328 29504
rect 29460 29452 29512 29504
rect 9138 29350 9190 29402
rect 9202 29350 9254 29402
rect 9266 29350 9318 29402
rect 9330 29350 9382 29402
rect 9394 29350 9446 29402
rect 17326 29350 17378 29402
rect 17390 29350 17442 29402
rect 17454 29350 17506 29402
rect 17518 29350 17570 29402
rect 17582 29350 17634 29402
rect 25514 29350 25566 29402
rect 25578 29350 25630 29402
rect 25642 29350 25694 29402
rect 25706 29350 25758 29402
rect 25770 29350 25822 29402
rect 33702 29350 33754 29402
rect 33766 29350 33818 29402
rect 33830 29350 33882 29402
rect 33894 29350 33946 29402
rect 33958 29350 34010 29402
rect 8024 29248 8076 29300
rect 28080 29248 28132 29300
rect 31116 29248 31168 29300
rect 32956 29180 33008 29232
rect 2872 29155 2924 29164
rect 2872 29121 2881 29155
rect 2881 29121 2915 29155
rect 2915 29121 2924 29155
rect 2872 29112 2924 29121
rect 3608 29112 3660 29164
rect 4436 29155 4488 29164
rect 4436 29121 4445 29155
rect 4445 29121 4479 29155
rect 4479 29121 4488 29155
rect 4436 29112 4488 29121
rect 6276 29112 6328 29164
rect 26976 29112 27028 29164
rect 29092 29112 29144 29164
rect 29184 29155 29236 29164
rect 29184 29121 29193 29155
rect 29193 29121 29227 29155
rect 29227 29121 29236 29155
rect 29184 29112 29236 29121
rect 31944 29155 31996 29164
rect 31944 29121 31953 29155
rect 31953 29121 31987 29155
rect 31987 29121 31996 29155
rect 31944 29112 31996 29121
rect 2780 29044 2832 29096
rect 3332 29087 3384 29096
rect 3332 29053 3341 29087
rect 3341 29053 3375 29087
rect 3375 29053 3384 29087
rect 3332 29044 3384 29053
rect 4344 29044 4396 29096
rect 26792 29087 26844 29096
rect 26792 29053 26801 29087
rect 26801 29053 26835 29087
rect 26835 29053 26844 29087
rect 26792 29044 26844 29053
rect 30380 29044 30432 29096
rect 31484 29087 31536 29096
rect 31484 29053 31493 29087
rect 31493 29053 31527 29087
rect 31527 29053 31536 29087
rect 31484 29044 31536 29053
rect 29368 28976 29420 29028
rect 32128 29087 32180 29096
rect 32128 29053 32137 29087
rect 32137 29053 32171 29087
rect 32171 29053 32180 29087
rect 32128 29044 32180 29053
rect 27160 28908 27212 28960
rect 28080 28908 28132 28960
rect 28724 28908 28776 28960
rect 30748 28908 30800 28960
rect 5044 28806 5096 28858
rect 5108 28806 5160 28858
rect 5172 28806 5224 28858
rect 5236 28806 5288 28858
rect 5300 28806 5352 28858
rect 13232 28806 13284 28858
rect 13296 28806 13348 28858
rect 13360 28806 13412 28858
rect 13424 28806 13476 28858
rect 13488 28806 13540 28858
rect 21420 28806 21472 28858
rect 21484 28806 21536 28858
rect 21548 28806 21600 28858
rect 21612 28806 21664 28858
rect 21676 28806 21728 28858
rect 29608 28806 29660 28858
rect 29672 28806 29724 28858
rect 29736 28806 29788 28858
rect 29800 28806 29852 28858
rect 29864 28806 29916 28858
rect 31576 28704 31628 28756
rect 4436 28611 4488 28620
rect 4436 28577 4445 28611
rect 4445 28577 4479 28611
rect 4479 28577 4488 28611
rect 4436 28568 4488 28577
rect 5908 28611 5960 28620
rect 5908 28577 5917 28611
rect 5917 28577 5951 28611
rect 5951 28577 5960 28611
rect 5908 28568 5960 28577
rect 6000 28611 6052 28620
rect 6000 28577 6009 28611
rect 6009 28577 6043 28611
rect 6043 28577 6052 28611
rect 6000 28568 6052 28577
rect 33508 28636 33560 28688
rect 30748 28568 30800 28620
rect 30840 28611 30892 28620
rect 30840 28577 30849 28611
rect 30849 28577 30883 28611
rect 30883 28577 30892 28611
rect 30840 28568 30892 28577
rect 31944 28568 31996 28620
rect 2964 28543 3016 28552
rect 2964 28509 2973 28543
rect 2973 28509 3007 28543
rect 3007 28509 3016 28543
rect 2964 28500 3016 28509
rect 3884 28543 3936 28552
rect 3884 28509 3893 28543
rect 3893 28509 3927 28543
rect 3927 28509 3936 28543
rect 3884 28500 3936 28509
rect 10416 28500 10468 28552
rect 24952 28500 25004 28552
rect 27988 28543 28040 28552
rect 27988 28509 27997 28543
rect 27997 28509 28031 28543
rect 28031 28509 28040 28543
rect 27988 28500 28040 28509
rect 28724 28543 28776 28552
rect 3792 28432 3844 28484
rect 28724 28509 28733 28543
rect 28733 28509 28767 28543
rect 28767 28509 28776 28543
rect 28724 28500 28776 28509
rect 30564 28543 30616 28552
rect 30564 28509 30573 28543
rect 30573 28509 30607 28543
rect 30607 28509 30616 28543
rect 30564 28500 30616 28509
rect 31852 28543 31904 28552
rect 31852 28509 31861 28543
rect 31861 28509 31895 28543
rect 31895 28509 31904 28543
rect 31852 28500 31904 28509
rect 2596 28364 2648 28416
rect 4344 28364 4396 28416
rect 4436 28364 4488 28416
rect 5724 28364 5776 28416
rect 6184 28364 6236 28416
rect 7104 28364 7156 28416
rect 27712 28364 27764 28416
rect 27896 28407 27948 28416
rect 27896 28373 27905 28407
rect 27905 28373 27939 28407
rect 27939 28373 27948 28407
rect 27896 28364 27948 28373
rect 29920 28407 29972 28416
rect 29920 28373 29929 28407
rect 29929 28373 29963 28407
rect 29963 28373 29972 28407
rect 29920 28364 29972 28373
rect 9138 28262 9190 28314
rect 9202 28262 9254 28314
rect 9266 28262 9318 28314
rect 9330 28262 9382 28314
rect 9394 28262 9446 28314
rect 17326 28262 17378 28314
rect 17390 28262 17442 28314
rect 17454 28262 17506 28314
rect 17518 28262 17570 28314
rect 17582 28262 17634 28314
rect 25514 28262 25566 28314
rect 25578 28262 25630 28314
rect 25642 28262 25694 28314
rect 25706 28262 25758 28314
rect 25770 28262 25822 28314
rect 33702 28262 33754 28314
rect 33766 28262 33818 28314
rect 33830 28262 33882 28314
rect 33894 28262 33946 28314
rect 33958 28262 34010 28314
rect 4896 28160 4948 28212
rect 26792 28160 26844 28212
rect 30104 28160 30156 28212
rect 30564 28160 30616 28212
rect 3608 28135 3660 28144
rect 3608 28101 3617 28135
rect 3617 28101 3651 28135
rect 3651 28101 3660 28135
rect 3608 28092 3660 28101
rect 2596 28067 2648 28076
rect 2596 28033 2605 28067
rect 2605 28033 2639 28067
rect 2639 28033 2648 28067
rect 2596 28024 2648 28033
rect 4160 28067 4212 28076
rect 4160 28033 4169 28067
rect 4169 28033 4203 28067
rect 4203 28033 4212 28067
rect 4160 28024 4212 28033
rect 5724 28067 5776 28076
rect 5724 28033 5733 28067
rect 5733 28033 5767 28067
rect 5767 28033 5776 28067
rect 5724 28024 5776 28033
rect 1584 27999 1636 28008
rect 1584 27965 1593 27999
rect 1593 27965 1627 27999
rect 1627 27965 1636 27999
rect 1584 27956 1636 27965
rect 4804 27956 4856 28008
rect 27896 28024 27948 28076
rect 29460 28024 29512 28076
rect 29920 28024 29972 28076
rect 31944 28067 31996 28076
rect 31944 28033 31953 28067
rect 31953 28033 31987 28067
rect 31987 28033 31996 28067
rect 31944 28024 31996 28033
rect 29184 27956 29236 28008
rect 31392 27956 31444 28008
rect 31484 27999 31536 28008
rect 31484 27965 31493 27999
rect 31493 27965 31527 27999
rect 31527 27965 31536 27999
rect 31484 27956 31536 27965
rect 31668 27956 31720 28008
rect 32128 27999 32180 28008
rect 32128 27965 32137 27999
rect 32137 27965 32171 27999
rect 32171 27965 32180 27999
rect 32128 27956 32180 27965
rect 27988 27888 28040 27940
rect 4896 27820 4948 27872
rect 26884 27820 26936 27872
rect 30104 27820 30156 27872
rect 5044 27718 5096 27770
rect 5108 27718 5160 27770
rect 5172 27718 5224 27770
rect 5236 27718 5288 27770
rect 5300 27718 5352 27770
rect 13232 27718 13284 27770
rect 13296 27718 13348 27770
rect 13360 27718 13412 27770
rect 13424 27718 13476 27770
rect 13488 27718 13540 27770
rect 21420 27718 21472 27770
rect 21484 27718 21536 27770
rect 21548 27718 21600 27770
rect 21612 27718 21664 27770
rect 21676 27718 21728 27770
rect 29608 27718 29660 27770
rect 29672 27718 29724 27770
rect 29736 27718 29788 27770
rect 29800 27718 29852 27770
rect 29864 27718 29916 27770
rect 2964 27616 3016 27668
rect 3884 27616 3936 27668
rect 4160 27616 4212 27668
rect 4804 27616 4856 27668
rect 24860 27548 24912 27600
rect 27160 27591 27212 27600
rect 27160 27557 27169 27591
rect 27169 27557 27203 27591
rect 27203 27557 27212 27591
rect 27160 27548 27212 27557
rect 28908 27616 28960 27668
rect 30288 27616 30340 27668
rect 28356 27548 28408 27600
rect 4436 27523 4488 27532
rect 4436 27489 4445 27523
rect 4445 27489 4479 27523
rect 4479 27489 4488 27523
rect 4436 27480 4488 27489
rect 4896 27480 4948 27532
rect 28172 27480 28224 27532
rect 30472 27548 30524 27600
rect 32220 27548 32272 27600
rect 1768 27455 1820 27464
rect 1768 27421 1777 27455
rect 1777 27421 1811 27455
rect 1811 27421 1820 27455
rect 1768 27412 1820 27421
rect 5816 27455 5868 27464
rect 5816 27421 5825 27455
rect 5825 27421 5859 27455
rect 5859 27421 5868 27455
rect 5816 27412 5868 27421
rect 28632 27412 28684 27464
rect 28724 27455 28776 27464
rect 28724 27421 28733 27455
rect 28733 27421 28767 27455
rect 28767 27421 28776 27455
rect 28724 27412 28776 27421
rect 29276 27455 29328 27464
rect 29276 27421 29285 27455
rect 29285 27421 29319 27455
rect 29319 27421 29328 27455
rect 29276 27412 29328 27421
rect 29552 27455 29604 27464
rect 29552 27421 29561 27455
rect 29561 27421 29595 27455
rect 29595 27421 29604 27455
rect 29552 27412 29604 27421
rect 31944 27480 31996 27532
rect 32220 27455 32272 27464
rect 32220 27421 32229 27455
rect 32229 27421 32263 27455
rect 32263 27421 32272 27455
rect 32220 27412 32272 27421
rect 3608 27344 3660 27396
rect 26884 27387 26936 27396
rect 26884 27353 26893 27387
rect 26893 27353 26927 27387
rect 26927 27353 26936 27387
rect 26884 27344 26936 27353
rect 28080 27344 28132 27396
rect 27988 27319 28040 27328
rect 27988 27285 27997 27319
rect 27997 27285 28031 27319
rect 28031 27285 28040 27319
rect 27988 27276 28040 27285
rect 9138 27174 9190 27226
rect 9202 27174 9254 27226
rect 9266 27174 9318 27226
rect 9330 27174 9382 27226
rect 9394 27174 9446 27226
rect 17326 27174 17378 27226
rect 17390 27174 17442 27226
rect 17454 27174 17506 27226
rect 17518 27174 17570 27226
rect 17582 27174 17634 27226
rect 25514 27174 25566 27226
rect 25578 27174 25630 27226
rect 25642 27174 25694 27226
rect 25706 27174 25758 27226
rect 25770 27174 25822 27226
rect 33702 27174 33754 27226
rect 33766 27174 33818 27226
rect 33830 27174 33882 27226
rect 33894 27174 33946 27226
rect 33958 27174 34010 27226
rect 3608 27072 3660 27124
rect 5816 27072 5868 27124
rect 10416 27115 10468 27124
rect 10416 27081 10425 27115
rect 10425 27081 10459 27115
rect 10459 27081 10468 27115
rect 10416 27072 10468 27081
rect 1768 26936 1820 26988
rect 2780 26936 2832 26988
rect 4160 26936 4212 26988
rect 4344 26979 4396 26988
rect 4344 26945 4353 26979
rect 4353 26945 4387 26979
rect 4387 26945 4396 26979
rect 4344 26936 4396 26945
rect 5724 27004 5776 27056
rect 6368 27004 6420 27056
rect 28356 27115 28408 27124
rect 28356 27081 28365 27115
rect 28365 27081 28399 27115
rect 28399 27081 28408 27115
rect 28356 27072 28408 27081
rect 30012 27072 30064 27124
rect 30196 27072 30248 27124
rect 32220 27072 32272 27124
rect 33416 27004 33468 27056
rect 5632 26936 5684 26988
rect 7104 26979 7156 26988
rect 7104 26945 7113 26979
rect 7113 26945 7147 26979
rect 7147 26945 7156 26979
rect 7104 26936 7156 26945
rect 27712 26936 27764 26988
rect 12072 26868 12124 26920
rect 26884 26868 26936 26920
rect 27804 26911 27856 26920
rect 27804 26877 27813 26911
rect 27813 26877 27847 26911
rect 27847 26877 27856 26911
rect 27804 26868 27856 26877
rect 27988 26936 28040 26988
rect 30104 26936 30156 26988
rect 30932 26936 30984 26988
rect 32312 26979 32364 26988
rect 32312 26945 32321 26979
rect 32321 26945 32355 26979
rect 32355 26945 32364 26979
rect 32312 26936 32364 26945
rect 29092 26911 29144 26920
rect 29092 26877 29101 26911
rect 29101 26877 29135 26911
rect 29135 26877 29144 26911
rect 29092 26868 29144 26877
rect 33324 26911 33376 26920
rect 33324 26877 33333 26911
rect 33333 26877 33367 26911
rect 33367 26877 33376 26911
rect 33324 26868 33376 26877
rect 4896 26800 4948 26852
rect 27620 26800 27672 26852
rect 29552 26800 29604 26852
rect 2596 26732 2648 26784
rect 4436 26732 4488 26784
rect 5044 26630 5096 26682
rect 5108 26630 5160 26682
rect 5172 26630 5224 26682
rect 5236 26630 5288 26682
rect 5300 26630 5352 26682
rect 13232 26630 13284 26682
rect 13296 26630 13348 26682
rect 13360 26630 13412 26682
rect 13424 26630 13476 26682
rect 13488 26630 13540 26682
rect 21420 26630 21472 26682
rect 21484 26630 21536 26682
rect 21548 26630 21600 26682
rect 21612 26630 21664 26682
rect 21676 26630 21728 26682
rect 29608 26630 29660 26682
rect 29672 26630 29724 26682
rect 29736 26630 29788 26682
rect 29800 26630 29852 26682
rect 29864 26630 29916 26682
rect 3792 26571 3844 26580
rect 3792 26537 3801 26571
rect 3801 26537 3835 26571
rect 3835 26537 3844 26571
rect 3792 26528 3844 26537
rect 4160 26528 4212 26580
rect 29368 26571 29420 26580
rect 29368 26537 29377 26571
rect 29377 26537 29411 26571
rect 29411 26537 29420 26571
rect 29368 26528 29420 26537
rect 4252 26460 4304 26512
rect 5448 26503 5500 26512
rect 5448 26469 5457 26503
rect 5457 26469 5491 26503
rect 5491 26469 5500 26503
rect 5448 26460 5500 26469
rect 29092 26460 29144 26512
rect 30104 26460 30156 26512
rect 2780 26392 2832 26444
rect 4436 26435 4488 26444
rect 4436 26401 4445 26435
rect 4445 26401 4479 26435
rect 4479 26401 4488 26435
rect 4436 26392 4488 26401
rect 5724 26435 5776 26444
rect 5724 26401 5733 26435
rect 5733 26401 5767 26435
rect 5767 26401 5776 26435
rect 5724 26392 5776 26401
rect 28080 26435 28132 26444
rect 28080 26401 28089 26435
rect 28089 26401 28123 26435
rect 28123 26401 28132 26435
rect 28080 26392 28132 26401
rect 30748 26392 30800 26444
rect 2596 26367 2648 26376
rect 2596 26333 2605 26367
rect 2605 26333 2639 26367
rect 2639 26333 2648 26367
rect 2596 26324 2648 26333
rect 3976 26324 4028 26376
rect 4160 26324 4212 26376
rect 18144 26367 18196 26376
rect 18144 26333 18153 26367
rect 18153 26333 18187 26367
rect 18187 26333 18196 26367
rect 18144 26324 18196 26333
rect 30196 26367 30248 26376
rect 30196 26333 30205 26367
rect 30205 26333 30239 26367
rect 30239 26333 30248 26367
rect 30196 26324 30248 26333
rect 30932 26367 30984 26376
rect 30932 26333 30941 26367
rect 30941 26333 30975 26367
rect 30975 26333 30984 26367
rect 30932 26324 30984 26333
rect 31668 26367 31720 26376
rect 31668 26333 31677 26367
rect 31677 26333 31711 26367
rect 31711 26333 31720 26367
rect 31668 26324 31720 26333
rect 27804 26256 27856 26308
rect 3792 26188 3844 26240
rect 16764 26188 16816 26240
rect 28816 26231 28868 26240
rect 28816 26197 28825 26231
rect 28825 26197 28859 26231
rect 28859 26197 28868 26231
rect 28816 26188 28868 26197
rect 30840 26231 30892 26240
rect 30840 26197 30849 26231
rect 30849 26197 30883 26231
rect 30883 26197 30892 26231
rect 30840 26188 30892 26197
rect 32220 26188 32272 26240
rect 33048 26231 33100 26240
rect 33048 26197 33057 26231
rect 33057 26197 33091 26231
rect 33091 26197 33100 26231
rect 33048 26188 33100 26197
rect 9138 26086 9190 26138
rect 9202 26086 9254 26138
rect 9266 26086 9318 26138
rect 9330 26086 9382 26138
rect 9394 26086 9446 26138
rect 17326 26086 17378 26138
rect 17390 26086 17442 26138
rect 17454 26086 17506 26138
rect 17518 26086 17570 26138
rect 17582 26086 17634 26138
rect 25514 26086 25566 26138
rect 25578 26086 25630 26138
rect 25642 26086 25694 26138
rect 25706 26086 25758 26138
rect 25770 26086 25822 26138
rect 33702 26086 33754 26138
rect 33766 26086 33818 26138
rect 33830 26086 33882 26138
rect 33894 26086 33946 26138
rect 33958 26086 34010 26138
rect 2872 25984 2924 26036
rect 3976 26027 4028 26036
rect 3976 25993 3985 26027
rect 3985 25993 4019 26027
rect 4019 25993 4028 26027
rect 3976 25984 4028 25993
rect 17132 25984 17184 26036
rect 30196 25984 30248 26036
rect 30380 25916 30432 25968
rect 1768 25891 1820 25900
rect 1768 25857 1777 25891
rect 1777 25857 1811 25891
rect 1811 25857 1820 25891
rect 1768 25848 1820 25857
rect 3792 25823 3844 25832
rect 3792 25789 3801 25823
rect 3801 25789 3835 25823
rect 3835 25789 3844 25823
rect 3792 25780 3844 25789
rect 4896 25780 4948 25832
rect 5908 25780 5960 25832
rect 16764 25823 16816 25832
rect 16764 25789 16773 25823
rect 16773 25789 16807 25823
rect 16807 25789 16816 25823
rect 16764 25780 16816 25789
rect 28816 25823 28868 25832
rect 28816 25789 28825 25823
rect 28825 25789 28859 25823
rect 28859 25789 28868 25823
rect 28816 25780 28868 25789
rect 33048 25984 33100 26036
rect 32312 25916 32364 25968
rect 32220 25891 32272 25900
rect 32220 25857 32229 25891
rect 32229 25857 32263 25891
rect 32263 25857 32272 25891
rect 32220 25848 32272 25857
rect 30564 25823 30616 25832
rect 30564 25789 30573 25823
rect 30573 25789 30607 25823
rect 30607 25789 30616 25823
rect 30564 25780 30616 25789
rect 31208 25823 31260 25832
rect 31208 25789 31217 25823
rect 31217 25789 31251 25823
rect 31251 25789 31260 25823
rect 31208 25780 31260 25789
rect 31300 25823 31352 25832
rect 31300 25789 31309 25823
rect 31309 25789 31343 25823
rect 31343 25789 31352 25823
rect 31300 25780 31352 25789
rect 4436 25712 4488 25764
rect 30840 25712 30892 25764
rect 31760 25644 31812 25696
rect 31944 25687 31996 25696
rect 31944 25653 31953 25687
rect 31953 25653 31987 25687
rect 31987 25653 31996 25687
rect 31944 25644 31996 25653
rect 5044 25542 5096 25594
rect 5108 25542 5160 25594
rect 5172 25542 5224 25594
rect 5236 25542 5288 25594
rect 5300 25542 5352 25594
rect 13232 25542 13284 25594
rect 13296 25542 13348 25594
rect 13360 25542 13412 25594
rect 13424 25542 13476 25594
rect 13488 25542 13540 25594
rect 21420 25542 21472 25594
rect 21484 25542 21536 25594
rect 21548 25542 21600 25594
rect 21612 25542 21664 25594
rect 21676 25542 21728 25594
rect 29608 25542 29660 25594
rect 29672 25542 29724 25594
rect 29736 25542 29788 25594
rect 29800 25542 29852 25594
rect 29864 25542 29916 25594
rect 3424 25440 3476 25492
rect 4160 25440 4212 25492
rect 29184 25440 29236 25492
rect 31208 25440 31260 25492
rect 3148 25279 3200 25288
rect 3148 25245 3157 25279
rect 3157 25245 3191 25279
rect 3191 25245 3200 25279
rect 3148 25236 3200 25245
rect 7012 25304 7064 25356
rect 26976 25304 27028 25356
rect 28540 25304 28592 25356
rect 4436 25279 4488 25288
rect 4436 25245 4445 25279
rect 4445 25245 4479 25279
rect 4479 25245 4488 25279
rect 4436 25236 4488 25245
rect 5448 25236 5500 25288
rect 28724 25279 28776 25288
rect 28724 25245 28733 25279
rect 28733 25245 28767 25279
rect 28767 25245 28776 25279
rect 28724 25236 28776 25245
rect 31576 25279 31628 25288
rect 31576 25245 31585 25279
rect 31585 25245 31619 25279
rect 31619 25245 31628 25279
rect 31576 25236 31628 25245
rect 31760 25236 31812 25288
rect 4068 25168 4120 25220
rect 31116 25168 31168 25220
rect 9138 24998 9190 25050
rect 9202 24998 9254 25050
rect 9266 24998 9318 25050
rect 9330 24998 9382 25050
rect 9394 24998 9446 25050
rect 17326 24998 17378 25050
rect 17390 24998 17442 25050
rect 17454 24998 17506 25050
rect 17518 24998 17570 25050
rect 17582 24998 17634 25050
rect 25514 24998 25566 25050
rect 25578 24998 25630 25050
rect 25642 24998 25694 25050
rect 25706 24998 25758 25050
rect 25770 24998 25822 25050
rect 33702 24998 33754 25050
rect 33766 24998 33818 25050
rect 33830 24998 33882 25050
rect 33894 24998 33946 25050
rect 33958 24998 34010 25050
rect 31300 24896 31352 24948
rect 4068 24871 4120 24880
rect 4068 24837 4077 24871
rect 4077 24837 4111 24871
rect 4111 24837 4120 24871
rect 4068 24828 4120 24837
rect 4896 24828 4948 24880
rect 31576 24828 31628 24880
rect 2596 24803 2648 24812
rect 2596 24769 2605 24803
rect 2605 24769 2639 24803
rect 2639 24769 2648 24803
rect 2596 24760 2648 24769
rect 940 24692 992 24744
rect 3332 24692 3384 24744
rect 15752 24760 15804 24812
rect 15936 24803 15988 24812
rect 15936 24769 15945 24803
rect 15945 24769 15979 24803
rect 15979 24769 15988 24803
rect 15936 24760 15988 24769
rect 30564 24803 30616 24812
rect 30564 24769 30573 24803
rect 30573 24769 30607 24803
rect 30607 24769 30616 24803
rect 30564 24760 30616 24769
rect 31944 24760 31996 24812
rect 3792 24667 3844 24676
rect 3792 24633 3801 24667
rect 3801 24633 3835 24667
rect 3835 24633 3844 24667
rect 3792 24624 3844 24633
rect 3516 24599 3568 24608
rect 3516 24565 3525 24599
rect 3525 24565 3559 24599
rect 3559 24565 3568 24599
rect 3516 24556 3568 24565
rect 3608 24599 3660 24608
rect 3608 24565 3617 24599
rect 3617 24565 3651 24599
rect 3651 24565 3660 24599
rect 3608 24556 3660 24565
rect 12072 24599 12124 24608
rect 12072 24565 12081 24599
rect 12081 24565 12115 24599
rect 12115 24565 12124 24599
rect 12072 24556 12124 24565
rect 13084 24556 13136 24608
rect 16764 24692 16816 24744
rect 31852 24735 31904 24744
rect 31852 24701 31861 24735
rect 31861 24701 31895 24735
rect 31895 24701 31904 24735
rect 31852 24692 31904 24701
rect 15752 24599 15804 24608
rect 15752 24565 15761 24599
rect 15761 24565 15795 24599
rect 15795 24565 15804 24599
rect 15752 24556 15804 24565
rect 30656 24556 30708 24608
rect 5044 24454 5096 24506
rect 5108 24454 5160 24506
rect 5172 24454 5224 24506
rect 5236 24454 5288 24506
rect 5300 24454 5352 24506
rect 13232 24454 13284 24506
rect 13296 24454 13348 24506
rect 13360 24454 13412 24506
rect 13424 24454 13476 24506
rect 13488 24454 13540 24506
rect 21420 24454 21472 24506
rect 21484 24454 21536 24506
rect 21548 24454 21600 24506
rect 21612 24454 21664 24506
rect 21676 24454 21728 24506
rect 29608 24454 29660 24506
rect 29672 24454 29724 24506
rect 29736 24454 29788 24506
rect 29800 24454 29852 24506
rect 29864 24454 29916 24506
rect 2596 24352 2648 24404
rect 2964 24395 3016 24404
rect 2964 24361 2973 24395
rect 2973 24361 3007 24395
rect 3007 24361 3016 24395
rect 2964 24352 3016 24361
rect 3332 24352 3384 24404
rect 15752 24395 15804 24404
rect 15752 24361 15761 24395
rect 15761 24361 15795 24395
rect 15795 24361 15804 24395
rect 15752 24352 15804 24361
rect 30748 24395 30800 24404
rect 30748 24361 30757 24395
rect 30757 24361 30791 24395
rect 30791 24361 30800 24395
rect 30748 24352 30800 24361
rect 3700 24216 3752 24268
rect 31300 24284 31352 24336
rect 2964 24148 3016 24200
rect 4344 24191 4396 24200
rect 4344 24157 4353 24191
rect 4353 24157 4387 24191
rect 4387 24157 4396 24191
rect 4344 24148 4396 24157
rect 4712 24148 4764 24200
rect 31392 24191 31444 24200
rect 31392 24157 31401 24191
rect 31401 24157 31435 24191
rect 31435 24157 31444 24191
rect 31392 24148 31444 24157
rect 32312 24191 32364 24200
rect 32312 24157 32321 24191
rect 32321 24157 32355 24191
rect 32355 24157 32364 24191
rect 32312 24148 32364 24157
rect 33324 24123 33376 24132
rect 33324 24089 33333 24123
rect 33333 24089 33367 24123
rect 33367 24089 33376 24123
rect 33324 24080 33376 24089
rect 31300 24055 31352 24064
rect 31300 24021 31309 24055
rect 31309 24021 31343 24055
rect 31343 24021 31352 24055
rect 31300 24012 31352 24021
rect 32036 24055 32088 24064
rect 32036 24021 32045 24055
rect 32045 24021 32079 24055
rect 32079 24021 32088 24055
rect 32036 24012 32088 24021
rect 9138 23910 9190 23962
rect 9202 23910 9254 23962
rect 9266 23910 9318 23962
rect 9330 23910 9382 23962
rect 9394 23910 9446 23962
rect 17326 23910 17378 23962
rect 17390 23910 17442 23962
rect 17454 23910 17506 23962
rect 17518 23910 17570 23962
rect 17582 23910 17634 23962
rect 25514 23910 25566 23962
rect 25578 23910 25630 23962
rect 25642 23910 25694 23962
rect 25706 23910 25758 23962
rect 25770 23910 25822 23962
rect 33702 23910 33754 23962
rect 33766 23910 33818 23962
rect 33830 23910 33882 23962
rect 33894 23910 33946 23962
rect 33958 23910 34010 23962
rect 3608 23808 3660 23860
rect 4344 23808 4396 23860
rect 2596 23715 2648 23724
rect 2596 23681 2605 23715
rect 2605 23681 2639 23715
rect 2639 23681 2648 23715
rect 2596 23672 2648 23681
rect 1584 23647 1636 23656
rect 1584 23613 1593 23647
rect 1593 23613 1627 23647
rect 1627 23613 1636 23647
rect 1584 23604 1636 23613
rect 13084 23808 13136 23860
rect 27620 23851 27672 23860
rect 27620 23817 27629 23851
rect 27629 23817 27663 23851
rect 27663 23817 27672 23851
rect 27620 23808 27672 23817
rect 31392 23808 31444 23860
rect 31852 23808 31904 23860
rect 31300 23740 31352 23792
rect 3148 23468 3200 23520
rect 25412 23604 25464 23656
rect 31668 23672 31720 23724
rect 30656 23647 30708 23656
rect 30656 23613 30665 23647
rect 30665 23613 30699 23647
rect 30699 23613 30708 23647
rect 30656 23604 30708 23613
rect 9588 23468 9640 23520
rect 25872 23468 25924 23520
rect 31300 23511 31352 23520
rect 31300 23477 31309 23511
rect 31309 23477 31343 23511
rect 31343 23477 31352 23511
rect 31300 23468 31352 23477
rect 33048 23468 33100 23520
rect 5044 23366 5096 23418
rect 5108 23366 5160 23418
rect 5172 23366 5224 23418
rect 5236 23366 5288 23418
rect 5300 23366 5352 23418
rect 13232 23366 13284 23418
rect 13296 23366 13348 23418
rect 13360 23366 13412 23418
rect 13424 23366 13476 23418
rect 13488 23366 13540 23418
rect 21420 23366 21472 23418
rect 21484 23366 21536 23418
rect 21548 23366 21600 23418
rect 21612 23366 21664 23418
rect 21676 23366 21728 23418
rect 29608 23366 29660 23418
rect 29672 23366 29724 23418
rect 29736 23366 29788 23418
rect 29800 23366 29852 23418
rect 29864 23366 29916 23418
rect 2964 23307 3016 23316
rect 2964 23273 2973 23307
rect 2973 23273 3007 23307
rect 3007 23273 3016 23307
rect 2964 23264 3016 23273
rect 4436 23307 4488 23316
rect 4436 23273 4445 23307
rect 4445 23273 4479 23307
rect 4479 23273 4488 23307
rect 4436 23264 4488 23273
rect 18144 23307 18196 23316
rect 18144 23273 18153 23307
rect 18153 23273 18187 23307
rect 18187 23273 18196 23307
rect 18144 23264 18196 23273
rect 26976 23264 27028 23316
rect 30748 23307 30800 23316
rect 30748 23273 30757 23307
rect 30757 23273 30791 23307
rect 30791 23273 30800 23307
rect 30748 23264 30800 23273
rect 4620 23239 4672 23248
rect 4620 23205 4629 23239
rect 4629 23205 4663 23239
rect 4663 23205 4672 23239
rect 4620 23196 4672 23205
rect 2596 23128 2648 23180
rect 3516 23171 3568 23180
rect 3516 23137 3525 23171
rect 3525 23137 3559 23171
rect 3559 23137 3568 23171
rect 3516 23128 3568 23137
rect 31392 23196 31444 23248
rect 31300 23128 31352 23180
rect 32312 23128 32364 23180
rect 3240 23060 3292 23112
rect 3792 23103 3844 23112
rect 3792 23069 3801 23103
rect 3801 23069 3835 23103
rect 3835 23069 3844 23103
rect 3792 23060 3844 23069
rect 17224 23060 17276 23112
rect 32220 23103 32272 23112
rect 32220 23069 32229 23103
rect 32229 23069 32263 23103
rect 32263 23069 32272 23103
rect 32220 23060 32272 23069
rect 4896 22992 4948 23044
rect 4528 22967 4580 22976
rect 4528 22933 4537 22967
rect 4537 22933 4571 22967
rect 4571 22933 4580 22967
rect 4528 22924 4580 22933
rect 25872 22967 25924 22976
rect 25872 22933 25881 22967
rect 25881 22933 25915 22967
rect 25915 22933 25924 22967
rect 25872 22924 25924 22933
rect 31300 22967 31352 22976
rect 31300 22933 31309 22967
rect 31309 22933 31343 22967
rect 31343 22933 31352 22967
rect 31300 22924 31352 22933
rect 31392 22967 31444 22976
rect 31392 22933 31401 22967
rect 31401 22933 31435 22967
rect 31435 22933 31444 22967
rect 31392 22924 31444 22933
rect 9138 22822 9190 22874
rect 9202 22822 9254 22874
rect 9266 22822 9318 22874
rect 9330 22822 9382 22874
rect 9394 22822 9446 22874
rect 17326 22822 17378 22874
rect 17390 22822 17442 22874
rect 17454 22822 17506 22874
rect 17518 22822 17570 22874
rect 17582 22822 17634 22874
rect 25514 22822 25566 22874
rect 25578 22822 25630 22874
rect 25642 22822 25694 22874
rect 25706 22822 25758 22874
rect 25770 22822 25822 22874
rect 33702 22822 33754 22874
rect 33766 22822 33818 22874
rect 33830 22822 33882 22874
rect 33894 22822 33946 22874
rect 33958 22822 34010 22874
rect 3516 22720 3568 22772
rect 28724 22720 28776 22772
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 4896 22516 4948 22568
rect 26792 22516 26844 22568
rect 31484 22559 31536 22568
rect 31484 22525 31493 22559
rect 31493 22525 31527 22559
rect 31527 22525 31536 22559
rect 31484 22516 31536 22525
rect 32036 22584 32088 22636
rect 4344 22380 4396 22432
rect 5044 22278 5096 22330
rect 5108 22278 5160 22330
rect 5172 22278 5224 22330
rect 5236 22278 5288 22330
rect 5300 22278 5352 22330
rect 13232 22278 13284 22330
rect 13296 22278 13348 22330
rect 13360 22278 13412 22330
rect 13424 22278 13476 22330
rect 13488 22278 13540 22330
rect 21420 22278 21472 22330
rect 21484 22278 21536 22330
rect 21548 22278 21600 22330
rect 21612 22278 21664 22330
rect 21676 22278 21728 22330
rect 29608 22278 29660 22330
rect 29672 22278 29724 22330
rect 29736 22278 29788 22330
rect 29800 22278 29852 22330
rect 29864 22278 29916 22330
rect 3240 22176 3292 22228
rect 32036 22176 32088 22228
rect 33048 22219 33100 22228
rect 33048 22185 33057 22219
rect 33057 22185 33091 22219
rect 33091 22185 33100 22219
rect 33048 22176 33100 22185
rect 1768 22083 1820 22092
rect 1768 22049 1777 22083
rect 1777 22049 1811 22083
rect 1811 22049 1820 22083
rect 1768 22040 1820 22049
rect 4344 22083 4396 22092
rect 4344 22049 4353 22083
rect 4353 22049 4387 22083
rect 4387 22049 4396 22083
rect 4344 22040 4396 22049
rect 31392 22040 31444 22092
rect 4528 21972 4580 22024
rect 31668 22015 31720 22024
rect 31668 21981 31677 22015
rect 31677 21981 31711 22015
rect 31711 21981 31720 22015
rect 31668 21972 31720 21981
rect 31300 21904 31352 21956
rect 4620 21836 4672 21888
rect 9138 21734 9190 21786
rect 9202 21734 9254 21786
rect 9266 21734 9318 21786
rect 9330 21734 9382 21786
rect 9394 21734 9446 21786
rect 17326 21734 17378 21786
rect 17390 21734 17442 21786
rect 17454 21734 17506 21786
rect 17518 21734 17570 21786
rect 17582 21734 17634 21786
rect 25514 21734 25566 21786
rect 25578 21734 25630 21786
rect 25642 21734 25694 21786
rect 25706 21734 25758 21786
rect 25770 21734 25822 21786
rect 33702 21734 33754 21786
rect 33766 21734 33818 21786
rect 33830 21734 33882 21786
rect 33894 21734 33946 21786
rect 33958 21734 34010 21786
rect 30748 21607 30800 21616
rect 30748 21573 30757 21607
rect 30757 21573 30791 21607
rect 30791 21573 30800 21607
rect 30748 21564 30800 21573
rect 2596 21539 2648 21548
rect 2596 21505 2605 21539
rect 2605 21505 2639 21539
rect 2639 21505 2648 21539
rect 2596 21496 2648 21505
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 940 21428 992 21480
rect 3700 21428 3752 21480
rect 4344 21428 4396 21480
rect 4804 21471 4856 21480
rect 4804 21437 4813 21471
rect 4813 21437 4847 21471
rect 4847 21437 4856 21471
rect 4804 21428 4856 21437
rect 31944 21471 31996 21480
rect 31944 21437 31953 21471
rect 31953 21437 31987 21471
rect 31987 21437 31996 21471
rect 31944 21428 31996 21437
rect 33324 21471 33376 21480
rect 33324 21437 33333 21471
rect 33333 21437 33367 21471
rect 33367 21437 33376 21471
rect 33324 21428 33376 21437
rect 31392 21360 31444 21412
rect 3516 21335 3568 21344
rect 3516 21301 3525 21335
rect 3525 21301 3559 21335
rect 3559 21301 3568 21335
rect 3516 21292 3568 21301
rect 3608 21292 3660 21344
rect 31208 21335 31260 21344
rect 31208 21301 31217 21335
rect 31217 21301 31251 21335
rect 31251 21301 31260 21335
rect 31208 21292 31260 21301
rect 31300 21335 31352 21344
rect 31300 21301 31309 21335
rect 31309 21301 31343 21335
rect 31343 21301 31352 21335
rect 31300 21292 31352 21301
rect 5044 21190 5096 21242
rect 5108 21190 5160 21242
rect 5172 21190 5224 21242
rect 5236 21190 5288 21242
rect 5300 21190 5352 21242
rect 13232 21190 13284 21242
rect 13296 21190 13348 21242
rect 13360 21190 13412 21242
rect 13424 21190 13476 21242
rect 13488 21190 13540 21242
rect 21420 21190 21472 21242
rect 21484 21190 21536 21242
rect 21548 21190 21600 21242
rect 21612 21190 21664 21242
rect 21676 21190 21728 21242
rect 29608 21190 29660 21242
rect 29672 21190 29724 21242
rect 29736 21190 29788 21242
rect 29800 21190 29852 21242
rect 29864 21190 29916 21242
rect 3700 21088 3752 21140
rect 3792 21131 3844 21140
rect 3792 21097 3801 21131
rect 3801 21097 3835 21131
rect 3835 21097 3844 21131
rect 3792 21088 3844 21097
rect 25412 21131 25464 21140
rect 25412 21097 25421 21131
rect 25421 21097 25455 21131
rect 25455 21097 25464 21131
rect 25412 21088 25464 21097
rect 31944 21088 31996 21140
rect 1768 20995 1820 21004
rect 1768 20961 1777 20995
rect 1777 20961 1811 20995
rect 1811 20961 1820 20995
rect 1768 20952 1820 20961
rect 31300 20952 31352 21004
rect 3608 20884 3660 20936
rect 4528 20884 4580 20936
rect 24768 20927 24820 20936
rect 24768 20893 24777 20927
rect 24777 20893 24811 20927
rect 24811 20893 24820 20927
rect 24768 20884 24820 20893
rect 31208 20884 31260 20936
rect 31668 20927 31720 20936
rect 31668 20893 31677 20927
rect 31677 20893 31711 20927
rect 31711 20893 31720 20927
rect 31668 20884 31720 20893
rect 9588 20748 9640 20800
rect 10324 20748 10376 20800
rect 31576 20791 31628 20800
rect 31576 20757 31585 20791
rect 31585 20757 31619 20791
rect 31619 20757 31628 20791
rect 31576 20748 31628 20757
rect 9138 20646 9190 20698
rect 9202 20646 9254 20698
rect 9266 20646 9318 20698
rect 9330 20646 9382 20698
rect 9394 20646 9446 20698
rect 17326 20646 17378 20698
rect 17390 20646 17442 20698
rect 17454 20646 17506 20698
rect 17518 20646 17570 20698
rect 17582 20646 17634 20698
rect 25514 20646 25566 20698
rect 25578 20646 25630 20698
rect 25642 20646 25694 20698
rect 25706 20646 25758 20698
rect 25770 20646 25822 20698
rect 33702 20646 33754 20698
rect 33766 20646 33818 20698
rect 33830 20646 33882 20698
rect 33894 20646 33946 20698
rect 33958 20646 34010 20698
rect 2596 20476 2648 20528
rect 32312 20476 32364 20528
rect 3608 20383 3660 20392
rect 3608 20349 3617 20383
rect 3617 20349 3651 20383
rect 3651 20349 3660 20383
rect 3608 20340 3660 20349
rect 31576 20340 31628 20392
rect 31852 20340 31904 20392
rect 5044 20102 5096 20154
rect 5108 20102 5160 20154
rect 5172 20102 5224 20154
rect 5236 20102 5288 20154
rect 5300 20102 5352 20154
rect 13232 20102 13284 20154
rect 13296 20102 13348 20154
rect 13360 20102 13412 20154
rect 13424 20102 13476 20154
rect 13488 20102 13540 20154
rect 21420 20102 21472 20154
rect 21484 20102 21536 20154
rect 21548 20102 21600 20154
rect 21612 20102 21664 20154
rect 21676 20102 21728 20154
rect 29608 20102 29660 20154
rect 29672 20102 29724 20154
rect 29736 20102 29788 20154
rect 29800 20102 29852 20154
rect 29864 20102 29916 20154
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 30748 20000 30800 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 31852 19975 31904 19984
rect 31852 19941 31861 19975
rect 31861 19941 31895 19975
rect 31895 19941 31904 19975
rect 31852 19932 31904 19941
rect 4436 19839 4488 19848
rect 4436 19805 4445 19839
rect 4445 19805 4479 19839
rect 4479 19805 4488 19839
rect 4436 19796 4488 19805
rect 3240 19728 3292 19780
rect 18052 19728 18104 19780
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 3792 19703 3844 19712
rect 3792 19669 3801 19703
rect 3801 19669 3835 19703
rect 3835 19669 3844 19703
rect 3792 19660 3844 19669
rect 28540 19796 28592 19848
rect 32588 19771 32640 19780
rect 32588 19737 32597 19771
rect 32597 19737 32631 19771
rect 32631 19737 32640 19771
rect 32588 19728 32640 19737
rect 25412 19660 25464 19712
rect 26976 19660 27028 19712
rect 32036 19703 32088 19712
rect 32036 19669 32045 19703
rect 32045 19669 32079 19703
rect 32079 19669 32088 19703
rect 32036 19660 32088 19669
rect 9138 19558 9190 19610
rect 9202 19558 9254 19610
rect 9266 19558 9318 19610
rect 9330 19558 9382 19610
rect 9394 19558 9446 19610
rect 17326 19558 17378 19610
rect 17390 19558 17442 19610
rect 17454 19558 17506 19610
rect 17518 19558 17570 19610
rect 17582 19558 17634 19610
rect 25514 19558 25566 19610
rect 25578 19558 25630 19610
rect 25642 19558 25694 19610
rect 25706 19558 25758 19610
rect 25770 19558 25822 19610
rect 33702 19558 33754 19610
rect 33766 19558 33818 19610
rect 33830 19558 33882 19610
rect 33894 19558 33946 19610
rect 33958 19558 34010 19610
rect 3240 19456 3292 19508
rect 26792 19499 26844 19508
rect 26792 19465 26801 19499
rect 26801 19465 26835 19499
rect 26835 19465 26844 19499
rect 26792 19456 26844 19465
rect 26976 19456 27028 19508
rect 25504 19388 25556 19440
rect 940 19320 992 19372
rect 2596 19363 2648 19372
rect 2596 19329 2605 19363
rect 2605 19329 2639 19363
rect 2639 19329 2648 19363
rect 2596 19320 2648 19329
rect 4436 19320 4488 19372
rect 25412 19363 25464 19372
rect 25412 19329 25428 19363
rect 25428 19329 25462 19363
rect 25462 19329 25464 19363
rect 25412 19320 25464 19329
rect 32588 19320 32640 19372
rect 33324 19363 33376 19372
rect 33324 19329 33333 19363
rect 33333 19329 33367 19363
rect 33367 19329 33376 19363
rect 33324 19320 33376 19329
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 3700 19295 3752 19304
rect 3700 19261 3709 19295
rect 3709 19261 3743 19295
rect 3743 19261 3752 19295
rect 3700 19252 3752 19261
rect 4804 19295 4856 19304
rect 4804 19261 4813 19295
rect 4813 19261 4847 19295
rect 4847 19261 4856 19295
rect 4804 19252 4856 19261
rect 31300 19295 31352 19304
rect 31300 19261 31309 19295
rect 31309 19261 31343 19295
rect 31343 19261 31352 19295
rect 31300 19252 31352 19261
rect 3608 19184 3660 19236
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 31944 19159 31996 19168
rect 31944 19125 31953 19159
rect 31953 19125 31987 19159
rect 31987 19125 31996 19159
rect 31944 19116 31996 19125
rect 5044 19014 5096 19066
rect 5108 19014 5160 19066
rect 5172 19014 5224 19066
rect 5236 19014 5288 19066
rect 5300 19014 5352 19066
rect 13232 19014 13284 19066
rect 13296 19014 13348 19066
rect 13360 19014 13412 19066
rect 13424 19014 13476 19066
rect 13488 19014 13540 19066
rect 21420 19014 21472 19066
rect 21484 19014 21536 19066
rect 21548 19014 21600 19066
rect 21612 19014 21664 19066
rect 21676 19014 21728 19066
rect 29608 19014 29660 19066
rect 29672 19014 29724 19066
rect 29736 19014 29788 19066
rect 29800 19014 29852 19066
rect 29864 19014 29916 19066
rect 2872 18955 2924 18964
rect 2872 18921 2881 18955
rect 2881 18921 2915 18955
rect 2915 18921 2924 18955
rect 2872 18912 2924 18921
rect 3700 18912 3752 18964
rect 1952 18887 2004 18896
rect 1952 18853 1961 18887
rect 1961 18853 1995 18887
rect 1995 18853 2004 18887
rect 8944 18912 8996 18964
rect 18052 18955 18104 18964
rect 18052 18921 18061 18955
rect 18061 18921 18095 18955
rect 18095 18921 18104 18955
rect 18052 18912 18104 18921
rect 1952 18844 2004 18853
rect 4712 18844 4764 18896
rect 19432 18844 19484 18896
rect 2596 18776 2648 18828
rect 3148 18776 3200 18828
rect 4252 18776 4304 18828
rect 4804 18776 4856 18828
rect 31668 18819 31720 18828
rect 31668 18785 31677 18819
rect 31677 18785 31711 18819
rect 31711 18785 31720 18819
rect 31668 18776 31720 18785
rect 3792 18708 3844 18760
rect 4160 18708 4212 18760
rect 30288 18640 30340 18692
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 3884 18572 3936 18624
rect 31576 18615 31628 18624
rect 31576 18581 31585 18615
rect 31585 18581 31619 18615
rect 31619 18581 31628 18615
rect 31576 18572 31628 18581
rect 32036 18640 32088 18692
rect 9138 18470 9190 18522
rect 9202 18470 9254 18522
rect 9266 18470 9318 18522
rect 9330 18470 9382 18522
rect 9394 18470 9446 18522
rect 17326 18470 17378 18522
rect 17390 18470 17442 18522
rect 17454 18470 17506 18522
rect 17518 18470 17570 18522
rect 17582 18470 17634 18522
rect 25514 18470 25566 18522
rect 25578 18470 25630 18522
rect 25642 18470 25694 18522
rect 25706 18470 25758 18522
rect 25770 18470 25822 18522
rect 33702 18470 33754 18522
rect 33766 18470 33818 18522
rect 33830 18470 33882 18522
rect 33894 18470 33946 18522
rect 33958 18470 34010 18522
rect 1952 18368 2004 18420
rect 3792 18368 3844 18420
rect 30380 18368 30432 18420
rect 30748 18368 30800 18420
rect 31024 18411 31076 18420
rect 31024 18377 31033 18411
rect 31033 18377 31067 18411
rect 31067 18377 31076 18411
rect 31024 18368 31076 18377
rect 31300 18411 31352 18420
rect 31300 18377 31309 18411
rect 31309 18377 31343 18411
rect 31343 18377 31352 18411
rect 31300 18368 31352 18377
rect 31576 18232 31628 18284
rect 31944 18232 31996 18284
rect 4804 18207 4856 18216
rect 1308 18096 1360 18148
rect 4804 18173 4813 18207
rect 4813 18173 4847 18207
rect 4847 18173 4856 18207
rect 4804 18164 4856 18173
rect 32496 18207 32548 18216
rect 32496 18173 32505 18207
rect 32505 18173 32539 18207
rect 32539 18173 32548 18207
rect 32496 18164 32548 18173
rect 4436 18139 4488 18148
rect 4436 18105 4445 18139
rect 4445 18105 4479 18139
rect 4479 18105 4488 18139
rect 4436 18096 4488 18105
rect 4252 18028 4304 18080
rect 5044 17926 5096 17978
rect 5108 17926 5160 17978
rect 5172 17926 5224 17978
rect 5236 17926 5288 17978
rect 5300 17926 5352 17978
rect 13232 17926 13284 17978
rect 13296 17926 13348 17978
rect 13360 17926 13412 17978
rect 13424 17926 13476 17978
rect 13488 17926 13540 17978
rect 21420 17926 21472 17978
rect 21484 17926 21536 17978
rect 21548 17926 21600 17978
rect 21612 17926 21664 17978
rect 21676 17926 21728 17978
rect 29608 17926 29660 17978
rect 29672 17926 29724 17978
rect 29736 17926 29788 17978
rect 29800 17926 29852 17978
rect 29864 17926 29916 17978
rect 4160 17824 4212 17876
rect 21824 17824 21876 17876
rect 4344 17756 4396 17808
rect 24768 17824 24820 17876
rect 31300 17756 31352 17808
rect 1768 17731 1820 17740
rect 1768 17697 1777 17731
rect 1777 17697 1811 17731
rect 1811 17697 1820 17731
rect 1768 17688 1820 17697
rect 4804 17688 4856 17740
rect 30288 17731 30340 17740
rect 30288 17697 30297 17731
rect 30297 17697 30331 17731
rect 30331 17697 30340 17731
rect 31024 17731 31076 17740
rect 30288 17688 30340 17697
rect 31024 17697 31033 17731
rect 31033 17697 31067 17731
rect 31067 17697 31076 17731
rect 31024 17688 31076 17697
rect 33324 17731 33376 17740
rect 33324 17697 33333 17731
rect 33333 17697 33367 17731
rect 33367 17697 33376 17731
rect 33324 17688 33376 17697
rect 4252 17620 4304 17672
rect 4620 17620 4672 17672
rect 10324 17620 10376 17672
rect 3516 17484 3568 17536
rect 4252 17484 4304 17536
rect 22008 17620 22060 17672
rect 24952 17663 25004 17672
rect 24952 17629 24961 17663
rect 24961 17629 24995 17663
rect 24995 17629 25004 17663
rect 24952 17620 25004 17629
rect 30380 17620 30432 17672
rect 32036 17663 32088 17672
rect 32036 17629 32045 17663
rect 32045 17629 32079 17663
rect 32079 17629 32088 17663
rect 32036 17620 32088 17629
rect 32496 17620 32548 17672
rect 19064 17595 19116 17604
rect 19064 17561 19073 17595
rect 19073 17561 19107 17595
rect 19107 17561 19116 17595
rect 19064 17552 19116 17561
rect 19156 17552 19208 17604
rect 25872 17552 25924 17604
rect 30748 17527 30800 17536
rect 30748 17493 30757 17527
rect 30757 17493 30791 17527
rect 30791 17493 30800 17527
rect 30748 17484 30800 17493
rect 31392 17527 31444 17536
rect 31392 17493 31401 17527
rect 31401 17493 31435 17527
rect 31435 17493 31444 17527
rect 31392 17484 31444 17493
rect 9138 17382 9190 17434
rect 9202 17382 9254 17434
rect 9266 17382 9318 17434
rect 9330 17382 9382 17434
rect 9394 17382 9446 17434
rect 17326 17382 17378 17434
rect 17390 17382 17442 17434
rect 17454 17382 17506 17434
rect 17518 17382 17570 17434
rect 17582 17382 17634 17434
rect 25514 17382 25566 17434
rect 25578 17382 25630 17434
rect 25642 17382 25694 17434
rect 25706 17382 25758 17434
rect 25770 17382 25822 17434
rect 33702 17382 33754 17434
rect 33766 17382 33818 17434
rect 33830 17382 33882 17434
rect 33894 17382 33946 17434
rect 33958 17382 34010 17434
rect 4528 17280 4580 17332
rect 32036 17280 32088 17332
rect 30748 17212 30800 17264
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 4160 17144 4212 17196
rect 31944 17187 31996 17196
rect 31944 17153 31953 17187
rect 31953 17153 31987 17187
rect 31987 17153 31996 17187
rect 31944 17144 31996 17153
rect 3332 17119 3384 17128
rect 3332 17085 3341 17119
rect 3341 17085 3375 17119
rect 3375 17085 3384 17119
rect 3332 17076 3384 17085
rect 4528 17119 4580 17128
rect 4528 17085 4537 17119
rect 4537 17085 4571 17119
rect 4571 17085 4580 17119
rect 4528 17076 4580 17085
rect 31484 17119 31536 17128
rect 31484 17085 31493 17119
rect 31493 17085 31527 17119
rect 31527 17085 31536 17119
rect 31484 17076 31536 17085
rect 31668 17076 31720 17128
rect 7472 17008 7524 17060
rect 3976 16983 4028 16992
rect 3976 16949 3985 16983
rect 3985 16949 4019 16983
rect 4019 16949 4028 16983
rect 3976 16940 4028 16949
rect 5044 16838 5096 16890
rect 5108 16838 5160 16890
rect 5172 16838 5224 16890
rect 5236 16838 5288 16890
rect 5300 16838 5352 16890
rect 13232 16838 13284 16890
rect 13296 16838 13348 16890
rect 13360 16838 13412 16890
rect 13424 16838 13476 16890
rect 13488 16838 13540 16890
rect 21420 16838 21472 16890
rect 21484 16838 21536 16890
rect 21548 16838 21600 16890
rect 21612 16838 21664 16890
rect 21676 16838 21728 16890
rect 29608 16838 29660 16890
rect 29672 16838 29724 16890
rect 29736 16838 29788 16890
rect 29800 16838 29852 16890
rect 29864 16838 29916 16890
rect 3332 16736 3384 16788
rect 4160 16736 4212 16788
rect 21824 16736 21876 16788
rect 31944 16736 31996 16788
rect 4620 16711 4672 16720
rect 4620 16677 4629 16711
rect 4629 16677 4663 16711
rect 4663 16677 4672 16711
rect 4620 16668 4672 16677
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 19524 16643 19576 16652
rect 19524 16609 19533 16643
rect 19533 16609 19567 16643
rect 19567 16609 19576 16643
rect 19524 16600 19576 16609
rect 3884 16532 3936 16584
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 20720 16532 20772 16584
rect 31392 16600 31444 16652
rect 32220 16575 32272 16584
rect 32220 16541 32229 16575
rect 32229 16541 32263 16575
rect 32263 16541 32272 16575
rect 32220 16532 32272 16541
rect 4528 16396 4580 16448
rect 4804 16396 4856 16448
rect 24952 16464 25004 16516
rect 28540 16396 28592 16448
rect 31392 16439 31444 16448
rect 31392 16405 31401 16439
rect 31401 16405 31435 16439
rect 31435 16405 31444 16439
rect 31392 16396 31444 16405
rect 9138 16294 9190 16346
rect 9202 16294 9254 16346
rect 9266 16294 9318 16346
rect 9330 16294 9382 16346
rect 9394 16294 9446 16346
rect 17326 16294 17378 16346
rect 17390 16294 17442 16346
rect 17454 16294 17506 16346
rect 17518 16294 17570 16346
rect 17582 16294 17634 16346
rect 25514 16294 25566 16346
rect 25578 16294 25630 16346
rect 25642 16294 25694 16346
rect 25706 16294 25758 16346
rect 25770 16294 25822 16346
rect 33702 16294 33754 16346
rect 33766 16294 33818 16346
rect 33830 16294 33882 16346
rect 33894 16294 33946 16346
rect 33958 16294 34010 16346
rect 4344 16192 4396 16244
rect 30380 16192 30432 16244
rect 4252 16124 4304 16176
rect 32220 16192 32272 16244
rect 3976 16056 4028 16108
rect 4896 16099 4948 16108
rect 4896 16065 4905 16099
rect 4905 16065 4939 16099
rect 4939 16065 4948 16099
rect 4896 16056 4948 16065
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 32312 16099 32364 16108
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 1768 15988 1820 16040
rect 4344 16031 4396 16040
rect 4344 15997 4353 16031
rect 4353 15997 4387 16031
rect 4387 15997 4396 16031
rect 4344 15988 4396 15997
rect 33324 16031 33376 16040
rect 33324 15997 33333 16031
rect 33333 15997 33367 16031
rect 33367 15997 33376 16031
rect 33324 15988 33376 15997
rect 3424 15852 3476 15904
rect 31760 15852 31812 15904
rect 5044 15750 5096 15802
rect 5108 15750 5160 15802
rect 5172 15750 5224 15802
rect 5236 15750 5288 15802
rect 5300 15750 5352 15802
rect 13232 15750 13284 15802
rect 13296 15750 13348 15802
rect 13360 15750 13412 15802
rect 13424 15750 13476 15802
rect 13488 15750 13540 15802
rect 21420 15750 21472 15802
rect 21484 15750 21536 15802
rect 21548 15750 21600 15802
rect 21612 15750 21664 15802
rect 21676 15750 21728 15802
rect 29608 15750 29660 15802
rect 29672 15750 29724 15802
rect 29736 15750 29788 15802
rect 29800 15750 29852 15802
rect 29864 15750 29916 15802
rect 4344 15648 4396 15700
rect 4896 15648 4948 15700
rect 25412 15648 25464 15700
rect 1584 15555 1636 15564
rect 1584 15521 1593 15555
rect 1593 15521 1627 15555
rect 1627 15521 1636 15555
rect 1584 15512 1636 15521
rect 24952 15623 25004 15632
rect 24952 15589 24961 15623
rect 24961 15589 24995 15623
rect 24995 15589 25004 15623
rect 24952 15580 25004 15589
rect 30288 15512 30340 15564
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 10600 15444 10652 15496
rect 30840 15487 30892 15496
rect 30840 15453 30849 15487
rect 30849 15453 30883 15487
rect 30883 15453 30892 15487
rect 30840 15444 30892 15453
rect 31668 15487 31720 15496
rect 31668 15453 31677 15487
rect 31677 15453 31711 15487
rect 31711 15453 31720 15487
rect 31668 15444 31720 15453
rect 31760 15444 31812 15496
rect 3976 15376 4028 15428
rect 24584 15419 24636 15428
rect 24584 15385 24593 15419
rect 24593 15385 24627 15419
rect 24627 15385 24636 15419
rect 24584 15376 24636 15385
rect 25228 15376 25280 15428
rect 2964 15351 3016 15360
rect 2964 15317 2973 15351
rect 2973 15317 3007 15351
rect 3007 15317 3016 15351
rect 2964 15308 3016 15317
rect 31576 15351 31628 15360
rect 31576 15317 31585 15351
rect 31585 15317 31619 15351
rect 31619 15317 31628 15351
rect 31576 15308 31628 15317
rect 33048 15351 33100 15360
rect 33048 15317 33057 15351
rect 33057 15317 33091 15351
rect 33091 15317 33100 15351
rect 33048 15308 33100 15317
rect 9138 15206 9190 15258
rect 9202 15206 9254 15258
rect 9266 15206 9318 15258
rect 9330 15206 9382 15258
rect 9394 15206 9446 15258
rect 17326 15206 17378 15258
rect 17390 15206 17442 15258
rect 17454 15206 17506 15258
rect 17518 15206 17570 15258
rect 17582 15206 17634 15258
rect 25514 15206 25566 15258
rect 25578 15206 25630 15258
rect 25642 15206 25694 15258
rect 25706 15206 25758 15258
rect 25770 15206 25822 15258
rect 33702 15206 33754 15258
rect 33766 15206 33818 15258
rect 33830 15206 33882 15258
rect 33894 15206 33946 15258
rect 33958 15206 34010 15258
rect 3792 15104 3844 15156
rect 1768 14900 1820 14952
rect 18512 15036 18564 15088
rect 24584 15104 24636 15156
rect 30840 15104 30892 15156
rect 32312 15036 32364 15088
rect 3700 14968 3752 15020
rect 11612 14968 11664 15020
rect 12716 14900 12768 14952
rect 20720 14968 20772 15020
rect 31576 14968 31628 15020
rect 33048 14968 33100 15020
rect 4344 14764 4396 14816
rect 5448 14764 5500 14816
rect 23480 14832 23532 14884
rect 30380 14900 30432 14952
rect 30564 14943 30616 14952
rect 30564 14909 30573 14943
rect 30573 14909 30607 14943
rect 30607 14909 30616 14943
rect 30564 14900 30616 14909
rect 30288 14875 30340 14884
rect 30288 14841 30297 14875
rect 30297 14841 30331 14875
rect 30331 14841 30340 14875
rect 30288 14832 30340 14841
rect 31760 14832 31812 14884
rect 18604 14807 18656 14816
rect 18604 14773 18613 14807
rect 18613 14773 18647 14807
rect 18647 14773 18656 14807
rect 18604 14764 18656 14773
rect 19524 14764 19576 14816
rect 19800 14807 19852 14816
rect 19800 14773 19809 14807
rect 19809 14773 19843 14807
rect 19843 14773 19852 14807
rect 19800 14764 19852 14773
rect 30012 14764 30064 14816
rect 31300 14764 31352 14816
rect 5044 14662 5096 14714
rect 5108 14662 5160 14714
rect 5172 14662 5224 14714
rect 5236 14662 5288 14714
rect 5300 14662 5352 14714
rect 13232 14662 13284 14714
rect 13296 14662 13348 14714
rect 13360 14662 13412 14714
rect 13424 14662 13476 14714
rect 13488 14662 13540 14714
rect 21420 14662 21472 14714
rect 21484 14662 21536 14714
rect 21548 14662 21600 14714
rect 21612 14662 21664 14714
rect 21676 14662 21728 14714
rect 29608 14662 29660 14714
rect 29672 14662 29724 14714
rect 29736 14662 29788 14714
rect 29800 14662 29852 14714
rect 29864 14662 29916 14714
rect 3700 14560 3752 14612
rect 4344 14603 4396 14612
rect 4344 14569 4353 14603
rect 4353 14569 4387 14603
rect 4387 14569 4396 14603
rect 4344 14560 4396 14569
rect 11612 14603 11664 14612
rect 11612 14569 11621 14603
rect 11621 14569 11655 14603
rect 11655 14569 11664 14603
rect 11612 14560 11664 14569
rect 18512 14603 18564 14612
rect 18512 14569 18521 14603
rect 18521 14569 18555 14603
rect 18555 14569 18564 14603
rect 18512 14560 18564 14569
rect 18604 14560 18656 14612
rect 19156 14560 19208 14612
rect 3976 14535 4028 14544
rect 3976 14501 3985 14535
rect 3985 14501 4019 14535
rect 4019 14501 4028 14535
rect 3976 14492 4028 14501
rect 4436 14535 4488 14544
rect 4436 14501 4445 14535
rect 4445 14501 4479 14535
rect 4479 14501 4488 14535
rect 4436 14492 4488 14501
rect 11428 14535 11480 14544
rect 11428 14501 11437 14535
rect 11437 14501 11471 14535
rect 11471 14501 11480 14535
rect 11428 14492 11480 14501
rect 1584 14467 1636 14476
rect 1584 14433 1593 14467
rect 1593 14433 1627 14467
rect 1627 14433 1636 14467
rect 1584 14424 1636 14433
rect 3424 14467 3476 14476
rect 3424 14433 3433 14467
rect 3433 14433 3467 14467
rect 3467 14433 3476 14467
rect 3424 14424 3476 14433
rect 2596 14399 2648 14408
rect 2596 14365 2605 14399
rect 2605 14365 2639 14399
rect 2639 14365 2648 14399
rect 2596 14356 2648 14365
rect 4804 14331 4856 14340
rect 4804 14297 4813 14331
rect 4813 14297 4847 14331
rect 4847 14297 4856 14331
rect 4804 14288 4856 14297
rect 18880 14535 18932 14544
rect 18880 14501 18889 14535
rect 18889 14501 18923 14535
rect 18923 14501 18932 14535
rect 18880 14492 18932 14501
rect 24400 14492 24452 14544
rect 31668 14467 31720 14476
rect 31668 14433 31677 14467
rect 31677 14433 31711 14467
rect 31711 14433 31720 14467
rect 31668 14424 31720 14433
rect 31576 14399 31628 14408
rect 31576 14365 31585 14399
rect 31585 14365 31619 14399
rect 31619 14365 31628 14399
rect 31576 14356 31628 14365
rect 31760 14356 31812 14408
rect 31116 14288 31168 14340
rect 2872 14263 2924 14272
rect 2872 14229 2881 14263
rect 2881 14229 2915 14263
rect 2915 14229 2924 14263
rect 2872 14220 2924 14229
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 20996 14263 21048 14272
rect 20996 14229 21005 14263
rect 21005 14229 21039 14263
rect 21039 14229 21048 14263
rect 20996 14220 21048 14229
rect 31024 14220 31076 14272
rect 9138 14118 9190 14170
rect 9202 14118 9254 14170
rect 9266 14118 9318 14170
rect 9330 14118 9382 14170
rect 9394 14118 9446 14170
rect 17326 14118 17378 14170
rect 17390 14118 17442 14170
rect 17454 14118 17506 14170
rect 17518 14118 17570 14170
rect 17582 14118 17634 14170
rect 25514 14118 25566 14170
rect 25578 14118 25630 14170
rect 25642 14118 25694 14170
rect 25706 14118 25758 14170
rect 25770 14118 25822 14170
rect 33702 14118 33754 14170
rect 33766 14118 33818 14170
rect 33830 14118 33882 14170
rect 33894 14118 33946 14170
rect 33958 14118 34010 14170
rect 2596 14016 2648 14068
rect 2964 14016 3016 14068
rect 19340 14016 19392 14068
rect 19800 14016 19852 14068
rect 30564 14059 30616 14068
rect 30564 14025 30573 14059
rect 30573 14025 30607 14059
rect 30607 14025 30616 14059
rect 30564 14016 30616 14025
rect 31576 13948 31628 14000
rect 2780 13880 2832 13932
rect 20996 13880 21048 13932
rect 22008 13880 22060 13932
rect 26516 13880 26568 13932
rect 31208 13880 31260 13932
rect 1308 13812 1360 13864
rect 3424 13744 3476 13796
rect 13636 13812 13688 13864
rect 15936 13812 15988 13864
rect 30012 13855 30064 13864
rect 30012 13821 30021 13855
rect 30021 13821 30055 13855
rect 30055 13821 30064 13855
rect 30012 13812 30064 13821
rect 30564 13812 30616 13864
rect 31024 13812 31076 13864
rect 31300 13855 31352 13864
rect 31300 13821 31309 13855
rect 31309 13821 31343 13855
rect 31343 13821 31352 13855
rect 31300 13812 31352 13821
rect 4344 13719 4396 13728
rect 4344 13685 4353 13719
rect 4353 13685 4387 13719
rect 4387 13685 4396 13719
rect 4344 13676 4396 13685
rect 4804 13676 4856 13728
rect 31760 13676 31812 13728
rect 5044 13574 5096 13626
rect 5108 13574 5160 13626
rect 5172 13574 5224 13626
rect 5236 13574 5288 13626
rect 5300 13574 5352 13626
rect 13232 13574 13284 13626
rect 13296 13574 13348 13626
rect 13360 13574 13412 13626
rect 13424 13574 13476 13626
rect 13488 13574 13540 13626
rect 21420 13574 21472 13626
rect 21484 13574 21536 13626
rect 21548 13574 21600 13626
rect 21612 13574 21664 13626
rect 21676 13574 21728 13626
rect 29608 13574 29660 13626
rect 29672 13574 29724 13626
rect 29736 13574 29788 13626
rect 29800 13574 29852 13626
rect 29864 13574 29916 13626
rect 10600 13447 10652 13456
rect 10600 13413 10609 13447
rect 10609 13413 10643 13447
rect 10643 13413 10652 13447
rect 10600 13404 10652 13413
rect 2780 13336 2832 13388
rect 4436 13379 4488 13388
rect 4436 13345 4445 13379
rect 4445 13345 4479 13379
rect 4479 13345 4488 13379
rect 4436 13336 4488 13345
rect 2872 13268 2924 13320
rect 4252 13268 4304 13320
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 19708 13268 19760 13320
rect 30932 13268 30984 13320
rect 31208 13268 31260 13320
rect 31760 13268 31812 13320
rect 2872 13175 2924 13184
rect 2872 13141 2881 13175
rect 2881 13141 2915 13175
rect 2915 13141 2924 13175
rect 2872 13132 2924 13141
rect 3424 13132 3476 13184
rect 11152 13132 11204 13184
rect 11980 13132 12032 13184
rect 13636 13132 13688 13184
rect 20352 13132 20404 13184
rect 30840 13175 30892 13184
rect 30840 13141 30849 13175
rect 30849 13141 30883 13175
rect 30883 13141 30892 13175
rect 30840 13132 30892 13141
rect 31576 13175 31628 13184
rect 31576 13141 31585 13175
rect 31585 13141 31619 13175
rect 31619 13141 31628 13175
rect 31576 13132 31628 13141
rect 9138 13030 9190 13082
rect 9202 13030 9254 13082
rect 9266 13030 9318 13082
rect 9330 13030 9382 13082
rect 9394 13030 9446 13082
rect 17326 13030 17378 13082
rect 17390 13030 17442 13082
rect 17454 13030 17506 13082
rect 17518 13030 17570 13082
rect 17582 13030 17634 13082
rect 25514 13030 25566 13082
rect 25578 13030 25630 13082
rect 25642 13030 25694 13082
rect 25706 13030 25758 13082
rect 25770 13030 25822 13082
rect 33702 13030 33754 13082
rect 33766 13030 33818 13082
rect 33830 13030 33882 13082
rect 33894 13030 33946 13082
rect 33958 13030 34010 13082
rect 4252 12928 4304 12980
rect 23480 12928 23532 12980
rect 31208 12971 31260 12980
rect 31208 12937 31217 12971
rect 31217 12937 31251 12971
rect 31251 12937 31260 12971
rect 31208 12928 31260 12937
rect 4344 12860 4396 12912
rect 4436 12860 4488 12912
rect 3516 12792 3568 12844
rect 26976 12792 27028 12844
rect 30840 12792 30892 12844
rect 30932 12792 30984 12844
rect 31576 12792 31628 12844
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 3976 12767 4028 12776
rect 3976 12733 3985 12767
rect 3985 12733 4019 12767
rect 4019 12733 4028 12767
rect 3976 12724 4028 12733
rect 32496 12767 32548 12776
rect 32496 12733 32505 12767
rect 32505 12733 32539 12767
rect 32539 12733 32548 12767
rect 32496 12724 32548 12733
rect 3148 12631 3200 12640
rect 3148 12597 3157 12631
rect 3157 12597 3191 12631
rect 3191 12597 3200 12631
rect 3148 12588 3200 12597
rect 4804 12588 4856 12640
rect 23664 12631 23716 12640
rect 23664 12597 23673 12631
rect 23673 12597 23707 12631
rect 23707 12597 23716 12631
rect 23664 12588 23716 12597
rect 5044 12486 5096 12538
rect 5108 12486 5160 12538
rect 5172 12486 5224 12538
rect 5236 12486 5288 12538
rect 5300 12486 5352 12538
rect 13232 12486 13284 12538
rect 13296 12486 13348 12538
rect 13360 12486 13412 12538
rect 13424 12486 13476 12538
rect 13488 12486 13540 12538
rect 21420 12486 21472 12538
rect 21484 12486 21536 12538
rect 21548 12486 21600 12538
rect 21612 12486 21664 12538
rect 21676 12486 21728 12538
rect 29608 12486 29660 12538
rect 29672 12486 29724 12538
rect 29736 12486 29788 12538
rect 29800 12486 29852 12538
rect 29864 12486 29916 12538
rect 3976 12384 4028 12436
rect 30564 12384 30616 12436
rect 4252 12316 4304 12368
rect 3148 12248 3200 12300
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 24400 12291 24452 12300
rect 24400 12257 24409 12291
rect 24409 12257 24443 12291
rect 24443 12257 24452 12291
rect 24400 12248 24452 12257
rect 30932 12316 30984 12368
rect 33324 12291 33376 12300
rect 33324 12257 33333 12291
rect 33333 12257 33367 12291
rect 33367 12257 33376 12291
rect 33324 12248 33376 12257
rect 2872 12180 2924 12232
rect 3792 12223 3844 12232
rect 3792 12189 3801 12223
rect 3801 12189 3835 12223
rect 3835 12189 3844 12223
rect 3792 12180 3844 12189
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 11428 12180 11480 12232
rect 32036 12223 32088 12232
rect 32036 12189 32045 12223
rect 32045 12189 32079 12223
rect 32079 12189 32088 12223
rect 32036 12180 32088 12189
rect 32496 12180 32548 12232
rect 4804 12112 4856 12164
rect 2596 12044 2648 12096
rect 4436 12087 4488 12096
rect 4436 12053 4445 12087
rect 4445 12053 4479 12087
rect 4479 12053 4488 12087
rect 4436 12044 4488 12053
rect 4528 12087 4580 12096
rect 4528 12053 4537 12087
rect 4537 12053 4571 12087
rect 4571 12053 4580 12087
rect 4528 12044 4580 12053
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 8944 12087 8996 12096
rect 8944 12053 8953 12087
rect 8953 12053 8987 12087
rect 8987 12053 8996 12087
rect 8944 12044 8996 12053
rect 25044 12087 25096 12096
rect 25044 12053 25053 12087
rect 25053 12053 25087 12087
rect 25087 12053 25096 12087
rect 25044 12044 25096 12053
rect 31300 12087 31352 12096
rect 31300 12053 31309 12087
rect 31309 12053 31343 12087
rect 31343 12053 31352 12087
rect 31300 12044 31352 12053
rect 31392 12087 31444 12096
rect 31392 12053 31401 12087
rect 31401 12053 31435 12087
rect 31435 12053 31444 12087
rect 31392 12044 31444 12053
rect 9138 11942 9190 11994
rect 9202 11942 9254 11994
rect 9266 11942 9318 11994
rect 9330 11942 9382 11994
rect 9394 11942 9446 11994
rect 17326 11942 17378 11994
rect 17390 11942 17442 11994
rect 17454 11942 17506 11994
rect 17518 11942 17570 11994
rect 17582 11942 17634 11994
rect 25514 11942 25566 11994
rect 25578 11942 25630 11994
rect 25642 11942 25694 11994
rect 25706 11942 25758 11994
rect 25770 11942 25822 11994
rect 33702 11942 33754 11994
rect 33766 11942 33818 11994
rect 33830 11942 33882 11994
rect 33894 11942 33946 11994
rect 33958 11942 34010 11994
rect 4436 11840 4488 11892
rect 32036 11840 32088 11892
rect 1584 11815 1636 11824
rect 1584 11781 1593 11815
rect 1593 11781 1627 11815
rect 1627 11781 1636 11815
rect 1584 11772 1636 11781
rect 2596 11747 2648 11756
rect 2596 11713 2605 11747
rect 2605 11713 2639 11747
rect 2639 11713 2648 11747
rect 2596 11704 2648 11713
rect 2872 11747 2924 11756
rect 2872 11713 2881 11747
rect 2881 11713 2915 11747
rect 2915 11713 2924 11747
rect 2872 11704 2924 11713
rect 11152 11772 11204 11824
rect 31300 11772 31352 11824
rect 12716 11704 12768 11756
rect 19340 11747 19392 11756
rect 19340 11713 19349 11747
rect 19349 11713 19383 11747
rect 19383 11713 19392 11747
rect 19340 11704 19392 11713
rect 31668 11704 31720 11756
rect 31944 11747 31996 11756
rect 31944 11713 31953 11747
rect 31953 11713 31987 11747
rect 31987 11713 31996 11747
rect 31944 11704 31996 11713
rect 1308 11636 1360 11688
rect 31484 11679 31536 11688
rect 31484 11645 31493 11679
rect 31493 11645 31527 11679
rect 31527 11645 31536 11679
rect 31484 11636 31536 11645
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 15476 11500 15528 11552
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 5044 11398 5096 11450
rect 5108 11398 5160 11450
rect 5172 11398 5224 11450
rect 5236 11398 5288 11450
rect 5300 11398 5352 11450
rect 13232 11398 13284 11450
rect 13296 11398 13348 11450
rect 13360 11398 13412 11450
rect 13424 11398 13476 11450
rect 13488 11398 13540 11450
rect 21420 11398 21472 11450
rect 21484 11398 21536 11450
rect 21548 11398 21600 11450
rect 21612 11398 21664 11450
rect 21676 11398 21728 11450
rect 29608 11398 29660 11450
rect 29672 11398 29724 11450
rect 29736 11398 29788 11450
rect 29800 11398 29852 11450
rect 29864 11398 29916 11450
rect 3792 11296 3844 11348
rect 4528 11296 4580 11348
rect 30564 11339 30616 11348
rect 30564 11305 30573 11339
rect 30573 11305 30607 11339
rect 30607 11305 30616 11339
rect 30564 11296 30616 11305
rect 31944 11296 31996 11348
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 31392 11160 31444 11212
rect 32220 11135 32272 11144
rect 32220 11101 32229 11135
rect 32229 11101 32263 11135
rect 32263 11101 32272 11135
rect 32220 11092 32272 11101
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 31392 10999 31444 11008
rect 31392 10965 31401 10999
rect 31401 10965 31435 10999
rect 31435 10965 31444 10999
rect 31392 10956 31444 10965
rect 9138 10854 9190 10906
rect 9202 10854 9254 10906
rect 9266 10854 9318 10906
rect 9330 10854 9382 10906
rect 9394 10854 9446 10906
rect 17326 10854 17378 10906
rect 17390 10854 17442 10906
rect 17454 10854 17506 10906
rect 17518 10854 17570 10906
rect 17582 10854 17634 10906
rect 25514 10854 25566 10906
rect 25578 10854 25630 10906
rect 25642 10854 25694 10906
rect 25706 10854 25758 10906
rect 25770 10854 25822 10906
rect 33702 10854 33754 10906
rect 33766 10854 33818 10906
rect 33830 10854 33882 10906
rect 33894 10854 33946 10906
rect 33958 10854 34010 10906
rect 2872 10684 2924 10736
rect 7840 10727 7892 10736
rect 7840 10693 7849 10727
rect 7849 10693 7883 10727
rect 7883 10693 7892 10727
rect 10324 10752 10376 10804
rect 32220 10752 32272 10804
rect 7840 10684 7892 10693
rect 31668 10684 31720 10736
rect 3792 10616 3844 10668
rect 4620 10616 4672 10668
rect 4344 10480 4396 10532
rect 4804 10548 4856 10600
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 12716 10548 12768 10600
rect 2964 10455 3016 10464
rect 2964 10421 2973 10455
rect 2973 10421 3007 10455
rect 3007 10421 3016 10455
rect 2964 10412 3016 10421
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 27804 10412 27856 10464
rect 30012 10548 30064 10600
rect 30564 10616 30616 10668
rect 31392 10659 31444 10668
rect 31392 10625 31401 10659
rect 31401 10625 31435 10659
rect 31435 10625 31444 10659
rect 31392 10616 31444 10625
rect 32312 10659 32364 10668
rect 32312 10625 32321 10659
rect 32321 10625 32355 10659
rect 32355 10625 32364 10659
rect 32312 10616 32364 10625
rect 33324 10591 33376 10600
rect 33324 10557 33333 10591
rect 33333 10557 33367 10591
rect 33367 10557 33376 10591
rect 33324 10548 33376 10557
rect 31208 10455 31260 10464
rect 31208 10421 31217 10455
rect 31217 10421 31251 10455
rect 31251 10421 31260 10455
rect 31208 10412 31260 10421
rect 5044 10310 5096 10362
rect 5108 10310 5160 10362
rect 5172 10310 5224 10362
rect 5236 10310 5288 10362
rect 5300 10310 5352 10362
rect 13232 10310 13284 10362
rect 13296 10310 13348 10362
rect 13360 10310 13412 10362
rect 13424 10310 13476 10362
rect 13488 10310 13540 10362
rect 21420 10310 21472 10362
rect 21484 10310 21536 10362
rect 21548 10310 21600 10362
rect 21612 10310 21664 10362
rect 21676 10310 21728 10362
rect 29608 10310 29660 10362
rect 29672 10310 29724 10362
rect 29736 10310 29788 10362
rect 29800 10310 29852 10362
rect 29864 10310 29916 10362
rect 1768 10047 1820 10056
rect 1768 10013 1777 10047
rect 1777 10013 1811 10047
rect 1811 10013 1820 10047
rect 1768 10004 1820 10013
rect 3700 10004 3752 10056
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 7840 10208 7892 10260
rect 25872 10251 25924 10260
rect 25872 10217 25881 10251
rect 25881 10217 25915 10251
rect 25915 10217 25924 10251
rect 25872 10208 25924 10217
rect 26516 10251 26568 10260
rect 26516 10217 26525 10251
rect 26525 10217 26559 10251
rect 26559 10217 26568 10251
rect 26516 10208 26568 10217
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 30380 10072 30432 10124
rect 31668 10115 31720 10124
rect 31668 10081 31677 10115
rect 31677 10081 31711 10115
rect 31711 10081 31720 10115
rect 31668 10072 31720 10081
rect 27804 10047 27856 10056
rect 27804 10013 27813 10047
rect 27813 10013 27847 10047
rect 27847 10013 27856 10047
rect 27804 10004 27856 10013
rect 30840 10047 30892 10056
rect 30840 10013 30849 10047
rect 30849 10013 30883 10047
rect 30883 10013 30892 10047
rect 30840 10004 30892 10013
rect 31208 10004 31260 10056
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 3792 9911 3844 9920
rect 3792 9877 3801 9911
rect 3801 9877 3835 9911
rect 3835 9877 3844 9911
rect 3792 9868 3844 9877
rect 16948 9868 17000 9920
rect 31576 9911 31628 9920
rect 31576 9877 31585 9911
rect 31585 9877 31619 9911
rect 31619 9877 31628 9911
rect 31576 9868 31628 9877
rect 33048 9911 33100 9920
rect 33048 9877 33057 9911
rect 33057 9877 33091 9911
rect 33091 9877 33100 9911
rect 33048 9868 33100 9877
rect 9138 9766 9190 9818
rect 9202 9766 9254 9818
rect 9266 9766 9318 9818
rect 9330 9766 9382 9818
rect 9394 9766 9446 9818
rect 17326 9766 17378 9818
rect 17390 9766 17442 9818
rect 17454 9766 17506 9818
rect 17518 9766 17570 9818
rect 17582 9766 17634 9818
rect 25514 9766 25566 9818
rect 25578 9766 25630 9818
rect 25642 9766 25694 9818
rect 25706 9766 25758 9818
rect 25770 9766 25822 9818
rect 33702 9766 33754 9818
rect 33766 9766 33818 9818
rect 33830 9766 33882 9818
rect 33894 9766 33946 9818
rect 33958 9766 34010 9818
rect 26976 9707 27028 9716
rect 26976 9673 26985 9707
rect 26985 9673 27019 9707
rect 27019 9673 27028 9707
rect 26976 9664 27028 9673
rect 30840 9664 30892 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 32312 9596 32364 9648
rect 2596 9571 2648 9580
rect 2596 9537 2605 9571
rect 2605 9537 2639 9571
rect 2639 9537 2648 9571
rect 2596 9528 2648 9537
rect 3148 9528 3200 9580
rect 4344 9460 4396 9512
rect 24952 9571 25004 9580
rect 24952 9537 24961 9571
rect 24961 9537 24995 9571
rect 24995 9537 25004 9571
rect 24952 9528 25004 9537
rect 25044 9528 25096 9580
rect 31576 9528 31628 9580
rect 33048 9528 33100 9580
rect 15200 9503 15252 9512
rect 15200 9469 15209 9503
rect 15209 9469 15243 9503
rect 15243 9469 15252 9503
rect 15200 9460 15252 9469
rect 18880 9460 18932 9512
rect 30012 9503 30064 9512
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 3608 9324 3660 9333
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 13912 9324 13964 9376
rect 23664 9324 23716 9376
rect 27620 9324 27672 9376
rect 30012 9469 30021 9503
rect 30021 9469 30055 9503
rect 30055 9469 30064 9503
rect 30012 9460 30064 9469
rect 31116 9503 31168 9512
rect 31116 9469 31125 9503
rect 31125 9469 31159 9503
rect 31159 9469 31168 9503
rect 31116 9460 31168 9469
rect 30380 9435 30432 9444
rect 30380 9401 30389 9435
rect 30389 9401 30423 9435
rect 30423 9401 30432 9435
rect 30380 9392 30432 9401
rect 30472 9367 30524 9376
rect 30472 9333 30481 9367
rect 30481 9333 30515 9367
rect 30515 9333 30524 9367
rect 30472 9324 30524 9333
rect 30564 9367 30616 9376
rect 30564 9333 30573 9367
rect 30573 9333 30607 9367
rect 30607 9333 30616 9367
rect 30564 9324 30616 9333
rect 5044 9222 5096 9274
rect 5108 9222 5160 9274
rect 5172 9222 5224 9274
rect 5236 9222 5288 9274
rect 5300 9222 5352 9274
rect 13232 9222 13284 9274
rect 13296 9222 13348 9274
rect 13360 9222 13412 9274
rect 13424 9222 13476 9274
rect 13488 9222 13540 9274
rect 21420 9222 21472 9274
rect 21484 9222 21536 9274
rect 21548 9222 21600 9274
rect 21612 9222 21664 9274
rect 21676 9222 21728 9274
rect 29608 9222 29660 9274
rect 29672 9222 29724 9274
rect 29736 9222 29788 9274
rect 29800 9222 29852 9274
rect 29864 9222 29916 9274
rect 2596 9120 2648 9172
rect 2872 9120 2924 9172
rect 4344 9120 4396 9172
rect 9496 9120 9548 9172
rect 19708 9163 19760 9172
rect 19708 9129 19717 9163
rect 19717 9129 19751 9163
rect 19751 9129 19760 9163
rect 19708 9120 19760 9129
rect 6000 8984 6052 9036
rect 19984 8984 20036 9036
rect 3792 8916 3844 8968
rect 4344 8959 4396 8968
rect 4344 8925 4353 8959
rect 4353 8925 4387 8959
rect 4387 8925 4396 8959
rect 4344 8916 4396 8925
rect 30472 8916 30524 8968
rect 31668 9027 31720 9036
rect 31668 8993 31677 9027
rect 31677 8993 31711 9027
rect 31711 8993 31720 9027
rect 31668 8984 31720 8993
rect 31300 8916 31352 8968
rect 31576 8959 31628 8968
rect 31576 8925 31585 8959
rect 31585 8925 31619 8959
rect 31619 8925 31628 8959
rect 31576 8916 31628 8925
rect 3148 8780 3200 8832
rect 31208 8780 31260 8832
rect 9138 8678 9190 8730
rect 9202 8678 9254 8730
rect 9266 8678 9318 8730
rect 9330 8678 9382 8730
rect 9394 8678 9446 8730
rect 17326 8678 17378 8730
rect 17390 8678 17442 8730
rect 17454 8678 17506 8730
rect 17518 8678 17570 8730
rect 17582 8678 17634 8730
rect 25514 8678 25566 8730
rect 25578 8678 25630 8730
rect 25642 8678 25694 8730
rect 25706 8678 25758 8730
rect 25770 8678 25822 8730
rect 33702 8678 33754 8730
rect 33766 8678 33818 8730
rect 33830 8678 33882 8730
rect 33894 8678 33946 8730
rect 33958 8678 34010 8730
rect 3608 8576 3660 8628
rect 31116 8576 31168 8628
rect 31576 8508 31628 8560
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 4436 8415 4488 8424
rect 4436 8381 4445 8415
rect 4445 8381 4479 8415
rect 4479 8381 4488 8415
rect 4436 8372 4488 8381
rect 3976 8347 4028 8356
rect 3976 8313 3985 8347
rect 3985 8313 4019 8347
rect 4019 8313 4028 8347
rect 3976 8304 4028 8313
rect 4344 8304 4396 8356
rect 30104 8372 30156 8424
rect 31208 8415 31260 8424
rect 31208 8381 31217 8415
rect 31217 8381 31251 8415
rect 31251 8381 31260 8415
rect 31208 8372 31260 8381
rect 31300 8415 31352 8424
rect 31300 8381 31309 8415
rect 31309 8381 31343 8415
rect 31343 8381 31352 8415
rect 31300 8372 31352 8381
rect 29000 8304 29052 8356
rect 3240 8279 3292 8288
rect 3240 8245 3249 8279
rect 3249 8245 3283 8279
rect 3283 8245 3292 8279
rect 3240 8236 3292 8245
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 4804 8236 4856 8245
rect 29460 8279 29512 8288
rect 29460 8245 29469 8279
rect 29469 8245 29503 8279
rect 29503 8245 29512 8279
rect 29460 8236 29512 8245
rect 5044 8134 5096 8186
rect 5108 8134 5160 8186
rect 5172 8134 5224 8186
rect 5236 8134 5288 8186
rect 5300 8134 5352 8186
rect 13232 8134 13284 8186
rect 13296 8134 13348 8186
rect 13360 8134 13412 8186
rect 13424 8134 13476 8186
rect 13488 8134 13540 8186
rect 21420 8134 21472 8186
rect 21484 8134 21536 8186
rect 21548 8134 21600 8186
rect 21612 8134 21664 8186
rect 21676 8134 21728 8186
rect 29608 8134 29660 8186
rect 29672 8134 29724 8186
rect 29736 8134 29788 8186
rect 29800 8134 29852 8186
rect 29864 8134 29916 8186
rect 4344 8032 4396 8084
rect 32036 8032 32088 8084
rect 4712 8007 4764 8016
rect 4712 7973 4721 8007
rect 4721 7973 4755 8007
rect 4755 7973 4764 8007
rect 4712 7964 4764 7973
rect 1584 7939 1636 7948
rect 1584 7905 1593 7939
rect 1593 7905 1627 7939
rect 1627 7905 1636 7939
rect 1584 7896 1636 7905
rect 3240 7896 3292 7948
rect 4160 7896 4212 7948
rect 30564 7964 30616 8016
rect 31300 7964 31352 8016
rect 29828 7896 29880 7948
rect 31668 7939 31720 7948
rect 31668 7905 31677 7939
rect 31677 7905 31711 7939
rect 31711 7905 31720 7939
rect 31668 7896 31720 7905
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 3792 7871 3844 7880
rect 3792 7837 3801 7871
rect 3801 7837 3835 7871
rect 3835 7837 3844 7871
rect 3792 7828 3844 7837
rect 4344 7760 4396 7812
rect 4804 7760 4856 7812
rect 4436 7735 4488 7744
rect 4436 7701 4445 7735
rect 4445 7701 4479 7735
rect 4479 7701 4488 7735
rect 4436 7692 4488 7701
rect 27252 7692 27304 7744
rect 29460 7760 29512 7812
rect 9138 7590 9190 7642
rect 9202 7590 9254 7642
rect 9266 7590 9318 7642
rect 9330 7590 9382 7642
rect 9394 7590 9446 7642
rect 17326 7590 17378 7642
rect 17390 7590 17442 7642
rect 17454 7590 17506 7642
rect 17518 7590 17570 7642
rect 17582 7590 17634 7642
rect 25514 7590 25566 7642
rect 25578 7590 25630 7642
rect 25642 7590 25694 7642
rect 25706 7590 25758 7642
rect 25770 7590 25822 7642
rect 33702 7590 33754 7642
rect 33766 7590 33818 7642
rect 33830 7590 33882 7642
rect 33894 7590 33946 7642
rect 33958 7590 34010 7642
rect 1768 7488 1820 7540
rect 2596 7420 2648 7472
rect 3148 7352 3200 7404
rect 3608 7352 3660 7404
rect 4436 7488 4488 7540
rect 16948 7352 17000 7404
rect 29000 7395 29052 7404
rect 29000 7361 29009 7395
rect 29009 7361 29043 7395
rect 29043 7361 29052 7395
rect 29000 7352 29052 7361
rect 29828 7395 29880 7404
rect 29828 7361 29837 7395
rect 29837 7361 29871 7395
rect 29871 7361 29880 7395
rect 29828 7352 29880 7361
rect 31024 7352 31076 7404
rect 27344 7284 27396 7336
rect 31208 7327 31260 7336
rect 31208 7293 31217 7327
rect 31217 7293 31251 7327
rect 31251 7293 31260 7327
rect 31208 7284 31260 7293
rect 32496 7327 32548 7336
rect 32496 7293 32505 7327
rect 32505 7293 32539 7327
rect 32539 7293 32548 7327
rect 32496 7284 32548 7293
rect 2872 7191 2924 7200
rect 2872 7157 2881 7191
rect 2881 7157 2915 7191
rect 2915 7157 2924 7191
rect 2872 7148 2924 7157
rect 4436 7148 4488 7200
rect 4712 7148 4764 7200
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 27528 7148 27580 7200
rect 28356 7191 28408 7200
rect 28356 7157 28365 7191
rect 28365 7157 28399 7191
rect 28399 7157 28408 7191
rect 28356 7148 28408 7157
rect 29092 7191 29144 7200
rect 29092 7157 29101 7191
rect 29101 7157 29135 7191
rect 29135 7157 29144 7191
rect 29092 7148 29144 7157
rect 5044 7046 5096 7098
rect 5108 7046 5160 7098
rect 5172 7046 5224 7098
rect 5236 7046 5288 7098
rect 5300 7046 5352 7098
rect 13232 7046 13284 7098
rect 13296 7046 13348 7098
rect 13360 7046 13412 7098
rect 13424 7046 13476 7098
rect 13488 7046 13540 7098
rect 21420 7046 21472 7098
rect 21484 7046 21536 7098
rect 21548 7046 21600 7098
rect 21612 7046 21664 7098
rect 21676 7046 21728 7098
rect 29608 7046 29660 7098
rect 29672 7046 29724 7098
rect 29736 7046 29788 7098
rect 29800 7046 29852 7098
rect 29864 7046 29916 7098
rect 3792 6944 3844 6996
rect 26240 6876 26292 6928
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 28080 6851 28132 6860
rect 28080 6817 28089 6851
rect 28089 6817 28123 6851
rect 28123 6817 28132 6851
rect 28080 6808 28132 6817
rect 29092 6808 29144 6860
rect 33324 6851 33376 6860
rect 33324 6817 33333 6851
rect 33333 6817 33367 6851
rect 33367 6817 33376 6851
rect 33324 6808 33376 6817
rect 3976 6740 4028 6792
rect 4528 6740 4580 6792
rect 29184 6740 29236 6792
rect 27528 6715 27580 6724
rect 27528 6681 27537 6715
rect 27537 6681 27571 6715
rect 27571 6681 27580 6715
rect 27528 6672 27580 6681
rect 30564 6783 30616 6792
rect 30564 6749 30573 6783
rect 30573 6749 30607 6783
rect 30607 6749 30616 6783
rect 30564 6740 30616 6749
rect 30748 6783 30800 6792
rect 30748 6749 30757 6783
rect 30757 6749 30791 6783
rect 30791 6749 30800 6783
rect 30748 6740 30800 6749
rect 31024 6740 31076 6792
rect 32496 6740 32548 6792
rect 32588 6672 32640 6724
rect 2780 6604 2832 6656
rect 4252 6604 4304 6656
rect 27620 6647 27672 6656
rect 27620 6613 27629 6647
rect 27629 6613 27663 6647
rect 27663 6613 27672 6647
rect 27620 6604 27672 6613
rect 30472 6604 30524 6656
rect 9138 6502 9190 6554
rect 9202 6502 9254 6554
rect 9266 6502 9318 6554
rect 9330 6502 9382 6554
rect 9394 6502 9446 6554
rect 17326 6502 17378 6554
rect 17390 6502 17442 6554
rect 17454 6502 17506 6554
rect 17518 6502 17570 6554
rect 17582 6502 17634 6554
rect 25514 6502 25566 6554
rect 25578 6502 25630 6554
rect 25642 6502 25694 6554
rect 25706 6502 25758 6554
rect 25770 6502 25822 6554
rect 33702 6502 33754 6554
rect 33766 6502 33818 6554
rect 33830 6502 33882 6554
rect 33894 6502 33946 6554
rect 33958 6502 34010 6554
rect 4712 6443 4764 6452
rect 4712 6409 4721 6443
rect 4721 6409 4755 6443
rect 4755 6409 4764 6443
rect 4712 6400 4764 6409
rect 25228 6400 25280 6452
rect 27252 6443 27304 6452
rect 27252 6409 27261 6443
rect 27261 6409 27295 6443
rect 27295 6409 27304 6443
rect 27252 6400 27304 6409
rect 30748 6400 30800 6452
rect 4160 6332 4212 6384
rect 27620 6332 27672 6384
rect 30564 6332 30616 6384
rect 32036 6332 32088 6384
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 30932 6264 30984 6316
rect 31668 6264 31720 6316
rect 31944 6307 31996 6316
rect 31944 6273 31953 6307
rect 31953 6273 31987 6307
rect 31987 6273 31996 6307
rect 31944 6264 31996 6273
rect 4344 6196 4396 6248
rect 1308 6060 1360 6112
rect 9864 6171 9916 6180
rect 9864 6137 9873 6171
rect 9873 6137 9907 6171
rect 9907 6137 9916 6171
rect 9864 6128 9916 6137
rect 27620 6239 27672 6248
rect 27620 6205 27629 6239
rect 27629 6205 27663 6239
rect 27663 6205 27672 6239
rect 27620 6196 27672 6205
rect 28816 6196 28868 6248
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 10232 6060 10284 6112
rect 10416 6103 10468 6112
rect 10416 6069 10425 6103
rect 10425 6069 10459 6103
rect 10459 6069 10468 6103
rect 10416 6060 10468 6069
rect 29092 6060 29144 6112
rect 31484 6239 31536 6248
rect 31484 6205 31493 6239
rect 31493 6205 31527 6239
rect 31527 6205 31536 6239
rect 31484 6196 31536 6205
rect 32128 6239 32180 6248
rect 32128 6205 32137 6239
rect 32137 6205 32171 6239
rect 32171 6205 32180 6239
rect 32128 6196 32180 6205
rect 34060 6060 34112 6112
rect 5044 5958 5096 6010
rect 5108 5958 5160 6010
rect 5172 5958 5224 6010
rect 5236 5958 5288 6010
rect 5300 5958 5352 6010
rect 13232 5958 13284 6010
rect 13296 5958 13348 6010
rect 13360 5958 13412 6010
rect 13424 5958 13476 6010
rect 13488 5958 13540 6010
rect 21420 5958 21472 6010
rect 21484 5958 21536 6010
rect 21548 5958 21600 6010
rect 21612 5958 21664 6010
rect 21676 5958 21728 6010
rect 29608 5958 29660 6010
rect 29672 5958 29724 6010
rect 29736 5958 29788 6010
rect 29800 5958 29852 6010
rect 29864 5958 29916 6010
rect 4344 5856 4396 5908
rect 4528 5856 4580 5908
rect 15200 5856 15252 5908
rect 26148 5856 26200 5908
rect 26516 5856 26568 5908
rect 27344 5899 27396 5908
rect 27344 5865 27353 5899
rect 27353 5865 27387 5899
rect 27387 5865 27396 5899
rect 27344 5856 27396 5865
rect 27620 5856 27672 5908
rect 11704 5831 11756 5840
rect 11704 5797 11713 5831
rect 11713 5797 11747 5831
rect 11747 5797 11756 5831
rect 11704 5788 11756 5797
rect 25228 5831 25280 5840
rect 25228 5797 25237 5831
rect 25237 5797 25271 5831
rect 25271 5797 25280 5831
rect 25228 5788 25280 5797
rect 31760 5856 31812 5908
rect 29092 5831 29144 5840
rect 29092 5797 29101 5831
rect 29101 5797 29135 5831
rect 29135 5797 29144 5831
rect 29092 5788 29144 5797
rect 30380 5788 30432 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 2872 5763 2924 5772
rect 2872 5729 2881 5763
rect 2881 5729 2915 5763
rect 2915 5729 2924 5763
rect 2872 5720 2924 5729
rect 8852 5720 8904 5772
rect 26792 5720 26844 5772
rect 28356 5720 28408 5772
rect 29460 5720 29512 5772
rect 30472 5763 30524 5772
rect 30472 5729 30481 5763
rect 30481 5729 30515 5763
rect 30515 5729 30524 5763
rect 30472 5720 30524 5729
rect 2596 5695 2648 5704
rect 2596 5661 2605 5695
rect 2605 5661 2639 5695
rect 2639 5661 2648 5695
rect 2596 5652 2648 5661
rect 3516 5652 3568 5704
rect 10048 5695 10100 5704
rect 10048 5661 10057 5695
rect 10057 5661 10091 5695
rect 10091 5661 10100 5695
rect 10048 5652 10100 5661
rect 10692 5652 10744 5704
rect 26700 5695 26752 5704
rect 26700 5661 26709 5695
rect 26709 5661 26743 5695
rect 26743 5661 26752 5695
rect 26700 5652 26752 5661
rect 8760 5627 8812 5636
rect 8760 5593 8769 5627
rect 8769 5593 8803 5627
rect 8803 5593 8812 5627
rect 8760 5584 8812 5593
rect 10416 5584 10468 5636
rect 28172 5695 28224 5704
rect 28172 5661 28181 5695
rect 28181 5661 28215 5695
rect 28215 5661 28224 5695
rect 28172 5652 28224 5661
rect 31116 5652 31168 5704
rect 31944 5720 31996 5772
rect 32036 5695 32088 5704
rect 32036 5661 32045 5695
rect 32045 5661 32079 5695
rect 32079 5661 32088 5695
rect 32036 5652 32088 5661
rect 32864 5695 32916 5704
rect 32864 5661 32873 5695
rect 32873 5661 32907 5695
rect 32907 5661 32916 5695
rect 32864 5652 32916 5661
rect 9036 5516 9088 5568
rect 29276 5584 29328 5636
rect 31576 5584 31628 5636
rect 12532 5516 12584 5568
rect 13728 5516 13780 5568
rect 28908 5559 28960 5568
rect 28908 5525 28917 5559
rect 28917 5525 28951 5559
rect 28951 5525 28960 5559
rect 28908 5516 28960 5525
rect 29920 5559 29972 5568
rect 29920 5525 29929 5559
rect 29929 5525 29963 5559
rect 29963 5525 29972 5559
rect 29920 5516 29972 5525
rect 9138 5414 9190 5466
rect 9202 5414 9254 5466
rect 9266 5414 9318 5466
rect 9330 5414 9382 5466
rect 9394 5414 9446 5466
rect 17326 5414 17378 5466
rect 17390 5414 17442 5466
rect 17454 5414 17506 5466
rect 17518 5414 17570 5466
rect 17582 5414 17634 5466
rect 25514 5414 25566 5466
rect 25578 5414 25630 5466
rect 25642 5414 25694 5466
rect 25706 5414 25758 5466
rect 25770 5414 25822 5466
rect 33702 5414 33754 5466
rect 33766 5414 33818 5466
rect 33830 5414 33882 5466
rect 33894 5414 33946 5466
rect 33958 5414 34010 5466
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 3608 5355 3660 5364
rect 3608 5321 3617 5355
rect 3617 5321 3651 5355
rect 3651 5321 3660 5355
rect 3608 5312 3660 5321
rect 10048 5355 10100 5364
rect 10048 5321 10057 5355
rect 10057 5321 10091 5355
rect 10091 5321 10100 5355
rect 10048 5312 10100 5321
rect 11704 5312 11756 5364
rect 12348 5355 12400 5364
rect 12348 5321 12357 5355
rect 12357 5321 12391 5355
rect 12391 5321 12400 5355
rect 12348 5312 12400 5321
rect 26056 5355 26108 5364
rect 26056 5321 26065 5355
rect 26065 5321 26099 5355
rect 26099 5321 26108 5355
rect 26056 5312 26108 5321
rect 30104 5355 30156 5364
rect 30104 5321 30113 5355
rect 30113 5321 30147 5355
rect 30147 5321 30156 5355
rect 30104 5312 30156 5321
rect 33508 5355 33560 5364
rect 33508 5321 33517 5355
rect 33517 5321 33551 5355
rect 33551 5321 33560 5355
rect 33508 5312 33560 5321
rect 2596 5244 2648 5296
rect 8392 5244 8444 5296
rect 8760 5244 8812 5296
rect 13636 5244 13688 5296
rect 15936 5287 15988 5296
rect 15936 5253 15945 5287
rect 15945 5253 15979 5287
rect 15979 5253 15988 5287
rect 15936 5244 15988 5253
rect 23388 5287 23440 5296
rect 23388 5253 23397 5287
rect 23397 5253 23431 5287
rect 23431 5253 23440 5287
rect 23388 5244 23440 5253
rect 25228 5244 25280 5296
rect 27068 5244 27120 5296
rect 29092 5244 29144 5296
rect 29184 5244 29236 5296
rect 2780 5176 2832 5228
rect 3148 5176 3200 5228
rect 4436 5176 4488 5228
rect 4528 5040 4580 5092
rect 9772 5176 9824 5228
rect 13728 5176 13780 5228
rect 16764 5219 16816 5228
rect 16764 5185 16773 5219
rect 16773 5185 16807 5219
rect 16807 5185 16816 5219
rect 16764 5176 16816 5185
rect 24308 5176 24360 5228
rect 26240 5219 26292 5228
rect 26240 5185 26249 5219
rect 26249 5185 26283 5219
rect 26283 5185 26292 5219
rect 26240 5176 26292 5185
rect 28816 5176 28868 5228
rect 31944 5176 31996 5228
rect 32128 5219 32180 5228
rect 32128 5185 32137 5219
rect 32137 5185 32171 5219
rect 32171 5185 32180 5219
rect 32128 5176 32180 5185
rect 8300 5108 8352 5160
rect 9036 5108 9088 5160
rect 10508 5108 10560 5160
rect 10784 5151 10836 5160
rect 10784 5117 10793 5151
rect 10793 5117 10827 5151
rect 10827 5117 10836 5151
rect 10784 5108 10836 5117
rect 12072 5151 12124 5160
rect 12072 5117 12081 5151
rect 12081 5117 12115 5151
rect 12115 5117 12124 5151
rect 12072 5108 12124 5117
rect 12440 5108 12492 5160
rect 16580 5108 16632 5160
rect 8484 5040 8536 5092
rect 24584 5151 24636 5160
rect 24584 5117 24593 5151
rect 24593 5117 24627 5151
rect 24627 5117 24636 5151
rect 24584 5108 24636 5117
rect 26976 5151 27028 5160
rect 26976 5117 26985 5151
rect 26985 5117 27019 5151
rect 27019 5117 27028 5151
rect 26976 5108 27028 5117
rect 28724 5151 28776 5160
rect 28724 5117 28733 5151
rect 28733 5117 28767 5151
rect 28767 5117 28776 5151
rect 28724 5108 28776 5117
rect 30104 5108 30156 5160
rect 4436 5015 4488 5024
rect 4436 4981 4445 5015
rect 4445 4981 4479 5015
rect 4479 4981 4488 5015
rect 4436 4972 4488 4981
rect 8576 5015 8628 5024
rect 8576 4981 8585 5015
rect 8585 4981 8619 5015
rect 8619 4981 8628 5015
rect 8576 4972 8628 4981
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 8760 4972 8812 5024
rect 9864 4972 9916 5024
rect 19340 4972 19392 5024
rect 24032 5015 24084 5024
rect 24032 4981 24041 5015
rect 24041 4981 24075 5015
rect 24075 4981 24084 5015
rect 24032 4972 24084 4981
rect 26608 4972 26660 5024
rect 27712 5015 27764 5024
rect 27712 4981 27721 5015
rect 27721 4981 27755 5015
rect 27755 4981 27764 5015
rect 27712 4972 27764 4981
rect 30012 5040 30064 5092
rect 5044 4870 5096 4922
rect 5108 4870 5160 4922
rect 5172 4870 5224 4922
rect 5236 4870 5288 4922
rect 5300 4870 5352 4922
rect 13232 4870 13284 4922
rect 13296 4870 13348 4922
rect 13360 4870 13412 4922
rect 13424 4870 13476 4922
rect 13488 4870 13540 4922
rect 21420 4870 21472 4922
rect 21484 4870 21536 4922
rect 21548 4870 21600 4922
rect 21612 4870 21664 4922
rect 21676 4870 21728 4922
rect 29608 4870 29660 4922
rect 29672 4870 29724 4922
rect 29736 4870 29788 4922
rect 29800 4870 29852 4922
rect 29864 4870 29916 4922
rect 4436 4768 4488 4820
rect 3240 4632 3292 4684
rect 4252 4564 4304 4616
rect 8484 4768 8536 4820
rect 8576 4768 8628 4820
rect 8760 4811 8812 4820
rect 8760 4777 8769 4811
rect 8769 4777 8803 4811
rect 8803 4777 8812 4811
rect 8760 4768 8812 4777
rect 8300 4700 8352 4752
rect 8392 4564 8444 4616
rect 9496 4768 9548 4820
rect 10508 4811 10560 4820
rect 10508 4777 10517 4811
rect 10517 4777 10551 4811
rect 10551 4777 10560 4811
rect 10508 4768 10560 4777
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 13728 4768 13780 4820
rect 24032 4768 24084 4820
rect 24584 4768 24636 4820
rect 11520 4632 11572 4684
rect 12348 4675 12400 4684
rect 12348 4641 12357 4675
rect 12357 4641 12391 4675
rect 12391 4641 12400 4675
rect 12348 4632 12400 4641
rect 14372 4743 14424 4752
rect 14372 4709 14381 4743
rect 14381 4709 14415 4743
rect 14415 4709 14424 4743
rect 14372 4700 14424 4709
rect 18696 4700 18748 4752
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 13820 4564 13872 4616
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 23388 4632 23440 4684
rect 16672 4564 16724 4616
rect 26424 4768 26476 4820
rect 26792 4768 26844 4820
rect 29092 4768 29144 4820
rect 30748 4768 30800 4820
rect 26516 4632 26568 4684
rect 27712 4632 27764 4684
rect 28908 4675 28960 4684
rect 28908 4641 28917 4675
rect 28917 4641 28951 4675
rect 28951 4641 28960 4675
rect 28908 4632 28960 4641
rect 30932 4675 30984 4684
rect 30932 4641 30941 4675
rect 30941 4641 30975 4675
rect 30975 4641 30984 4675
rect 30932 4632 30984 4641
rect 32036 4632 32088 4684
rect 24952 4607 25004 4616
rect 24952 4573 24961 4607
rect 24961 4573 24995 4607
rect 24995 4573 25004 4607
rect 24952 4564 25004 4573
rect 24860 4496 24912 4548
rect 25412 4564 25464 4616
rect 27528 4496 27580 4548
rect 27896 4539 27948 4548
rect 27896 4505 27905 4539
rect 27905 4505 27939 4539
rect 27939 4505 27948 4539
rect 27896 4496 27948 4505
rect 29552 4607 29604 4616
rect 29552 4573 29561 4607
rect 29561 4573 29595 4607
rect 29595 4573 29604 4607
rect 29552 4564 29604 4573
rect 29736 4564 29788 4616
rect 32220 4607 32272 4616
rect 32220 4573 32229 4607
rect 32229 4573 32263 4607
rect 32263 4573 32272 4607
rect 32220 4564 32272 4573
rect 31668 4496 31720 4548
rect 31852 4539 31904 4548
rect 31852 4505 31861 4539
rect 31861 4505 31895 4539
rect 31895 4505 31904 4539
rect 31852 4496 31904 4505
rect 9588 4428 9640 4480
rect 12992 4471 13044 4480
rect 12992 4437 13001 4471
rect 13001 4437 13035 4471
rect 13035 4437 13044 4471
rect 12992 4428 13044 4437
rect 13636 4428 13688 4480
rect 14464 4428 14516 4480
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 15476 4471 15528 4480
rect 15476 4437 15485 4471
rect 15485 4437 15519 4471
rect 15519 4437 15528 4471
rect 15476 4428 15528 4437
rect 16764 4471 16816 4480
rect 16764 4437 16773 4471
rect 16773 4437 16807 4471
rect 16807 4437 16816 4471
rect 16764 4428 16816 4437
rect 16856 4471 16908 4480
rect 16856 4437 16865 4471
rect 16865 4437 16899 4471
rect 16899 4437 16908 4471
rect 16856 4428 16908 4437
rect 22744 4471 22796 4480
rect 22744 4437 22753 4471
rect 22753 4437 22787 4471
rect 22787 4437 22796 4471
rect 22744 4428 22796 4437
rect 24216 4471 24268 4480
rect 24216 4437 24225 4471
rect 24225 4437 24259 4471
rect 24259 4437 24268 4471
rect 24216 4428 24268 4437
rect 26056 4428 26108 4480
rect 27344 4471 27396 4480
rect 27344 4437 27353 4471
rect 27353 4437 27387 4471
rect 27387 4437 27396 4471
rect 27344 4428 27396 4437
rect 27804 4428 27856 4480
rect 30196 4471 30248 4480
rect 30196 4437 30205 4471
rect 30205 4437 30239 4471
rect 30239 4437 30248 4471
rect 30196 4428 30248 4437
rect 9138 4326 9190 4378
rect 9202 4326 9254 4378
rect 9266 4326 9318 4378
rect 9330 4326 9382 4378
rect 9394 4326 9446 4378
rect 17326 4326 17378 4378
rect 17390 4326 17442 4378
rect 17454 4326 17506 4378
rect 17518 4326 17570 4378
rect 17582 4326 17634 4378
rect 25514 4326 25566 4378
rect 25578 4326 25630 4378
rect 25642 4326 25694 4378
rect 25706 4326 25758 4378
rect 25770 4326 25822 4378
rect 33702 4326 33754 4378
rect 33766 4326 33818 4378
rect 33830 4326 33882 4378
rect 33894 4326 33946 4378
rect 33958 4326 34010 4378
rect 9496 4224 9548 4276
rect 10784 4224 10836 4276
rect 12532 4224 12584 4276
rect 13820 4267 13872 4276
rect 13820 4233 13829 4267
rect 13829 4233 13863 4267
rect 13863 4233 13872 4267
rect 13820 4224 13872 4233
rect 24952 4224 25004 4276
rect 28172 4224 28224 4276
rect 29276 4224 29328 4276
rect 2964 4088 3016 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 9588 4131 9640 4140
rect 9588 4097 9622 4131
rect 9622 4097 9640 4131
rect 9588 4088 9640 4097
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 15384 4088 15436 4140
rect 16764 4131 16816 4140
rect 16764 4097 16773 4131
rect 16773 4097 16807 4131
rect 16807 4097 16816 4131
rect 16764 4088 16816 4097
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 24400 4088 24452 4140
rect 24584 4088 24636 4140
rect 26884 4088 26936 4140
rect 6736 4020 6788 4072
rect 7748 4020 7800 4072
rect 12624 4063 12676 4072
rect 12624 4029 12633 4063
rect 12633 4029 12667 4063
rect 12667 4029 12676 4063
rect 12624 4020 12676 4029
rect 13084 4020 13136 4072
rect 14096 4063 14148 4072
rect 14096 4029 14105 4063
rect 14105 4029 14139 4063
rect 14139 4029 14148 4063
rect 14096 4020 14148 4029
rect 16028 4063 16080 4072
rect 16028 4029 16037 4063
rect 16037 4029 16071 4063
rect 16071 4029 16080 4063
rect 16028 4020 16080 4029
rect 17040 4063 17092 4072
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 17040 4020 17092 4029
rect 19524 4063 19576 4072
rect 19524 4029 19533 4063
rect 19533 4029 19567 4063
rect 19567 4029 19576 4063
rect 19524 4020 19576 4029
rect 23204 4020 23256 4072
rect 13636 3952 13688 4004
rect 24768 4020 24820 4072
rect 26332 4020 26384 4072
rect 28724 4088 28776 4140
rect 29000 4131 29052 4140
rect 29000 4097 29018 4131
rect 29018 4097 29052 4131
rect 29000 4088 29052 4097
rect 30840 4088 30892 4140
rect 31760 4156 31812 4208
rect 32128 4088 32180 4140
rect 2596 3884 2648 3936
rect 6644 3884 6696 3936
rect 11336 3927 11388 3936
rect 11336 3893 11345 3927
rect 11345 3893 11379 3927
rect 11379 3893 11388 3927
rect 11336 3884 11388 3893
rect 14648 3927 14700 3936
rect 14648 3893 14657 3927
rect 14657 3893 14691 3927
rect 14691 3893 14700 3927
rect 14648 3884 14700 3893
rect 18144 3927 18196 3936
rect 18144 3893 18153 3927
rect 18153 3893 18187 3927
rect 18187 3893 18196 3927
rect 18144 3884 18196 3893
rect 23296 3927 23348 3936
rect 23296 3893 23305 3927
rect 23305 3893 23339 3927
rect 23339 3893 23348 3927
rect 23296 3884 23348 3893
rect 23388 3884 23440 3936
rect 26516 3995 26568 4004
rect 26516 3961 26525 3995
rect 26525 3961 26559 3995
rect 26559 3961 26568 3995
rect 26516 3952 26568 3961
rect 27160 4020 27212 4072
rect 27896 4020 27948 4072
rect 31116 4020 31168 4072
rect 31668 4020 31720 4072
rect 26240 3884 26292 3936
rect 27068 3884 27120 3936
rect 27620 3927 27672 3936
rect 27620 3893 27629 3927
rect 27629 3893 27663 3927
rect 27663 3893 27672 3927
rect 27620 3884 27672 3893
rect 29552 3884 29604 3936
rect 5044 3782 5096 3834
rect 5108 3782 5160 3834
rect 5172 3782 5224 3834
rect 5236 3782 5288 3834
rect 5300 3782 5352 3834
rect 13232 3782 13284 3834
rect 13296 3782 13348 3834
rect 13360 3782 13412 3834
rect 13424 3782 13476 3834
rect 13488 3782 13540 3834
rect 21420 3782 21472 3834
rect 21484 3782 21536 3834
rect 21548 3782 21600 3834
rect 21612 3782 21664 3834
rect 21676 3782 21728 3834
rect 29608 3782 29660 3834
rect 29672 3782 29724 3834
rect 29736 3782 29788 3834
rect 29800 3782 29852 3834
rect 29864 3782 29916 3834
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 6644 3587 6696 3596
rect 6644 3553 6653 3587
rect 6653 3553 6687 3587
rect 6687 3553 6696 3587
rect 6644 3544 6696 3553
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 8944 3680 8996 3732
rect 11520 3723 11572 3732
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 13912 3680 13964 3732
rect 14096 3723 14148 3732
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 19524 3680 19576 3732
rect 9496 3544 9548 3596
rect 8668 3519 8720 3528
rect 8668 3485 8677 3519
rect 8677 3485 8711 3519
rect 8711 3485 8720 3519
rect 8668 3476 8720 3485
rect 9864 3476 9916 3528
rect 13636 3587 13688 3596
rect 13636 3553 13645 3587
rect 13645 3553 13679 3587
rect 13679 3553 13688 3587
rect 13636 3544 13688 3553
rect 16580 3544 16632 3596
rect 23388 3680 23440 3732
rect 24308 3680 24360 3732
rect 24400 3723 24452 3732
rect 24400 3689 24409 3723
rect 24409 3689 24443 3723
rect 24443 3689 24452 3723
rect 24400 3680 24452 3689
rect 24584 3680 24636 3732
rect 24860 3680 24912 3732
rect 25412 3680 25464 3732
rect 27344 3680 27396 3732
rect 31852 3680 31904 3732
rect 32864 3723 32916 3732
rect 32864 3689 32873 3723
rect 32873 3689 32907 3723
rect 32907 3689 32916 3723
rect 32864 3680 32916 3689
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 8300 3451 8352 3460
rect 8300 3417 8309 3451
rect 8309 3417 8343 3451
rect 8343 3417 8352 3451
rect 8300 3408 8352 3417
rect 10232 3408 10284 3460
rect 11336 3408 11388 3460
rect 22192 3587 22244 3596
rect 22192 3553 22201 3587
rect 22201 3553 22235 3587
rect 22235 3553 22244 3587
rect 22192 3544 22244 3553
rect 20352 3519 20404 3528
rect 20352 3485 20361 3519
rect 20361 3485 20395 3519
rect 20395 3485 20404 3519
rect 20352 3476 20404 3485
rect 22744 3476 22796 3528
rect 22928 3476 22980 3528
rect 24768 3476 24820 3528
rect 16856 3408 16908 3460
rect 21916 3408 21968 3460
rect 23388 3408 23440 3460
rect 25320 3476 25372 3528
rect 26240 3476 26292 3528
rect 26332 3519 26384 3528
rect 26332 3485 26341 3519
rect 26341 3485 26375 3519
rect 26375 3485 26384 3519
rect 26332 3476 26384 3485
rect 26424 3519 26476 3528
rect 26424 3485 26433 3519
rect 26433 3485 26467 3519
rect 26467 3485 26476 3519
rect 26424 3476 26476 3485
rect 6000 3340 6052 3392
rect 8116 3340 8168 3392
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 12900 3340 12952 3392
rect 15476 3340 15528 3392
rect 16948 3383 17000 3392
rect 16948 3349 16957 3383
rect 16957 3349 16991 3383
rect 16991 3349 17000 3383
rect 16948 3340 17000 3349
rect 24124 3383 24176 3392
rect 24124 3349 24133 3383
rect 24133 3349 24167 3383
rect 24167 3349 24176 3383
rect 24124 3340 24176 3349
rect 24492 3340 24544 3392
rect 30012 3612 30064 3664
rect 29920 3476 29972 3528
rect 30196 3519 30248 3528
rect 30196 3485 30205 3519
rect 30205 3485 30239 3519
rect 30239 3485 30248 3519
rect 30196 3476 30248 3485
rect 31760 3519 31812 3528
rect 31760 3485 31769 3519
rect 31769 3485 31803 3519
rect 31803 3485 31812 3519
rect 31760 3476 31812 3485
rect 31944 3476 31996 3528
rect 31116 3408 31168 3460
rect 27896 3340 27948 3392
rect 31852 3340 31904 3392
rect 33508 3340 33560 3392
rect 9138 3238 9190 3290
rect 9202 3238 9254 3290
rect 9266 3238 9318 3290
rect 9330 3238 9382 3290
rect 9394 3238 9446 3290
rect 17326 3238 17378 3290
rect 17390 3238 17442 3290
rect 17454 3238 17506 3290
rect 17518 3238 17570 3290
rect 17582 3238 17634 3290
rect 25514 3238 25566 3290
rect 25578 3238 25630 3290
rect 25642 3238 25694 3290
rect 25706 3238 25758 3290
rect 25770 3238 25822 3290
rect 33702 3238 33754 3290
rect 33766 3238 33818 3290
rect 33830 3238 33882 3290
rect 33894 3238 33946 3290
rect 33958 3238 34010 3290
rect 8300 3136 8352 3188
rect 11428 3136 11480 3188
rect 12900 3136 12952 3188
rect 12992 3136 13044 3188
rect 13084 3136 13136 3188
rect 16028 3136 16080 3188
rect 16672 3179 16724 3188
rect 16672 3145 16681 3179
rect 16681 3145 16715 3179
rect 16715 3145 16724 3179
rect 16672 3136 16724 3145
rect 18144 3136 18196 3188
rect 22192 3136 22244 3188
rect 23204 3136 23256 3188
rect 3424 3000 3476 3052
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 8760 3043 8812 3052
rect 8760 3009 8794 3043
rect 8794 3009 8812 3043
rect 8760 3000 8812 3009
rect 9496 3000 9548 3052
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 14464 3000 14516 3052
rect 19708 3043 19760 3052
rect 19708 3009 19717 3043
rect 19717 3009 19751 3043
rect 19751 3009 19760 3043
rect 19708 3000 19760 3009
rect 2596 2932 2648 2984
rect 4988 2975 5040 2984
rect 4988 2941 4997 2975
rect 4997 2941 5031 2975
rect 5031 2941 5040 2975
rect 4988 2932 5040 2941
rect 10508 2975 10560 2984
rect 10508 2941 10517 2975
rect 10517 2941 10551 2975
rect 10551 2941 10560 2975
rect 10508 2932 10560 2941
rect 12532 2975 12584 2984
rect 12532 2941 12541 2975
rect 12541 2941 12575 2975
rect 12575 2941 12584 2975
rect 12532 2932 12584 2941
rect 14832 2932 14884 2984
rect 17316 2975 17368 2984
rect 17316 2941 17325 2975
rect 17325 2941 17359 2975
rect 17359 2941 17368 2975
rect 17316 2932 17368 2941
rect 17684 2975 17736 2984
rect 17684 2941 17693 2975
rect 17693 2941 17727 2975
rect 17727 2941 17736 2975
rect 17684 2932 17736 2941
rect 18788 2932 18840 2984
rect 23664 3000 23716 3052
rect 21824 2864 21876 2916
rect 24124 3136 24176 3188
rect 26976 3179 27028 3188
rect 26976 3145 26985 3179
rect 26985 3145 27019 3179
rect 27019 3145 27028 3179
rect 26976 3136 27028 3145
rect 30840 3136 30892 3188
rect 32588 3136 32640 3188
rect 26332 3068 26384 3120
rect 27068 3000 27120 3052
rect 27804 3000 27856 3052
rect 26332 2975 26384 2984
rect 26332 2941 26341 2975
rect 26341 2941 26375 2975
rect 26375 2941 26384 2975
rect 31852 3111 31904 3120
rect 31852 3077 31861 3111
rect 31861 3077 31895 3111
rect 31895 3077 31904 3111
rect 31852 3068 31904 3077
rect 26332 2932 26384 2941
rect 28356 2975 28408 2984
rect 28356 2941 28365 2975
rect 28365 2941 28399 2975
rect 28399 2941 28408 2975
rect 28356 2932 28408 2941
rect 28632 2975 28684 2984
rect 28632 2941 28641 2975
rect 28641 2941 28675 2975
rect 28675 2941 28684 2975
rect 28632 2932 28684 2941
rect 29920 3043 29972 3052
rect 29920 3009 29929 3043
rect 29929 3009 29963 3043
rect 29963 3009 29972 3043
rect 29920 3000 29972 3009
rect 32128 3043 32180 3052
rect 32128 3009 32137 3043
rect 32137 3009 32171 3043
rect 32171 3009 32180 3043
rect 32128 3000 32180 3009
rect 30012 2932 30064 2984
rect 30196 2932 30248 2984
rect 26700 2907 26752 2916
rect 26700 2873 26709 2907
rect 26709 2873 26743 2907
rect 26743 2873 26752 2907
rect 26700 2864 26752 2873
rect 28816 2864 28868 2916
rect 9128 2796 9180 2848
rect 5044 2694 5096 2746
rect 5108 2694 5160 2746
rect 5172 2694 5224 2746
rect 5236 2694 5288 2746
rect 5300 2694 5352 2746
rect 13232 2694 13284 2746
rect 13296 2694 13348 2746
rect 13360 2694 13412 2746
rect 13424 2694 13476 2746
rect 13488 2694 13540 2746
rect 21420 2694 21472 2746
rect 21484 2694 21536 2746
rect 21548 2694 21600 2746
rect 21612 2694 21664 2746
rect 21676 2694 21728 2746
rect 29608 2694 29660 2746
rect 29672 2694 29724 2746
rect 29736 2694 29788 2746
rect 29800 2694 29852 2746
rect 29864 2694 29916 2746
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12440 2592 12492 2601
rect 14372 2635 14424 2644
rect 14372 2601 14381 2635
rect 14381 2601 14415 2635
rect 14415 2601 14424 2635
rect 14372 2592 14424 2601
rect 17316 2635 17368 2644
rect 17316 2601 17325 2635
rect 17325 2601 17359 2635
rect 17359 2601 17368 2635
rect 17316 2592 17368 2601
rect 19064 2592 19116 2644
rect 29552 2592 29604 2644
rect 31760 2592 31812 2644
rect 2504 2524 2556 2576
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 7840 2456 7892 2508
rect 9956 2456 10008 2508
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 848 2320 900 2372
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 8116 2388 8168 2440
rect 9772 2431 9824 2440
rect 9772 2397 9781 2431
rect 9781 2397 9815 2431
rect 9815 2397 9824 2431
rect 9772 2388 9824 2397
rect 11612 2456 11664 2508
rect 13268 2499 13320 2508
rect 13268 2465 13277 2499
rect 13277 2465 13311 2499
rect 13311 2465 13320 2499
rect 13268 2456 13320 2465
rect 14648 2456 14700 2508
rect 16028 2499 16080 2508
rect 16028 2465 16037 2499
rect 16037 2465 16071 2499
rect 16071 2465 16080 2499
rect 16028 2456 16080 2465
rect 16948 2456 17000 2508
rect 17960 2456 18012 2508
rect 19708 2499 19760 2508
rect 19708 2465 19717 2499
rect 19717 2465 19751 2499
rect 19751 2465 19760 2499
rect 19708 2456 19760 2465
rect 11888 2388 11940 2440
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 12624 2388 12676 2440
rect 17040 2388 17092 2440
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 19340 2431 19392 2440
rect 19340 2397 19349 2431
rect 19349 2397 19383 2431
rect 19383 2397 19392 2431
rect 19340 2388 19392 2397
rect 22008 2456 22060 2508
rect 23296 2499 23348 2508
rect 23296 2465 23305 2499
rect 23305 2465 23339 2499
rect 23339 2465 23348 2499
rect 23296 2456 23348 2465
rect 24952 2524 25004 2576
rect 25320 2524 25372 2576
rect 26332 2524 26384 2576
rect 26424 2524 26476 2576
rect 27620 2524 27672 2576
rect 28356 2524 28408 2576
rect 26884 2456 26936 2508
rect 27528 2456 27580 2508
rect 21916 2431 21968 2440
rect 21916 2397 21925 2431
rect 21925 2397 21959 2431
rect 21959 2397 21968 2431
rect 21916 2388 21968 2397
rect 23848 2388 23900 2440
rect 24216 2388 24268 2440
rect 24676 2388 24728 2440
rect 26056 2388 26108 2440
rect 26608 2388 26660 2440
rect 30012 2499 30064 2508
rect 30012 2465 30021 2499
rect 30021 2465 30055 2499
rect 30055 2465 30064 2499
rect 30012 2456 30064 2465
rect 26792 2320 26844 2372
rect 27160 2320 27212 2372
rect 28540 2320 28592 2372
rect 30472 2388 30524 2440
rect 31116 2388 31168 2440
rect 23388 2252 23440 2304
rect 28908 2252 28960 2304
rect 32588 2252 32640 2304
rect 9138 2150 9190 2202
rect 9202 2150 9254 2202
rect 9266 2150 9318 2202
rect 9330 2150 9382 2202
rect 9394 2150 9446 2202
rect 17326 2150 17378 2202
rect 17390 2150 17442 2202
rect 17454 2150 17506 2202
rect 17518 2150 17570 2202
rect 17582 2150 17634 2202
rect 25514 2150 25566 2202
rect 25578 2150 25630 2202
rect 25642 2150 25694 2202
rect 25706 2150 25758 2202
rect 25770 2150 25822 2202
rect 33702 2150 33754 2202
rect 33766 2150 33818 2202
rect 33830 2150 33882 2202
rect 33894 2150 33946 2202
rect 33958 2150 34010 2202
rect 23848 2048 23900 2100
rect 28080 2048 28132 2100
rect 27068 1504 27120 1556
rect 30196 1504 30248 1556
rect 25688 1436 25740 1488
rect 28632 1436 28684 1488
rect 20352 1368 20404 1420
rect 22008 1368 22060 1420
<< metal2 >>
rect 1030 34200 1086 35000
rect 2594 34354 2650 35000
rect 2516 34326 2650 34354
rect 1044 30190 1072 34200
rect 1584 32360 1636 32366
rect 1584 32302 1636 32308
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 30297 1440 31758
rect 1596 31482 1624 32302
rect 2136 32224 2188 32230
rect 2136 32166 2188 32172
rect 2148 32026 2176 32166
rect 2136 32020 2188 32026
rect 2136 31962 2188 31968
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1768 31272 1820 31278
rect 1768 31214 1820 31220
rect 1780 30734 1808 31214
rect 1768 30728 1820 30734
rect 1768 30670 1820 30676
rect 1398 30288 1454 30297
rect 1398 30223 1454 30232
rect 1032 30184 1084 30190
rect 1032 30126 1084 30132
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1596 26217 1624 27950
rect 1780 27470 1808 30670
rect 2516 30394 2544 34326
rect 2594 34200 2650 34326
rect 4158 34200 4214 35000
rect 5722 34200 5778 35000
rect 7286 34200 7342 35000
rect 8850 34200 8906 35000
rect 10414 34200 10470 35000
rect 11978 34200 12034 35000
rect 13542 34200 13598 35000
rect 15106 34200 15162 35000
rect 16670 34354 16726 35000
rect 18234 34354 18290 35000
rect 19798 34354 19854 35000
rect 16670 34326 17080 34354
rect 16670 34200 16726 34326
rect 2872 32428 2924 32434
rect 2872 32370 2924 32376
rect 2884 32026 2912 32370
rect 2872 32020 2924 32026
rect 2872 31962 2924 31968
rect 4172 31890 4200 34200
rect 5736 32502 5764 34200
rect 5724 32496 5776 32502
rect 5724 32438 5776 32444
rect 7012 32496 7064 32502
rect 7012 32438 7064 32444
rect 6736 32360 6788 32366
rect 6736 32302 6788 32308
rect 4344 32224 4396 32230
rect 4344 32166 4396 32172
rect 6276 32224 6328 32230
rect 6276 32166 6328 32172
rect 6552 32224 6604 32230
rect 6552 32166 6604 32172
rect 4160 31884 4212 31890
rect 4160 31826 4212 31832
rect 4356 31822 4384 32166
rect 5044 32124 5352 32133
rect 5044 32122 5050 32124
rect 5106 32122 5130 32124
rect 5186 32122 5210 32124
rect 5266 32122 5290 32124
rect 5346 32122 5352 32124
rect 5106 32070 5108 32122
rect 5288 32070 5290 32122
rect 5044 32068 5050 32070
rect 5106 32068 5130 32070
rect 5186 32068 5210 32070
rect 5266 32068 5290 32070
rect 5346 32068 5352 32070
rect 5044 32059 5352 32068
rect 2596 31816 2648 31822
rect 2596 31758 2648 31764
rect 4344 31816 4396 31822
rect 4344 31758 4396 31764
rect 6184 31816 6236 31822
rect 6184 31758 6236 31764
rect 2504 30388 2556 30394
rect 2504 30330 2556 30336
rect 2608 30326 2636 31758
rect 3792 31680 3844 31686
rect 3792 31622 3844 31628
rect 4066 31648 4122 31657
rect 3804 31414 3832 31622
rect 4066 31583 4122 31592
rect 4080 31498 4108 31583
rect 4080 31470 4384 31498
rect 3792 31408 3844 31414
rect 3792 31350 3844 31356
rect 4160 30660 4212 30666
rect 4160 30602 4212 30608
rect 2596 30320 2648 30326
rect 2596 30262 2648 30268
rect 2964 30252 3016 30258
rect 3016 30212 3096 30240
rect 2964 30194 3016 30200
rect 2872 29504 2924 29510
rect 2872 29446 2924 29452
rect 2884 29170 2912 29446
rect 2872 29164 2924 29170
rect 2872 29106 2924 29112
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2596 28416 2648 28422
rect 2596 28358 2648 28364
rect 2608 28082 2636 28358
rect 2596 28076 2648 28082
rect 2596 28018 2648 28024
rect 2792 27577 2820 29038
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 2976 27674 3004 28494
rect 2964 27668 3016 27674
rect 2964 27610 3016 27616
rect 2778 27568 2834 27577
rect 2778 27503 2834 27512
rect 1768 27464 1820 27470
rect 1768 27406 1820 27412
rect 1780 26994 1808 27406
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 1582 26208 1638 26217
rect 1582 26143 1638 26152
rect 1780 25906 1808 26930
rect 2596 26784 2648 26790
rect 2596 26726 2648 26732
rect 2608 26382 2636 26726
rect 2792 26602 2820 26930
rect 2792 26574 2912 26602
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2596 26376 2648 26382
rect 2596 26318 2648 26324
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 940 24744 992 24750
rect 940 24686 992 24692
rect 952 23497 980 24686
rect 1584 23656 1636 23662
rect 1584 23598 1636 23604
rect 938 23488 994 23497
rect 938 23423 994 23432
rect 1596 22409 1624 23598
rect 1780 22642 1808 25842
rect 2792 24857 2820 26386
rect 2884 26042 2912 26574
rect 3068 26234 3096 30212
rect 4172 29850 4200 30602
rect 4160 29844 4212 29850
rect 4160 29786 4212 29792
rect 3424 29708 3476 29714
rect 3424 29650 3476 29656
rect 3332 29096 3384 29102
rect 3332 29038 3384 29044
rect 3344 28937 3372 29038
rect 3330 28928 3386 28937
rect 3330 28863 3386 28872
rect 2976 26206 3096 26234
rect 2872 26036 2924 26042
rect 2872 25978 2924 25984
rect 2778 24848 2834 24857
rect 2596 24812 2648 24818
rect 2778 24783 2834 24792
rect 2596 24754 2648 24760
rect 2608 24410 2636 24754
rect 2976 24410 3004 26206
rect 3436 25498 3464 29650
rect 4252 29640 4304 29646
rect 4252 29582 4304 29588
rect 3516 29504 3568 29510
rect 3516 29446 3568 29452
rect 3528 26234 3556 29446
rect 3608 29164 3660 29170
rect 3608 29106 3660 29112
rect 3620 28150 3648 29106
rect 3884 28552 3936 28558
rect 3884 28494 3936 28500
rect 3792 28484 3844 28490
rect 3792 28426 3844 28432
rect 3608 28144 3660 28150
rect 3608 28086 3660 28092
rect 3608 27396 3660 27402
rect 3608 27338 3660 27344
rect 3620 27130 3648 27338
rect 3608 27124 3660 27130
rect 3608 27066 3660 27072
rect 3804 26586 3832 28426
rect 3896 27674 3924 28494
rect 4160 28076 4212 28082
rect 4160 28018 4212 28024
rect 4172 27674 4200 28018
rect 3884 27668 3936 27674
rect 3884 27610 3936 27616
rect 4160 27668 4212 27674
rect 4160 27610 4212 27616
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4172 26586 4200 26930
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 4160 26580 4212 26586
rect 4160 26522 4212 26528
rect 4264 26518 4292 29582
rect 4356 29102 4384 31470
rect 6196 31414 6224 31758
rect 6000 31408 6052 31414
rect 6000 31350 6052 31356
rect 6184 31408 6236 31414
rect 6184 31350 6236 31356
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5724 31136 5776 31142
rect 5724 31078 5776 31084
rect 5044 31036 5352 31045
rect 5044 31034 5050 31036
rect 5106 31034 5130 31036
rect 5186 31034 5210 31036
rect 5266 31034 5290 31036
rect 5346 31034 5352 31036
rect 5106 30982 5108 31034
rect 5288 30982 5290 31034
rect 5044 30980 5050 30982
rect 5106 30980 5130 30982
rect 5186 30980 5210 30982
rect 5266 30980 5290 30982
rect 5346 30980 5352 30982
rect 5044 30971 5352 30980
rect 5460 30802 5488 31078
rect 5448 30796 5500 30802
rect 5448 30738 5500 30744
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5540 30660 5592 30666
rect 5540 30602 5592 30608
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4528 30048 4580 30054
rect 4528 29990 4580 29996
rect 4540 29714 4568 29990
rect 4632 29714 4660 30534
rect 5552 30258 5580 30602
rect 5540 30252 5592 30258
rect 5540 30194 5592 30200
rect 5044 29948 5352 29957
rect 5044 29946 5050 29948
rect 5106 29946 5130 29948
rect 5186 29946 5210 29948
rect 5266 29946 5290 29948
rect 5346 29946 5352 29948
rect 5106 29894 5108 29946
rect 5288 29894 5290 29946
rect 5044 29892 5050 29894
rect 5106 29892 5130 29894
rect 5186 29892 5210 29894
rect 5266 29892 5290 29894
rect 5346 29892 5352 29894
rect 5044 29883 5352 29892
rect 4528 29708 4580 29714
rect 4528 29650 4580 29656
rect 4620 29708 4672 29714
rect 4620 29650 4672 29656
rect 4896 29640 4948 29646
rect 4896 29582 4948 29588
rect 4436 29164 4488 29170
rect 4436 29106 4488 29112
rect 4344 29096 4396 29102
rect 4344 29038 4396 29044
rect 4448 28626 4476 29106
rect 4436 28620 4488 28626
rect 4436 28562 4488 28568
rect 4344 28416 4396 28422
rect 4344 28358 4396 28364
rect 4436 28416 4488 28422
rect 4436 28358 4488 28364
rect 4356 26994 4384 28358
rect 4448 27538 4476 28358
rect 4908 28218 4936 29582
rect 5044 28860 5352 28869
rect 5044 28858 5050 28860
rect 5106 28858 5130 28860
rect 5186 28858 5210 28860
rect 5266 28858 5290 28860
rect 5346 28858 5352 28860
rect 5106 28806 5108 28858
rect 5288 28806 5290 28858
rect 5044 28804 5050 28806
rect 5106 28804 5130 28806
rect 5186 28804 5210 28806
rect 5266 28804 5290 28806
rect 5346 28804 5352 28806
rect 5044 28795 5352 28804
rect 4896 28212 4948 28218
rect 4896 28154 4948 28160
rect 4804 28008 4856 28014
rect 4804 27950 4856 27956
rect 4816 27674 4844 27950
rect 4896 27872 4948 27878
rect 4896 27814 4948 27820
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4908 27538 4936 27814
rect 5044 27772 5352 27781
rect 5044 27770 5050 27772
rect 5106 27770 5130 27772
rect 5186 27770 5210 27772
rect 5266 27770 5290 27772
rect 5346 27770 5352 27772
rect 5106 27718 5108 27770
rect 5288 27718 5290 27770
rect 5044 27716 5050 27718
rect 5106 27716 5130 27718
rect 5186 27716 5210 27718
rect 5266 27716 5290 27718
rect 5346 27716 5352 27718
rect 5044 27707 5352 27716
rect 4436 27532 4488 27538
rect 4436 27474 4488 27480
rect 4896 27532 4948 27538
rect 4896 27474 4948 27480
rect 4448 27418 4476 27474
rect 4448 27390 4660 27418
rect 4344 26988 4396 26994
rect 4344 26930 4396 26936
rect 4436 26784 4488 26790
rect 4436 26726 4488 26732
rect 4252 26512 4304 26518
rect 4252 26454 4304 26460
rect 4448 26450 4476 26726
rect 4436 26444 4488 26450
rect 4436 26386 4488 26392
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 4160 26376 4212 26382
rect 4160 26318 4212 26324
rect 3792 26240 3844 26246
rect 3528 26206 3740 26234
rect 3424 25492 3476 25498
rect 3424 25434 3476 25440
rect 3148 25288 3200 25294
rect 3148 25230 3200 25236
rect 2596 24404 2648 24410
rect 2596 24346 2648 24352
rect 2964 24404 3016 24410
rect 2964 24346 3016 24352
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 2596 23724 2648 23730
rect 2596 23666 2648 23672
rect 2608 23186 2636 23666
rect 2976 23322 3004 24142
rect 3160 23526 3188 25230
rect 3332 24744 3384 24750
rect 3332 24686 3384 24692
rect 3344 24410 3372 24686
rect 3516 24608 3568 24614
rect 3516 24550 3568 24556
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2964 23316 3016 23322
rect 2964 23258 3016 23264
rect 3528 23186 3556 24550
rect 3620 23866 3648 24550
rect 3712 24274 3740 26206
rect 3792 26182 3844 26188
rect 3804 25838 3832 26182
rect 3988 26042 4016 26318
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 3792 25832 3844 25838
rect 3792 25774 3844 25780
rect 3804 24682 3832 25774
rect 4172 25498 4200 26318
rect 4448 25770 4476 26386
rect 4436 25764 4488 25770
rect 4436 25706 4488 25712
rect 4160 25492 4212 25498
rect 4160 25434 4212 25440
rect 4436 25288 4488 25294
rect 4436 25230 4488 25236
rect 4068 25220 4120 25226
rect 4068 25162 4120 25168
rect 4080 24886 4108 25162
rect 4068 24880 4120 24886
rect 4068 24822 4120 24828
rect 3792 24676 3844 24682
rect 3792 24618 3844 24624
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 4344 24200 4396 24206
rect 4344 24142 4396 24148
rect 4356 23866 4384 24142
rect 3608 23860 3660 23866
rect 3608 23802 3660 23808
rect 4344 23860 4396 23866
rect 4344 23802 4396 23808
rect 4448 23322 4476 25230
rect 4436 23316 4488 23322
rect 4436 23258 4488 23264
rect 4632 23254 4660 27390
rect 4908 26858 4936 27474
rect 5644 26994 5672 30670
rect 5736 30666 5764 31078
rect 5724 30660 5776 30666
rect 5724 30602 5776 30608
rect 5908 29504 5960 29510
rect 5908 29446 5960 29452
rect 5920 28626 5948 29446
rect 6012 28626 6040 31350
rect 6196 30326 6224 31350
rect 6288 31210 6316 32166
rect 6564 31890 6592 32166
rect 6748 32026 6776 32302
rect 6736 32020 6788 32026
rect 6736 31962 6788 31968
rect 6552 31884 6604 31890
rect 6552 31826 6604 31832
rect 6828 31340 6880 31346
rect 6828 31282 6880 31288
rect 6276 31204 6328 31210
rect 6276 31146 6328 31152
rect 6184 30320 6236 30326
rect 6184 30262 6236 30268
rect 6184 29776 6236 29782
rect 6184 29718 6236 29724
rect 5908 28620 5960 28626
rect 5908 28562 5960 28568
rect 6000 28620 6052 28626
rect 6000 28562 6052 28568
rect 6196 28422 6224 29718
rect 6288 29170 6316 31146
rect 6840 30394 6868 31282
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6828 30388 6880 30394
rect 6828 30330 6880 30336
rect 6368 30320 6420 30326
rect 6368 30262 6420 30268
rect 6380 29714 6408 30262
rect 6932 30258 6960 30534
rect 6920 30252 6972 30258
rect 6920 30194 6972 30200
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6656 29714 6684 29990
rect 7024 29850 7052 32438
rect 7300 31890 7328 34200
rect 8668 32428 8720 32434
rect 8668 32370 8720 32376
rect 8392 32360 8444 32366
rect 8392 32302 8444 32308
rect 8300 32224 8352 32230
rect 8300 32166 8352 32172
rect 7288 31884 7340 31890
rect 7288 31826 7340 31832
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 7472 31816 7524 31822
rect 7472 31758 7524 31764
rect 7116 29850 7144 31758
rect 7484 30802 7512 31758
rect 8312 31210 8340 32166
rect 8300 31204 8352 31210
rect 8300 31146 8352 31152
rect 7840 31136 7892 31142
rect 7840 31078 7892 31084
rect 7472 30796 7524 30802
rect 7472 30738 7524 30744
rect 7012 29844 7064 29850
rect 7012 29786 7064 29792
rect 7104 29844 7156 29850
rect 7104 29786 7156 29792
rect 7852 29714 7880 31078
rect 8024 30728 8076 30734
rect 8024 30670 8076 30676
rect 6368 29708 6420 29714
rect 6368 29650 6420 29656
rect 6644 29708 6696 29714
rect 6644 29650 6696 29656
rect 7840 29708 7892 29714
rect 7840 29650 7892 29656
rect 6276 29164 6328 29170
rect 6276 29106 6328 29112
rect 5724 28416 5776 28422
rect 5724 28358 5776 28364
rect 6184 28416 6236 28422
rect 6184 28358 6236 28364
rect 5736 28082 5764 28358
rect 5724 28076 5776 28082
rect 5724 28018 5776 28024
rect 5816 27464 5868 27470
rect 5816 27406 5868 27412
rect 5828 27130 5856 27406
rect 5816 27124 5868 27130
rect 5816 27066 5868 27072
rect 6380 27062 6408 29650
rect 8036 29306 8064 30670
rect 8312 30394 8340 31146
rect 8404 30734 8432 32302
rect 8392 30728 8444 30734
rect 8392 30670 8444 30676
rect 8300 30388 8352 30394
rect 8300 30330 8352 30336
rect 8680 30326 8708 32370
rect 8864 30802 8892 34200
rect 9138 32668 9446 32677
rect 9138 32666 9144 32668
rect 9200 32666 9224 32668
rect 9280 32666 9304 32668
rect 9360 32666 9384 32668
rect 9440 32666 9446 32668
rect 9200 32614 9202 32666
rect 9382 32614 9384 32666
rect 9138 32612 9144 32614
rect 9200 32612 9224 32614
rect 9280 32612 9304 32614
rect 9360 32612 9384 32614
rect 9440 32612 9446 32614
rect 9138 32603 9446 32612
rect 10428 32502 10456 34200
rect 10416 32496 10468 32502
rect 10416 32438 10468 32444
rect 11152 32428 11204 32434
rect 11152 32370 11204 32376
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9404 32292 9456 32298
rect 9404 32234 9456 32240
rect 9416 32026 9444 32234
rect 9404 32020 9456 32026
rect 9404 31962 9456 31968
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 8944 31680 8996 31686
rect 8944 31622 8996 31628
rect 8956 31278 8984 31622
rect 9138 31580 9446 31589
rect 9138 31578 9144 31580
rect 9200 31578 9224 31580
rect 9280 31578 9304 31580
rect 9360 31578 9384 31580
rect 9440 31578 9446 31580
rect 9200 31526 9202 31578
rect 9382 31526 9384 31578
rect 9138 31524 9144 31526
rect 9200 31524 9224 31526
rect 9280 31524 9304 31526
rect 9360 31524 9384 31526
rect 9440 31524 9446 31526
rect 9138 31515 9446 31524
rect 8944 31272 8996 31278
rect 8944 31214 8996 31220
rect 8852 30796 8904 30802
rect 8852 30738 8904 30744
rect 8956 30598 8984 31214
rect 8944 30592 8996 30598
rect 8944 30534 8996 30540
rect 8668 30320 8720 30326
rect 8668 30262 8720 30268
rect 8956 29714 8984 30534
rect 9138 30492 9446 30501
rect 9138 30490 9144 30492
rect 9200 30490 9224 30492
rect 9280 30490 9304 30492
rect 9360 30490 9384 30492
rect 9440 30490 9446 30492
rect 9200 30438 9202 30490
rect 9382 30438 9384 30490
rect 9138 30436 9144 30438
rect 9200 30436 9224 30438
rect 9280 30436 9304 30438
rect 9360 30436 9384 30438
rect 9440 30436 9446 30438
rect 9138 30427 9446 30436
rect 9692 30122 9720 31826
rect 9876 30326 9904 32302
rect 11164 32026 11192 32370
rect 11152 32020 11204 32026
rect 11152 31962 11204 31968
rect 11060 31952 11112 31958
rect 11060 31894 11112 31900
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 10140 31340 10192 31346
rect 10140 31282 10192 31288
rect 9864 30320 9916 30326
rect 9864 30262 9916 30268
rect 9680 30116 9732 30122
rect 9680 30058 9732 30064
rect 10152 29850 10180 31282
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 10428 30258 10456 31078
rect 10416 30252 10468 30258
rect 10416 30194 10468 30200
rect 10140 29844 10192 29850
rect 10140 29786 10192 29792
rect 10704 29782 10732 31078
rect 10876 30592 10928 30598
rect 10876 30534 10928 30540
rect 10888 30258 10916 30534
rect 10876 30252 10928 30258
rect 10876 30194 10928 30200
rect 10980 29850 11008 31758
rect 11072 30734 11100 31894
rect 11992 31754 12020 34200
rect 13556 32434 13584 34200
rect 15120 32586 15148 34200
rect 15120 32558 15240 32586
rect 15212 32502 15240 32558
rect 15200 32496 15252 32502
rect 15200 32438 15252 32444
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 14280 32428 14332 32434
rect 14280 32370 14332 32376
rect 15292 32428 15344 32434
rect 15292 32370 15344 32376
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 11980 31748 12032 31754
rect 11980 31690 12032 31696
rect 11336 31272 11388 31278
rect 11336 31214 11388 31220
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 11348 30394 11376 31214
rect 12360 30938 12388 31758
rect 12544 31482 12572 32302
rect 12900 32292 12952 32298
rect 12900 32234 12952 32240
rect 12532 31476 12584 31482
rect 12532 31418 12584 31424
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 12348 30932 12400 30938
rect 12348 30874 12400 30880
rect 11336 30388 11388 30394
rect 11336 30330 11388 30336
rect 12452 30258 12480 31078
rect 12912 30734 12940 32234
rect 13636 32224 13688 32230
rect 13636 32166 13688 32172
rect 13232 32124 13540 32133
rect 13232 32122 13238 32124
rect 13294 32122 13318 32124
rect 13374 32122 13398 32124
rect 13454 32122 13478 32124
rect 13534 32122 13540 32124
rect 13294 32070 13296 32122
rect 13476 32070 13478 32122
rect 13232 32068 13238 32070
rect 13294 32068 13318 32070
rect 13374 32068 13398 32070
rect 13454 32068 13478 32070
rect 13534 32068 13540 32070
rect 13232 32059 13540 32068
rect 12992 31340 13044 31346
rect 12992 31282 13044 31288
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 13004 30394 13032 31282
rect 13084 31272 13136 31278
rect 13084 31214 13136 31220
rect 13096 30734 13124 31214
rect 13232 31036 13540 31045
rect 13232 31034 13238 31036
rect 13294 31034 13318 31036
rect 13374 31034 13398 31036
rect 13454 31034 13478 31036
rect 13534 31034 13540 31036
rect 13294 30982 13296 31034
rect 13476 30982 13478 31034
rect 13232 30980 13238 30982
rect 13294 30980 13318 30982
rect 13374 30980 13398 30982
rect 13454 30980 13478 30982
rect 13534 30980 13540 30982
rect 13232 30971 13540 30980
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 12992 30388 13044 30394
rect 12992 30330 13044 30336
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 11152 30184 11204 30190
rect 11152 30126 11204 30132
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 10692 29776 10744 29782
rect 10692 29718 10744 29724
rect 11164 29714 11192 30126
rect 8944 29708 8996 29714
rect 8944 29650 8996 29656
rect 11152 29708 11204 29714
rect 11152 29650 11204 29656
rect 8024 29300 8076 29306
rect 8024 29242 8076 29248
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 5724 27056 5776 27062
rect 5724 26998 5776 27004
rect 6368 27056 6420 27062
rect 6368 26998 6420 27004
rect 5632 26988 5684 26994
rect 5632 26930 5684 26936
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 5044 26684 5352 26693
rect 5044 26682 5050 26684
rect 5106 26682 5130 26684
rect 5186 26682 5210 26684
rect 5266 26682 5290 26684
rect 5346 26682 5352 26684
rect 5106 26630 5108 26682
rect 5288 26630 5290 26682
rect 5044 26628 5050 26630
rect 5106 26628 5130 26630
rect 5186 26628 5210 26630
rect 5266 26628 5290 26630
rect 5346 26628 5352 26630
rect 5044 26619 5352 26628
rect 5448 26512 5500 26518
rect 5448 26454 5500 26460
rect 4896 25832 4948 25838
rect 4896 25774 4948 25780
rect 4908 24886 4936 25774
rect 5044 25596 5352 25605
rect 5044 25594 5050 25596
rect 5106 25594 5130 25596
rect 5186 25594 5210 25596
rect 5266 25594 5290 25596
rect 5346 25594 5352 25596
rect 5106 25542 5108 25594
rect 5288 25542 5290 25594
rect 5044 25540 5050 25542
rect 5106 25540 5130 25542
rect 5186 25540 5210 25542
rect 5266 25540 5290 25542
rect 5346 25540 5352 25542
rect 5044 25531 5352 25540
rect 5460 25294 5488 26454
rect 5736 26450 5764 26998
rect 7116 26994 7144 28358
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 5724 26444 5776 26450
rect 5724 26386 5776 26392
rect 5736 26234 5764 26386
rect 7116 26234 7144 26930
rect 5736 26206 5948 26234
rect 5920 25838 5948 26206
rect 7024 26206 7144 26234
rect 5908 25832 5960 25838
rect 5908 25774 5960 25780
rect 7024 25362 7052 26206
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 5448 25288 5500 25294
rect 5448 25230 5500 25236
rect 4896 24880 4948 24886
rect 4896 24822 4948 24828
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4620 23248 4672 23254
rect 4620 23190 4672 23196
rect 2596 23180 2648 23186
rect 2596 23122 2648 23128
rect 3516 23180 3568 23186
rect 3516 23122 3568 23128
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1582 22400 1638 22409
rect 1582 22335 1638 22344
rect 1780 22098 1808 22578
rect 3252 22234 3280 23054
rect 3528 22778 3556 23122
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 1768 22092 1820 22098
rect 1768 22034 1820 22040
rect 940 21480 992 21486
rect 940 21422 992 21428
rect 952 20777 980 21422
rect 1780 21010 1808 22034
rect 2596 21548 2648 21554
rect 2596 21490 2648 21496
rect 1768 21004 1820 21010
rect 1768 20946 1820 20952
rect 938 20768 994 20777
rect 938 20703 994 20712
rect 1780 19922 1808 20946
rect 2608 20534 2636 21490
rect 3700 21480 3752 21486
rect 3700 21422 3752 21428
rect 3516 21344 3568 21350
rect 3516 21286 3568 21292
rect 3608 21344 3660 21350
rect 3608 21286 3660 21292
rect 2596 20528 2648 20534
rect 2596 20470 2648 20476
rect 3528 20482 3556 21286
rect 3620 20942 3648 21286
rect 3712 21146 3740 21422
rect 3804 21146 3832 23054
rect 4528 22976 4580 22982
rect 4528 22918 4580 22924
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 4356 22098 4384 22374
rect 4344 22092 4396 22098
rect 4344 22034 4396 22040
rect 4356 21486 4384 22034
rect 4540 22030 4568 22918
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 4344 21480 4396 21486
rect 4344 21422 4396 21428
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 3528 20454 3648 20482
rect 3620 20398 3648 20454
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 938 19408 994 19417
rect 938 19343 940 19352
rect 992 19343 994 19352
rect 940 19314 992 19320
rect 1308 18148 1360 18154
rect 1308 18090 1360 18096
rect 1320 18057 1348 18090
rect 1306 18048 1362 18057
rect 1306 17983 1362 17992
rect 1780 17746 1808 19858
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 1952 18896 2004 18902
rect 1952 18838 2004 18844
rect 1964 18426 1992 18838
rect 2608 18834 2636 19314
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2884 18970 2912 19246
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 3160 18834 3188 19654
rect 3252 19514 3280 19722
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3620 19242 3648 20334
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3608 19236 3660 19242
rect 3608 19178 3660 19184
rect 3712 18970 3740 19246
rect 3700 18964 3752 18970
rect 3700 18906 3752 18912
rect 2596 18828 2648 18834
rect 2596 18770 2648 18776
rect 3148 18828 3200 18834
rect 3148 18770 3200 18776
rect 3804 18766 3832 19654
rect 4448 19378 4476 19790
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 4264 18834 4292 19110
rect 4252 18828 4304 18834
rect 4252 18770 4304 18776
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3804 18426 3832 18566
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 1768 17740 1820 17746
rect 1768 17682 1820 17688
rect 1780 17202 1808 17682
rect 3516 17536 3568 17542
rect 3516 17478 3568 17484
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1582 16688 1638 16697
rect 1780 16658 1808 17138
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3344 16794 3372 17070
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 1582 16623 1638 16632
rect 1768 16652 1820 16658
rect 1596 15570 1624 16623
rect 1768 16594 1820 16600
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 1596 14482 1624 15263
rect 1780 14958 1808 15982
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1306 13968 1362 13977
rect 1306 13903 1362 13912
rect 1320 13870 1348 13903
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1780 12782 1808 14894
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2608 14074 2636 14350
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13394 2820 13874
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2884 13326 2912 14214
rect 2976 14074 3004 15302
rect 3436 14482 3464 15846
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 3436 13802 3464 14418
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2872 13184 2924 13190
rect 2872 13126 2924 13132
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1582 12472 1638 12481
rect 1582 12407 1638 12416
rect 1596 11830 1624 12407
rect 1584 11824 1636 11830
rect 1584 11766 1636 11772
rect 1308 11688 1360 11694
rect 1308 11630 1360 11636
rect 1320 11257 1348 11630
rect 1306 11248 1362 11257
rect 1306 11183 1362 11192
rect 1780 11150 1808 12718
rect 2884 12238 2912 13126
rect 3148 12640 3200 12646
rect 3148 12582 3200 12588
rect 3160 12306 3188 12582
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11762 2636 12038
rect 2596 11756 2648 11762
rect 2596 11698 2648 11704
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10062 1808 11086
rect 2884 10742 2912 11698
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 1768 10056 1820 10062
rect 1768 9998 1820 10004
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1596 9654 1624 9687
rect 1584 9648 1636 9654
rect 1584 9590 1636 9596
rect 1780 8430 1808 9998
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2608 9178 2636 9522
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 9178 2912 9318
rect 2596 9172 2648 9178
rect 2596 9114 2648 9120
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 1768 8424 1820 8430
rect 1582 8392 1638 8401
rect 1768 8366 1820 8372
rect 1582 8327 1638 8336
rect 1596 7954 1624 8327
rect 1584 7948 1636 7954
rect 1584 7890 1636 7896
rect 1780 7546 1808 8366
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1582 7032 1638 7041
rect 1582 6967 1638 6976
rect 1308 6112 1360 6118
rect 1308 6054 1360 6060
rect 1320 5817 1348 6054
rect 1306 5808 1362 5817
rect 1596 5778 1624 6967
rect 1780 6866 1808 7482
rect 2608 7478 2636 7822
rect 2596 7472 2648 7478
rect 2596 7414 2648 7420
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6322 1808 6802
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1306 5743 1362 5752
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2608 5302 2636 5646
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2792 5234 2820 6598
rect 2884 5778 2912 7142
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 1582 4176 1638 4185
rect 2976 4146 3004 10406
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9586 3188 9862
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 7410 3188 8774
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 7954 3280 8230
rect 3240 7948 3292 7954
rect 3240 7890 3292 7896
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5234 3188 6054
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 3252 4690 3280 6258
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 1582 4111 1638 4120
rect 2964 4140 3016 4146
rect 1596 3602 1624 4111
rect 2964 4082 3016 4088
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 2608 3534 2636 3878
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 3436 3058 3464 13126
rect 3528 12850 3556 17478
rect 3896 16590 3924 18566
rect 4172 17882 4200 18702
rect 4264 18170 4292 18770
rect 4264 18142 4384 18170
rect 4448 18154 4476 19314
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 4264 17678 4292 18022
rect 4356 17814 4384 18142
rect 4436 18148 4488 18154
rect 4436 18090 4488 18096
rect 4344 17808 4396 17814
rect 4344 17750 4396 17756
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3988 16114 4016 16934
rect 4172 16794 4200 17138
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4264 16182 4292 17478
rect 4540 17338 4568 20878
rect 4632 17678 4660 21830
rect 4724 18902 4752 24142
rect 4908 23050 4936 24822
rect 5044 24508 5352 24517
rect 5044 24506 5050 24508
rect 5106 24506 5130 24508
rect 5186 24506 5210 24508
rect 5266 24506 5290 24508
rect 5346 24506 5352 24508
rect 5106 24454 5108 24506
rect 5288 24454 5290 24506
rect 5044 24452 5050 24454
rect 5106 24452 5130 24454
rect 5186 24452 5210 24454
rect 5266 24452 5290 24454
rect 5346 24452 5352 24454
rect 5044 24443 5352 24452
rect 5044 23420 5352 23429
rect 5044 23418 5050 23420
rect 5106 23418 5130 23420
rect 5186 23418 5210 23420
rect 5266 23418 5290 23420
rect 5346 23418 5352 23420
rect 5106 23366 5108 23418
rect 5288 23366 5290 23418
rect 5044 23364 5050 23366
rect 5106 23364 5130 23366
rect 5186 23364 5210 23366
rect 5266 23364 5290 23366
rect 5346 23364 5352 23366
rect 5044 23355 5352 23364
rect 4896 23044 4948 23050
rect 4896 22986 4948 22992
rect 4908 22574 4936 22986
rect 4896 22568 4948 22574
rect 4816 22516 4896 22522
rect 4816 22510 4948 22516
rect 4816 22494 4936 22510
rect 4816 21486 4844 22494
rect 5044 22332 5352 22341
rect 5044 22330 5050 22332
rect 5106 22330 5130 22332
rect 5186 22330 5210 22332
rect 5266 22330 5290 22332
rect 5346 22330 5352 22332
rect 5106 22278 5108 22330
rect 5288 22278 5290 22330
rect 5044 22276 5050 22278
rect 5106 22276 5130 22278
rect 5186 22276 5210 22278
rect 5266 22276 5290 22278
rect 5346 22276 5352 22278
rect 5044 22267 5352 22276
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4816 19310 4844 21422
rect 5044 21244 5352 21253
rect 5044 21242 5050 21244
rect 5106 21242 5130 21244
rect 5186 21242 5210 21244
rect 5266 21242 5290 21244
rect 5346 21242 5352 21244
rect 5106 21190 5108 21242
rect 5288 21190 5290 21242
rect 5044 21188 5050 21190
rect 5106 21188 5130 21190
rect 5186 21188 5210 21190
rect 5266 21188 5290 21190
rect 5346 21188 5352 21190
rect 5044 21179 5352 21188
rect 5044 20156 5352 20165
rect 5044 20154 5050 20156
rect 5106 20154 5130 20156
rect 5186 20154 5210 20156
rect 5266 20154 5290 20156
rect 5346 20154 5352 20156
rect 5106 20102 5108 20154
rect 5288 20102 5290 20154
rect 5044 20100 5050 20102
rect 5106 20100 5130 20102
rect 5186 20100 5210 20102
rect 5266 20100 5290 20102
rect 5346 20100 5352 20102
rect 5044 20091 5352 20100
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 4816 18834 4844 19246
rect 5044 19068 5352 19077
rect 5044 19066 5050 19068
rect 5106 19066 5130 19068
rect 5186 19066 5210 19068
rect 5266 19066 5290 19068
rect 5346 19066 5352 19068
rect 5106 19014 5108 19066
rect 5288 19014 5290 19066
rect 5044 19012 5050 19014
rect 5106 19012 5130 19014
rect 5186 19012 5210 19014
rect 5266 19012 5290 19014
rect 5346 19012 5352 19014
rect 5044 19003 5352 19012
rect 8956 18970 8984 29650
rect 9138 29404 9446 29413
rect 9138 29402 9144 29404
rect 9200 29402 9224 29404
rect 9280 29402 9304 29404
rect 9360 29402 9384 29404
rect 9440 29402 9446 29404
rect 9200 29350 9202 29402
rect 9382 29350 9384 29402
rect 9138 29348 9144 29350
rect 9200 29348 9224 29350
rect 9280 29348 9304 29350
rect 9360 29348 9384 29350
rect 9440 29348 9446 29350
rect 9138 29339 9446 29348
rect 10416 28552 10468 28558
rect 10416 28494 10468 28500
rect 9138 28316 9446 28325
rect 9138 28314 9144 28316
rect 9200 28314 9224 28316
rect 9280 28314 9304 28316
rect 9360 28314 9384 28316
rect 9440 28314 9446 28316
rect 9200 28262 9202 28314
rect 9382 28262 9384 28314
rect 9138 28260 9144 28262
rect 9200 28260 9224 28262
rect 9280 28260 9304 28262
rect 9360 28260 9384 28262
rect 9440 28260 9446 28262
rect 9138 28251 9446 28260
rect 9138 27228 9446 27237
rect 9138 27226 9144 27228
rect 9200 27226 9224 27228
rect 9280 27226 9304 27228
rect 9360 27226 9384 27228
rect 9440 27226 9446 27228
rect 9200 27174 9202 27226
rect 9382 27174 9384 27226
rect 9138 27172 9144 27174
rect 9200 27172 9224 27174
rect 9280 27172 9304 27174
rect 9360 27172 9384 27174
rect 9440 27172 9446 27174
rect 9138 27163 9446 27172
rect 10428 27130 10456 28494
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 12072 26920 12124 26926
rect 12072 26862 12124 26868
rect 9138 26140 9446 26149
rect 9138 26138 9144 26140
rect 9200 26138 9224 26140
rect 9280 26138 9304 26140
rect 9360 26138 9384 26140
rect 9440 26138 9446 26140
rect 9200 26086 9202 26138
rect 9382 26086 9384 26138
rect 9138 26084 9144 26086
rect 9200 26084 9224 26086
rect 9280 26084 9304 26086
rect 9360 26084 9384 26086
rect 9440 26084 9446 26086
rect 9138 26075 9446 26084
rect 9138 25052 9446 25061
rect 9138 25050 9144 25052
rect 9200 25050 9224 25052
rect 9280 25050 9304 25052
rect 9360 25050 9384 25052
rect 9440 25050 9446 25052
rect 9200 24998 9202 25050
rect 9382 24998 9384 25050
rect 9138 24996 9144 24998
rect 9200 24996 9224 24998
rect 9280 24996 9304 24998
rect 9360 24996 9384 24998
rect 9440 24996 9446 24998
rect 9138 24987 9446 24996
rect 12084 24614 12112 26862
rect 13096 24614 13124 30670
rect 13648 30054 13676 32166
rect 14292 30734 14320 32370
rect 14464 32360 14516 32366
rect 14464 32302 14516 32308
rect 14476 31482 14504 32302
rect 15304 32026 15332 32370
rect 16120 32224 16172 32230
rect 16120 32166 16172 32172
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 15292 32020 15344 32026
rect 15292 31962 15344 31968
rect 14556 31816 14608 31822
rect 14556 31758 14608 31764
rect 14464 31476 14516 31482
rect 14464 31418 14516 31424
rect 14464 31340 14516 31346
rect 14464 31282 14516 31288
rect 13728 30728 13780 30734
rect 13728 30670 13780 30676
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 13740 30394 13768 30670
rect 14476 30394 14504 31282
rect 14568 30870 14596 31758
rect 14556 30864 14608 30870
rect 14556 30806 14608 30812
rect 13728 30388 13780 30394
rect 13728 30330 13780 30336
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 13740 30122 13768 30330
rect 14568 30122 14596 30806
rect 16132 30802 16160 32166
rect 16868 32026 16896 32166
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16120 30796 16172 30802
rect 16120 30738 16172 30744
rect 16316 30394 16344 31282
rect 16672 31136 16724 31142
rect 16672 31078 16724 31084
rect 16684 30938 16712 31078
rect 16672 30932 16724 30938
rect 16672 30874 16724 30880
rect 17052 30802 17080 34326
rect 18234 34326 18552 34354
rect 18234 34200 18290 34326
rect 17326 32668 17634 32677
rect 17326 32666 17332 32668
rect 17388 32666 17412 32668
rect 17468 32666 17492 32668
rect 17548 32666 17572 32668
rect 17628 32666 17634 32668
rect 17388 32614 17390 32666
rect 17570 32614 17572 32666
rect 17326 32612 17332 32614
rect 17388 32612 17412 32614
rect 17468 32612 17492 32614
rect 17548 32612 17572 32614
rect 17628 32612 17634 32614
rect 17326 32603 17634 32612
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 17040 30796 17092 30802
rect 17040 30738 17092 30744
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 14556 30116 14608 30122
rect 14556 30058 14608 30064
rect 13636 30048 13688 30054
rect 13636 29990 13688 29996
rect 15752 30048 15804 30054
rect 15752 29990 15804 29996
rect 13232 29948 13540 29957
rect 13232 29946 13238 29948
rect 13294 29946 13318 29948
rect 13374 29946 13398 29948
rect 13454 29946 13478 29948
rect 13534 29946 13540 29948
rect 13294 29894 13296 29946
rect 13476 29894 13478 29946
rect 13232 29892 13238 29894
rect 13294 29892 13318 29894
rect 13374 29892 13398 29894
rect 13454 29892 13478 29894
rect 13534 29892 13540 29894
rect 13232 29883 13540 29892
rect 13232 28860 13540 28869
rect 13232 28858 13238 28860
rect 13294 28858 13318 28860
rect 13374 28858 13398 28860
rect 13454 28858 13478 28860
rect 13534 28858 13540 28860
rect 13294 28806 13296 28858
rect 13476 28806 13478 28858
rect 13232 28804 13238 28806
rect 13294 28804 13318 28806
rect 13374 28804 13398 28806
rect 13454 28804 13478 28806
rect 13534 28804 13540 28806
rect 13232 28795 13540 28804
rect 13232 27772 13540 27781
rect 13232 27770 13238 27772
rect 13294 27770 13318 27772
rect 13374 27770 13398 27772
rect 13454 27770 13478 27772
rect 13534 27770 13540 27772
rect 13294 27718 13296 27770
rect 13476 27718 13478 27770
rect 13232 27716 13238 27718
rect 13294 27716 13318 27718
rect 13374 27716 13398 27718
rect 13454 27716 13478 27718
rect 13534 27716 13540 27718
rect 13232 27707 13540 27716
rect 13232 26684 13540 26693
rect 13232 26682 13238 26684
rect 13294 26682 13318 26684
rect 13374 26682 13398 26684
rect 13454 26682 13478 26684
rect 13534 26682 13540 26684
rect 13294 26630 13296 26682
rect 13476 26630 13478 26682
rect 13232 26628 13238 26630
rect 13294 26628 13318 26630
rect 13374 26628 13398 26630
rect 13454 26628 13478 26630
rect 13534 26628 13540 26630
rect 13232 26619 13540 26628
rect 13232 25596 13540 25605
rect 13232 25594 13238 25596
rect 13294 25594 13318 25596
rect 13374 25594 13398 25596
rect 13454 25594 13478 25596
rect 13534 25594 13540 25596
rect 13294 25542 13296 25594
rect 13476 25542 13478 25594
rect 13232 25540 13238 25542
rect 13294 25540 13318 25542
rect 13374 25540 13398 25542
rect 13454 25540 13478 25542
rect 13534 25540 13540 25542
rect 13232 25531 13540 25540
rect 15764 24818 15792 29990
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16776 25838 16804 26182
rect 17144 26042 17172 32370
rect 18524 32366 18552 34326
rect 19798 34326 20208 34354
rect 19798 34200 19854 34326
rect 17684 32360 17736 32366
rect 17684 32302 17736 32308
rect 18512 32360 18564 32366
rect 18512 32302 18564 32308
rect 17224 31748 17276 31754
rect 17224 31690 17276 31696
rect 17236 30734 17264 31690
rect 17326 31580 17634 31589
rect 17326 31578 17332 31580
rect 17388 31578 17412 31580
rect 17468 31578 17492 31580
rect 17548 31578 17572 31580
rect 17628 31578 17634 31580
rect 17388 31526 17390 31578
rect 17570 31526 17572 31578
rect 17326 31524 17332 31526
rect 17388 31524 17412 31526
rect 17468 31524 17492 31526
rect 17548 31524 17572 31526
rect 17628 31524 17634 31526
rect 17326 31515 17634 31524
rect 17696 31142 17724 32302
rect 20180 32298 20208 34326
rect 21362 34200 21418 35000
rect 22926 34354 22982 35000
rect 24490 34354 24546 35000
rect 22926 34326 23336 34354
rect 22926 34200 22982 34326
rect 21376 32502 21404 34200
rect 21364 32496 21416 32502
rect 21364 32438 21416 32444
rect 21824 32428 21876 32434
rect 21824 32370 21876 32376
rect 20904 32360 20956 32366
rect 20904 32302 20956 32308
rect 20168 32292 20220 32298
rect 20168 32234 20220 32240
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 18524 31890 18552 32166
rect 18512 31884 18564 31890
rect 18512 31826 18564 31832
rect 18144 31680 18196 31686
rect 18144 31622 18196 31628
rect 18156 31346 18184 31622
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 18144 31340 18196 31346
rect 18144 31282 18196 31288
rect 17684 31136 17736 31142
rect 17684 31078 17736 31084
rect 17224 30728 17276 30734
rect 17224 30670 17276 30676
rect 17326 30492 17634 30501
rect 17326 30490 17332 30492
rect 17388 30490 17412 30492
rect 17468 30490 17492 30492
rect 17548 30490 17572 30492
rect 17628 30490 17634 30492
rect 17388 30438 17390 30490
rect 17570 30438 17572 30490
rect 17326 30436 17332 30438
rect 17388 30436 17412 30438
rect 17468 30436 17492 30438
rect 17548 30436 17572 30438
rect 17628 30436 17634 30438
rect 17326 30427 17634 30436
rect 17696 30122 17724 31078
rect 17972 30394 18000 31282
rect 17960 30388 18012 30394
rect 17960 30330 18012 30336
rect 18524 30122 18552 31826
rect 20260 31680 20312 31686
rect 20260 31622 20312 31628
rect 20272 31346 20300 31622
rect 20260 31340 20312 31346
rect 20260 31282 20312 31288
rect 18696 31272 18748 31278
rect 18696 31214 18748 31220
rect 18708 30938 18736 31214
rect 18880 31136 18932 31142
rect 18880 31078 18932 31084
rect 18892 30938 18920 31078
rect 20272 30938 20300 31282
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18880 30932 18932 30938
rect 18880 30874 18932 30880
rect 20260 30932 20312 30938
rect 20260 30874 20312 30880
rect 20916 30734 20944 32302
rect 21420 32124 21728 32133
rect 21420 32122 21426 32124
rect 21482 32122 21506 32124
rect 21562 32122 21586 32124
rect 21642 32122 21666 32124
rect 21722 32122 21728 32124
rect 21482 32070 21484 32122
rect 21664 32070 21666 32122
rect 21420 32068 21426 32070
rect 21482 32068 21506 32070
rect 21562 32068 21586 32070
rect 21642 32068 21666 32070
rect 21722 32068 21728 32070
rect 21420 32059 21728 32068
rect 21836 32026 21864 32370
rect 22008 32360 22060 32366
rect 22008 32302 22060 32308
rect 21824 32020 21876 32026
rect 21824 31962 21876 31968
rect 21272 31680 21324 31686
rect 21272 31622 21324 31628
rect 21284 31278 21312 31622
rect 21272 31272 21324 31278
rect 21272 31214 21324 31220
rect 21916 31272 21968 31278
rect 21916 31214 21968 31220
rect 20904 30728 20956 30734
rect 20904 30670 20956 30676
rect 21180 30660 21232 30666
rect 21180 30602 21232 30608
rect 21192 30394 21220 30602
rect 21180 30388 21232 30394
rect 21180 30330 21232 30336
rect 21284 30258 21312 31214
rect 21420 31036 21728 31045
rect 21420 31034 21426 31036
rect 21482 31034 21506 31036
rect 21562 31034 21586 31036
rect 21642 31034 21666 31036
rect 21722 31034 21728 31036
rect 21482 30982 21484 31034
rect 21664 30982 21666 31034
rect 21420 30980 21426 30982
rect 21482 30980 21506 30982
rect 21562 30980 21586 30982
rect 21642 30980 21666 30982
rect 21722 30980 21728 30982
rect 21420 30971 21728 30980
rect 21928 30938 21956 31214
rect 21916 30932 21968 30938
rect 21916 30874 21968 30880
rect 21272 30252 21324 30258
rect 21272 30194 21324 30200
rect 22020 30190 22048 32302
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22388 31260 22416 31758
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22388 31232 22508 31260
rect 22100 31136 22152 31142
rect 22100 31078 22152 31084
rect 22112 30938 22140 31078
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 22480 30394 22508 31232
rect 22468 30388 22520 30394
rect 22468 30330 22520 30336
rect 22008 30184 22060 30190
rect 22008 30126 22060 30132
rect 22940 30122 22968 31282
rect 23308 30666 23336 34326
rect 24490 34326 24808 34354
rect 24490 34200 24546 34326
rect 24780 32586 24808 34326
rect 26054 34200 26110 35000
rect 27618 34200 27674 35000
rect 29182 34200 29238 35000
rect 30746 34354 30802 35000
rect 32310 34354 32366 35000
rect 33874 34354 33930 35000
rect 30746 34326 30880 34354
rect 30746 34200 30802 34326
rect 25514 32668 25822 32677
rect 25514 32666 25520 32668
rect 25576 32666 25600 32668
rect 25656 32666 25680 32668
rect 25736 32666 25760 32668
rect 25816 32666 25822 32668
rect 25576 32614 25578 32666
rect 25758 32614 25760 32666
rect 25514 32612 25520 32614
rect 25576 32612 25600 32614
rect 25656 32612 25680 32614
rect 25736 32612 25760 32614
rect 25816 32612 25822 32614
rect 25514 32603 25822 32612
rect 24780 32558 24992 32586
rect 24400 32428 24452 32434
rect 24964 32416 24992 32558
rect 25044 32428 25096 32434
rect 24964 32388 25044 32416
rect 24400 32370 24452 32376
rect 25044 32370 25096 32376
rect 24412 32026 24440 32370
rect 26068 32366 26096 34200
rect 26976 32428 27028 32434
rect 26976 32370 27028 32376
rect 26056 32360 26108 32366
rect 26056 32302 26108 32308
rect 26424 32360 26476 32366
rect 26424 32302 26476 32308
rect 26148 32224 26200 32230
rect 26148 32166 26200 32172
rect 24400 32020 24452 32026
rect 24400 31962 24452 31968
rect 26160 31822 26188 32166
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 24676 31816 24728 31822
rect 24676 31758 24728 31764
rect 26148 31816 26200 31822
rect 26148 31758 26200 31764
rect 23400 31482 23428 31758
rect 23388 31476 23440 31482
rect 23388 31418 23440 31424
rect 23388 31340 23440 31346
rect 23388 31282 23440 31288
rect 23296 30660 23348 30666
rect 23296 30602 23348 30608
rect 23400 30394 23428 31282
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23676 30938 23704 31078
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23388 30388 23440 30394
rect 23388 30330 23440 30336
rect 24688 30326 24716 31758
rect 25412 31680 25464 31686
rect 25412 31622 25464 31628
rect 25424 31346 25452 31622
rect 25514 31580 25822 31589
rect 25514 31578 25520 31580
rect 25576 31578 25600 31580
rect 25656 31578 25680 31580
rect 25736 31578 25760 31580
rect 25816 31578 25822 31580
rect 25576 31526 25578 31578
rect 25758 31526 25760 31578
rect 25514 31524 25520 31526
rect 25576 31524 25600 31526
rect 25656 31524 25680 31526
rect 25736 31524 25760 31526
rect 25816 31524 25822 31526
rect 25514 31515 25822 31524
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 25412 31340 25464 31346
rect 25412 31282 25464 31288
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 24964 30938 24992 31282
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 26240 30864 26292 30870
rect 26240 30806 26292 30812
rect 25320 30660 25372 30666
rect 25320 30602 25372 30608
rect 24676 30320 24728 30326
rect 24676 30262 24728 30268
rect 23572 30184 23624 30190
rect 23572 30126 23624 30132
rect 17684 30116 17736 30122
rect 17684 30058 17736 30064
rect 18512 30116 18564 30122
rect 18512 30058 18564 30064
rect 22928 30116 22980 30122
rect 22928 30058 22980 30064
rect 21420 29948 21728 29957
rect 21420 29946 21426 29948
rect 21482 29946 21506 29948
rect 21562 29946 21586 29948
rect 21642 29946 21666 29948
rect 21722 29946 21728 29948
rect 21482 29894 21484 29946
rect 21664 29894 21666 29946
rect 21420 29892 21426 29894
rect 21482 29892 21506 29894
rect 21562 29892 21586 29894
rect 21642 29892 21666 29894
rect 21722 29892 21728 29894
rect 21420 29883 21728 29892
rect 23584 29646 23612 30126
rect 24952 30116 25004 30122
rect 24952 30058 25004 30064
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 23572 29640 23624 29646
rect 23572 29582 23624 29588
rect 17326 29404 17634 29413
rect 17326 29402 17332 29404
rect 17388 29402 17412 29404
rect 17468 29402 17492 29404
rect 17548 29402 17572 29404
rect 17628 29402 17634 29404
rect 17388 29350 17390 29402
rect 17570 29350 17572 29402
rect 17326 29348 17332 29350
rect 17388 29348 17412 29350
rect 17468 29348 17492 29350
rect 17548 29348 17572 29350
rect 17628 29348 17634 29350
rect 17326 29339 17634 29348
rect 21420 28860 21728 28869
rect 21420 28858 21426 28860
rect 21482 28858 21506 28860
rect 21562 28858 21586 28860
rect 21642 28858 21666 28860
rect 21722 28858 21728 28860
rect 21482 28806 21484 28858
rect 21664 28806 21666 28858
rect 21420 28804 21426 28806
rect 21482 28804 21506 28806
rect 21562 28804 21586 28806
rect 21642 28804 21666 28806
rect 21722 28804 21728 28806
rect 21420 28795 21728 28804
rect 17326 28316 17634 28325
rect 17326 28314 17332 28316
rect 17388 28314 17412 28316
rect 17468 28314 17492 28316
rect 17548 28314 17572 28316
rect 17628 28314 17634 28316
rect 17388 28262 17390 28314
rect 17570 28262 17572 28314
rect 17326 28260 17332 28262
rect 17388 28260 17412 28262
rect 17468 28260 17492 28262
rect 17548 28260 17572 28262
rect 17628 28260 17634 28262
rect 17326 28251 17634 28260
rect 21420 27772 21728 27781
rect 21420 27770 21426 27772
rect 21482 27770 21506 27772
rect 21562 27770 21586 27772
rect 21642 27770 21666 27772
rect 21722 27770 21728 27772
rect 21482 27718 21484 27770
rect 21664 27718 21666 27770
rect 21420 27716 21426 27718
rect 21482 27716 21506 27718
rect 21562 27716 21586 27718
rect 21642 27716 21666 27718
rect 21722 27716 21728 27718
rect 21420 27707 21728 27716
rect 24872 27606 24900 29650
rect 24964 28558 24992 30058
rect 25332 29646 25360 30602
rect 25412 30592 25464 30598
rect 25412 30534 25464 30540
rect 25424 30258 25452 30534
rect 25514 30492 25822 30501
rect 25514 30490 25520 30492
rect 25576 30490 25600 30492
rect 25656 30490 25680 30492
rect 25736 30490 25760 30492
rect 25816 30490 25822 30492
rect 25576 30438 25578 30490
rect 25758 30438 25760 30490
rect 25514 30436 25520 30438
rect 25576 30436 25600 30438
rect 25656 30436 25680 30438
rect 25736 30436 25760 30438
rect 25816 30436 25822 30438
rect 25514 30427 25822 30436
rect 25412 30252 25464 30258
rect 25412 30194 25464 30200
rect 26252 30190 26280 30806
rect 26344 30190 26372 31282
rect 26436 30938 26464 32302
rect 26884 32224 26936 32230
rect 26884 32166 26936 32172
rect 26516 31748 26568 31754
rect 26516 31690 26568 31696
rect 26424 30932 26476 30938
rect 26424 30874 26476 30880
rect 26528 30734 26556 31690
rect 26516 30728 26568 30734
rect 26516 30670 26568 30676
rect 26700 30592 26752 30598
rect 26700 30534 26752 30540
rect 26240 30184 26292 30190
rect 26240 30126 26292 30132
rect 26332 30184 26384 30190
rect 26332 30126 26384 30132
rect 26252 29850 26280 30126
rect 26240 29844 26292 29850
rect 26240 29786 26292 29792
rect 26712 29646 26740 30534
rect 26896 29646 26924 32166
rect 26988 31890 27016 32370
rect 27632 32026 27660 34200
rect 29196 32502 29224 34200
rect 29184 32496 29236 32502
rect 29184 32438 29236 32444
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 27620 32020 27672 32026
rect 27620 31962 27672 31968
rect 28184 31890 28212 32370
rect 29000 32360 29052 32366
rect 29000 32302 29052 32308
rect 30380 32360 30432 32366
rect 30380 32302 30432 32308
rect 26976 31884 27028 31890
rect 26976 31826 27028 31832
rect 28172 31884 28224 31890
rect 28172 31826 28224 31832
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 27160 31680 27212 31686
rect 27160 31622 27212 31628
rect 26976 31136 27028 31142
rect 26976 31078 27028 31084
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 26700 29640 26752 29646
rect 26700 29582 26752 29588
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 25514 29404 25822 29413
rect 25514 29402 25520 29404
rect 25576 29402 25600 29404
rect 25656 29402 25680 29404
rect 25736 29402 25760 29404
rect 25816 29402 25822 29404
rect 25576 29350 25578 29402
rect 25758 29350 25760 29402
rect 25514 29348 25520 29350
rect 25576 29348 25600 29350
rect 25656 29348 25680 29350
rect 25736 29348 25760 29350
rect 25816 29348 25822 29350
rect 25514 29339 25822 29348
rect 26988 29170 27016 31078
rect 27172 30666 27200 31622
rect 27434 31376 27490 31385
rect 27434 31311 27490 31320
rect 27448 30802 27476 31311
rect 27436 30796 27488 30802
rect 27436 30738 27488 30744
rect 27160 30660 27212 30666
rect 27160 30602 27212 30608
rect 27436 30660 27488 30666
rect 27436 30602 27488 30608
rect 27448 30190 27476 30602
rect 27632 30394 27660 31758
rect 28540 31680 28592 31686
rect 28540 31622 28592 31628
rect 28264 31340 28316 31346
rect 28264 31282 28316 31288
rect 28448 31340 28500 31346
rect 28448 31282 28500 31288
rect 28080 30728 28132 30734
rect 28080 30670 28132 30676
rect 27620 30388 27672 30394
rect 27620 30330 27672 30336
rect 27436 30184 27488 30190
rect 27436 30126 27488 30132
rect 27988 30184 28040 30190
rect 27988 30126 28040 30132
rect 27344 30116 27396 30122
rect 27344 30058 27396 30064
rect 27356 29646 27384 30058
rect 27344 29640 27396 29646
rect 27344 29582 27396 29588
rect 28000 29186 28028 30126
rect 28092 29306 28120 30670
rect 28172 30388 28224 30394
rect 28172 30330 28224 30336
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 26976 29164 27028 29170
rect 28000 29158 28120 29186
rect 26976 29106 27028 29112
rect 26792 29096 26844 29102
rect 26792 29038 26844 29044
rect 24952 28552 25004 28558
rect 24952 28494 25004 28500
rect 25514 28316 25822 28325
rect 25514 28314 25520 28316
rect 25576 28314 25600 28316
rect 25656 28314 25680 28316
rect 25736 28314 25760 28316
rect 25816 28314 25822 28316
rect 25576 28262 25578 28314
rect 25758 28262 25760 28314
rect 25514 28260 25520 28262
rect 25576 28260 25600 28262
rect 25656 28260 25680 28262
rect 25736 28260 25760 28262
rect 25816 28260 25822 28262
rect 25514 28251 25822 28260
rect 26804 28218 26832 29038
rect 28092 28966 28120 29158
rect 27160 28960 27212 28966
rect 27160 28902 27212 28908
rect 28080 28960 28132 28966
rect 28080 28902 28132 28908
rect 26792 28212 26844 28218
rect 26792 28154 26844 28160
rect 26884 27872 26936 27878
rect 26884 27814 26936 27820
rect 24860 27600 24912 27606
rect 24860 27542 24912 27548
rect 26896 27402 26924 27814
rect 27172 27606 27200 28902
rect 27988 28552 28040 28558
rect 27988 28494 28040 28500
rect 27712 28416 27764 28422
rect 27712 28358 27764 28364
rect 27896 28416 27948 28422
rect 27896 28358 27948 28364
rect 27160 27600 27212 27606
rect 27160 27542 27212 27548
rect 26884 27396 26936 27402
rect 26884 27338 26936 27344
rect 17326 27228 17634 27237
rect 17326 27226 17332 27228
rect 17388 27226 17412 27228
rect 17468 27226 17492 27228
rect 17548 27226 17572 27228
rect 17628 27226 17634 27228
rect 17388 27174 17390 27226
rect 17570 27174 17572 27226
rect 17326 27172 17332 27174
rect 17388 27172 17412 27174
rect 17468 27172 17492 27174
rect 17548 27172 17572 27174
rect 17628 27172 17634 27174
rect 17326 27163 17634 27172
rect 25514 27228 25822 27237
rect 25514 27226 25520 27228
rect 25576 27226 25600 27228
rect 25656 27226 25680 27228
rect 25736 27226 25760 27228
rect 25816 27226 25822 27228
rect 25576 27174 25578 27226
rect 25758 27174 25760 27226
rect 25514 27172 25520 27174
rect 25576 27172 25600 27174
rect 25656 27172 25680 27174
rect 25736 27172 25760 27174
rect 25816 27172 25822 27174
rect 25514 27163 25822 27172
rect 26896 26926 26924 27338
rect 27724 26994 27752 28358
rect 27908 28082 27936 28358
rect 27896 28076 27948 28082
rect 27896 28018 27948 28024
rect 28000 27946 28028 28494
rect 27988 27940 28040 27946
rect 27988 27882 28040 27888
rect 28092 27402 28120 28902
rect 28184 27538 28212 30330
rect 28276 29782 28304 31282
rect 28460 29850 28488 31282
rect 28448 29844 28500 29850
rect 28448 29786 28500 29792
rect 28264 29776 28316 29782
rect 28264 29718 28316 29724
rect 28356 27600 28408 27606
rect 28356 27542 28408 27548
rect 28172 27532 28224 27538
rect 28172 27474 28224 27480
rect 28080 27396 28132 27402
rect 28080 27338 28132 27344
rect 27988 27328 28040 27334
rect 27988 27270 28040 27276
rect 28000 26994 28028 27270
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27988 26988 28040 26994
rect 27988 26930 28040 26936
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 27804 26920 27856 26926
rect 27804 26862 27856 26868
rect 27620 26852 27672 26858
rect 27620 26794 27672 26800
rect 21420 26684 21728 26693
rect 21420 26682 21426 26684
rect 21482 26682 21506 26684
rect 21562 26682 21586 26684
rect 21642 26682 21666 26684
rect 21722 26682 21728 26684
rect 21482 26630 21484 26682
rect 21664 26630 21666 26682
rect 21420 26628 21426 26630
rect 21482 26628 21506 26630
rect 21562 26628 21586 26630
rect 21642 26628 21666 26630
rect 21722 26628 21728 26630
rect 21420 26619 21728 26628
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 17326 26140 17634 26149
rect 17326 26138 17332 26140
rect 17388 26138 17412 26140
rect 17468 26138 17492 26140
rect 17548 26138 17572 26140
rect 17628 26138 17634 26140
rect 17388 26086 17390 26138
rect 17570 26086 17572 26138
rect 17326 26084 17332 26086
rect 17388 26084 17412 26086
rect 17468 26084 17492 26086
rect 17548 26084 17572 26086
rect 17628 26084 17634 26086
rect 17326 26075 17634 26084
rect 17132 26036 17184 26042
rect 17132 25978 17184 25984
rect 16764 25832 16816 25838
rect 16764 25774 16816 25780
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 15764 24614 15792 24754
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 15752 24608 15804 24614
rect 15752 24550 15804 24556
rect 9138 23964 9446 23973
rect 9138 23962 9144 23964
rect 9200 23962 9224 23964
rect 9280 23962 9304 23964
rect 9360 23962 9384 23964
rect 9440 23962 9446 23964
rect 9200 23910 9202 23962
rect 9382 23910 9384 23962
rect 9138 23908 9144 23910
rect 9200 23908 9224 23910
rect 9280 23908 9304 23910
rect 9360 23908 9384 23910
rect 9440 23908 9446 23910
rect 9138 23899 9446 23908
rect 13096 23866 13124 24550
rect 13232 24508 13540 24517
rect 13232 24506 13238 24508
rect 13294 24506 13318 24508
rect 13374 24506 13398 24508
rect 13454 24506 13478 24508
rect 13534 24506 13540 24508
rect 13294 24454 13296 24506
rect 13476 24454 13478 24506
rect 13232 24452 13238 24454
rect 13294 24452 13318 24454
rect 13374 24452 13398 24454
rect 13454 24452 13478 24454
rect 13534 24452 13540 24454
rect 13232 24443 13540 24452
rect 15764 24410 15792 24550
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9138 22876 9446 22885
rect 9138 22874 9144 22876
rect 9200 22874 9224 22876
rect 9280 22874 9304 22876
rect 9360 22874 9384 22876
rect 9440 22874 9446 22876
rect 9200 22822 9202 22874
rect 9382 22822 9384 22874
rect 9138 22820 9144 22822
rect 9200 22820 9224 22822
rect 9280 22820 9304 22822
rect 9360 22820 9384 22822
rect 9440 22820 9446 22822
rect 9138 22811 9446 22820
rect 9138 21788 9446 21797
rect 9138 21786 9144 21788
rect 9200 21786 9224 21788
rect 9280 21786 9304 21788
rect 9360 21786 9384 21788
rect 9440 21786 9446 21788
rect 9200 21734 9202 21786
rect 9382 21734 9384 21786
rect 9138 21732 9144 21734
rect 9200 21732 9224 21734
rect 9280 21732 9304 21734
rect 9360 21732 9384 21734
rect 9440 21732 9446 21734
rect 9138 21723 9446 21732
rect 9600 20806 9628 23462
rect 13232 23420 13540 23429
rect 13232 23418 13238 23420
rect 13294 23418 13318 23420
rect 13374 23418 13398 23420
rect 13454 23418 13478 23420
rect 13534 23418 13540 23420
rect 13294 23366 13296 23418
rect 13476 23366 13478 23418
rect 13232 23364 13238 23366
rect 13294 23364 13318 23366
rect 13374 23364 13398 23366
rect 13454 23364 13478 23366
rect 13534 23364 13540 23366
rect 13232 23355 13540 23364
rect 13232 22332 13540 22341
rect 13232 22330 13238 22332
rect 13294 22330 13318 22332
rect 13374 22330 13398 22332
rect 13454 22330 13478 22332
rect 13534 22330 13540 22332
rect 13294 22278 13296 22330
rect 13476 22278 13478 22330
rect 13232 22276 13238 22278
rect 13294 22276 13318 22278
rect 13374 22276 13398 22278
rect 13454 22276 13478 22278
rect 13534 22276 13540 22278
rect 13232 22267 13540 22276
rect 13232 21244 13540 21253
rect 13232 21242 13238 21244
rect 13294 21242 13318 21244
rect 13374 21242 13398 21244
rect 13454 21242 13478 21244
rect 13534 21242 13540 21244
rect 13294 21190 13296 21242
rect 13476 21190 13478 21242
rect 13232 21188 13238 21190
rect 13294 21188 13318 21190
rect 13374 21188 13398 21190
rect 13454 21188 13478 21190
rect 13534 21188 13540 21190
rect 13232 21179 13540 21188
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 9138 20700 9446 20709
rect 9138 20698 9144 20700
rect 9200 20698 9224 20700
rect 9280 20698 9304 20700
rect 9360 20698 9384 20700
rect 9440 20698 9446 20700
rect 9200 20646 9202 20698
rect 9382 20646 9384 20698
rect 9138 20644 9144 20646
rect 9200 20644 9224 20646
rect 9280 20644 9304 20646
rect 9360 20644 9384 20646
rect 9440 20644 9446 20646
rect 9138 20635 9446 20644
rect 9138 19612 9446 19621
rect 9138 19610 9144 19612
rect 9200 19610 9224 19612
rect 9280 19610 9304 19612
rect 9360 19610 9384 19612
rect 9440 19610 9446 19612
rect 9200 19558 9202 19610
rect 9382 19558 9384 19610
rect 9138 19556 9144 19558
rect 9200 19556 9224 19558
rect 9280 19556 9304 19558
rect 9360 19556 9384 19558
rect 9440 19556 9446 19558
rect 9138 19547 9446 19556
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4816 18222 4844 18770
rect 9138 18524 9446 18533
rect 9138 18522 9144 18524
rect 9200 18522 9224 18524
rect 9280 18522 9304 18524
rect 9360 18522 9384 18524
rect 9440 18522 9446 18524
rect 9200 18470 9202 18522
rect 9382 18470 9384 18522
rect 9138 18468 9144 18470
rect 9200 18468 9224 18470
rect 9280 18468 9304 18470
rect 9360 18468 9384 18470
rect 9440 18468 9446 18470
rect 9138 18459 9446 18468
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4816 17746 4844 18158
rect 5044 17980 5352 17989
rect 5044 17978 5050 17980
rect 5106 17978 5130 17980
rect 5186 17978 5210 17980
rect 5266 17978 5290 17980
rect 5346 17978 5352 17980
rect 5106 17926 5108 17978
rect 5288 17926 5290 17978
rect 5044 17924 5050 17926
rect 5106 17924 5130 17926
rect 5186 17924 5210 17926
rect 5266 17924 5290 17926
rect 5346 17924 5352 17926
rect 5044 17915 5352 17924
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 10336 17678 10364 20742
rect 13232 20156 13540 20165
rect 13232 20154 13238 20156
rect 13294 20154 13318 20156
rect 13374 20154 13398 20156
rect 13454 20154 13478 20156
rect 13534 20154 13540 20156
rect 13294 20102 13296 20154
rect 13476 20102 13478 20154
rect 13232 20100 13238 20102
rect 13294 20100 13318 20102
rect 13374 20100 13398 20102
rect 13454 20100 13478 20102
rect 13534 20100 13540 20102
rect 13232 20091 13540 20100
rect 13232 19068 13540 19077
rect 13232 19066 13238 19068
rect 13294 19066 13318 19068
rect 13374 19066 13398 19068
rect 13454 19066 13478 19068
rect 13534 19066 13540 19068
rect 13294 19014 13296 19066
rect 13476 19014 13478 19066
rect 13232 19012 13238 19014
rect 13294 19012 13318 19014
rect 13374 19012 13398 19014
rect 13454 19012 13478 19014
rect 13534 19012 13540 19014
rect 13232 19003 13540 19012
rect 13232 17980 13540 17989
rect 13232 17978 13238 17980
rect 13294 17978 13318 17980
rect 13374 17978 13398 17980
rect 13454 17978 13478 17980
rect 13534 17978 13540 17980
rect 13294 17926 13296 17978
rect 13476 17926 13478 17978
rect 13232 17924 13238 17926
rect 13294 17924 13318 17926
rect 13374 17924 13398 17926
rect 13454 17924 13478 17926
rect 13534 17924 13540 17926
rect 13232 17915 13540 17924
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 9138 17436 9446 17445
rect 9138 17434 9144 17436
rect 9200 17434 9224 17436
rect 9280 17434 9304 17436
rect 9360 17434 9384 17436
rect 9440 17434 9446 17436
rect 9200 17382 9202 17434
rect 9382 17382 9384 17434
rect 9138 17380 9144 17382
rect 9200 17380 9224 17382
rect 9280 17380 9304 17382
rect 9360 17380 9384 17382
rect 9440 17380 9446 17382
rect 9138 17371 9446 17380
rect 4528 17332 4580 17338
rect 4528 17274 4580 17280
rect 4528 17128 4580 17134
rect 4528 17070 4580 17076
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 16250 4384 16526
rect 4540 16454 4568 17070
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 5044 16892 5352 16901
rect 5044 16890 5050 16892
rect 5106 16890 5130 16892
rect 5186 16890 5210 16892
rect 5266 16890 5290 16892
rect 5346 16890 5352 16892
rect 5106 16838 5108 16890
rect 5288 16838 5290 16890
rect 5044 16836 5050 16838
rect 5106 16836 5130 16838
rect 5186 16836 5210 16838
rect 5266 16836 5290 16838
rect 5346 16836 5352 16838
rect 5044 16827 5352 16836
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4356 15706 4384 15982
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 3804 15162 3832 15438
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3712 14618 3740 14962
rect 3700 14612 3752 14618
rect 3700 14554 3752 14560
rect 3988 14550 4016 15370
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4356 14618 4384 14758
rect 4344 14612 4396 14618
rect 4344 14554 4396 14560
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4264 12986 4292 13262
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3988 12442 4016 12718
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 4264 12374 4292 12922
rect 4356 12918 4384 13670
rect 4448 13394 4476 14486
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4448 12918 4476 13330
rect 4344 12912 4396 12918
rect 4344 12854 4396 12860
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3804 11354 3832 12174
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4448 11898 4476 12038
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 4356 11218 4384 11494
rect 4540 11354 4568 12038
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10674 3832 10950
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 4356 10538 4384 11154
rect 4632 10674 4660 16662
rect 7484 16574 7512 17002
rect 7484 16546 7604 16574
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 14346 4844 16390
rect 4896 16108 4948 16114
rect 4896 16050 4948 16056
rect 4908 15706 4936 16050
rect 5044 15804 5352 15813
rect 5044 15802 5050 15804
rect 5106 15802 5130 15804
rect 5186 15802 5210 15804
rect 5266 15802 5290 15804
rect 5346 15802 5352 15804
rect 5106 15750 5108 15802
rect 5288 15750 5290 15802
rect 5044 15748 5050 15750
rect 5106 15748 5130 15750
rect 5186 15748 5210 15750
rect 5266 15748 5290 15750
rect 5346 15748 5352 15750
rect 5044 15739 5352 15748
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 7576 15502 7604 16546
rect 9138 16348 9446 16357
rect 9138 16346 9144 16348
rect 9200 16346 9224 16348
rect 9280 16346 9304 16348
rect 9360 16346 9384 16348
rect 9440 16346 9446 16348
rect 9200 16294 9202 16346
rect 9382 16294 9384 16346
rect 9138 16292 9144 16294
rect 9200 16292 9224 16294
rect 9280 16292 9304 16294
rect 9360 16292 9384 16294
rect 9440 16292 9446 16294
rect 9138 16283 9446 16292
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 9138 15260 9446 15269
rect 9138 15258 9144 15260
rect 9200 15258 9224 15260
rect 9280 15258 9304 15260
rect 9360 15258 9384 15260
rect 9440 15258 9446 15260
rect 9200 15206 9202 15258
rect 9382 15206 9384 15258
rect 9138 15204 9144 15206
rect 9200 15204 9224 15206
rect 9280 15204 9304 15206
rect 9360 15204 9384 15206
rect 9440 15204 9446 15206
rect 9138 15195 9446 15204
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5044 14716 5352 14725
rect 5044 14714 5050 14716
rect 5106 14714 5130 14716
rect 5186 14714 5210 14716
rect 5266 14714 5290 14716
rect 5346 14714 5352 14716
rect 5106 14662 5108 14714
rect 5288 14662 5290 14714
rect 5044 14660 5050 14662
rect 5106 14660 5130 14662
rect 5186 14660 5210 14662
rect 5266 14660 5290 14662
rect 5346 14660 5352 14662
rect 5044 14651 5352 14660
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4816 13734 4844 14282
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 12646 4844 13670
rect 5044 13628 5352 13637
rect 5044 13626 5050 13628
rect 5106 13626 5130 13628
rect 5186 13626 5210 13628
rect 5266 13626 5290 13628
rect 5346 13626 5352 13628
rect 5106 13574 5108 13626
rect 5288 13574 5290 13626
rect 5044 13572 5050 13574
rect 5106 13572 5130 13574
rect 5186 13572 5210 13574
rect 5266 13572 5290 13574
rect 5346 13572 5352 13574
rect 5044 13563 5352 13572
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4816 12170 4844 12582
rect 5044 12540 5352 12549
rect 5044 12538 5050 12540
rect 5106 12538 5130 12540
rect 5186 12538 5210 12540
rect 5266 12538 5290 12540
rect 5346 12538 5352 12540
rect 5106 12486 5108 12538
rect 5288 12486 5290 12538
rect 5044 12484 5050 12486
rect 5106 12484 5130 12486
rect 5186 12484 5210 12486
rect 5266 12484 5290 12486
rect 5346 12484 5352 12486
rect 5044 12475 5352 12484
rect 5460 12306 5488 14758
rect 9138 14172 9446 14181
rect 9138 14170 9144 14172
rect 9200 14170 9224 14172
rect 9280 14170 9304 14172
rect 9360 14170 9384 14172
rect 9440 14170 9446 14172
rect 9200 14118 9202 14170
rect 9382 14118 9384 14170
rect 9138 14116 9144 14118
rect 9200 14116 9224 14118
rect 9280 14116 9304 14118
rect 9360 14116 9384 14118
rect 9440 14116 9446 14118
rect 9138 14107 9446 14116
rect 9138 13084 9446 13093
rect 9138 13082 9144 13084
rect 9200 13082 9224 13084
rect 9280 13082 9304 13084
rect 9360 13082 9384 13084
rect 9440 13082 9446 13084
rect 9200 13030 9202 13082
rect 9382 13030 9384 13082
rect 9138 13028 9144 13030
rect 9200 13028 9224 13030
rect 9280 13028 9304 13030
rect 9360 13028 9384 13030
rect 9440 13028 9446 13030
rect 9138 13019 9446 13028
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4344 10532 4396 10538
rect 4344 10474 4396 10480
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 3712 10062 3740 10406
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 8634 3648 9318
rect 3804 8974 3832 9862
rect 4356 9518 4384 9998
rect 4344 9512 4396 9518
rect 4344 9454 4396 9460
rect 4356 9178 4384 9454
rect 4448 9382 4476 10406
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 4356 8362 4384 8910
rect 4448 8430 4476 9318
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 5370 3556 5646
rect 3620 5370 3648 7346
rect 3804 7002 3832 7822
rect 3792 6996 3844 7002
rect 3792 6938 3844 6944
rect 3988 6798 4016 8298
rect 4356 8090 4384 8298
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4172 6390 4200 7890
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 4264 4622 4292 6598
rect 4356 6338 4384 7754
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4448 7546 4476 7686
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4448 6866 4476 7142
rect 4632 6914 4660 10610
rect 4816 10606 4844 12106
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 5044 11452 5352 11461
rect 5044 11450 5050 11452
rect 5106 11450 5130 11452
rect 5186 11450 5210 11452
rect 5266 11450 5290 11452
rect 5346 11450 5352 11452
rect 5106 11398 5108 11450
rect 5288 11398 5290 11450
rect 5044 11396 5050 11398
rect 5106 11396 5130 11398
rect 5186 11396 5210 11398
rect 5266 11396 5290 11398
rect 5346 11396 5352 11398
rect 5044 11387 5352 11396
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 5044 10364 5352 10373
rect 5044 10362 5050 10364
rect 5106 10362 5130 10364
rect 5186 10362 5210 10364
rect 5266 10362 5290 10364
rect 5346 10362 5352 10364
rect 5106 10310 5108 10362
rect 5288 10310 5290 10362
rect 5044 10308 5050 10310
rect 5106 10308 5130 10310
rect 5186 10308 5210 10310
rect 5266 10308 5290 10310
rect 5346 10308 5352 10310
rect 5044 10299 5352 10308
rect 5044 9276 5352 9285
rect 5044 9274 5050 9276
rect 5106 9274 5130 9276
rect 5186 9274 5210 9276
rect 5266 9274 5290 9276
rect 5346 9274 5352 9276
rect 5106 9222 5108 9274
rect 5288 9222 5290 9274
rect 5044 9220 5050 9222
rect 5106 9220 5130 9222
rect 5186 9220 5210 9222
rect 5266 9220 5290 9222
rect 5346 9220 5352 9222
rect 5044 9211 5352 9220
rect 6012 9042 6040 12038
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7852 10266 7880 10678
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4724 7206 4752 7958
rect 4816 7818 4844 8230
rect 5044 8188 5352 8197
rect 5044 8186 5050 8188
rect 5106 8186 5130 8188
rect 5186 8186 5210 8188
rect 5266 8186 5290 8188
rect 5346 8186 5352 8188
rect 5106 8134 5108 8186
rect 5288 8134 5290 8186
rect 5044 8132 5050 8134
rect 5106 8132 5130 8134
rect 5186 8132 5210 8134
rect 5266 8132 5290 8134
rect 5346 8132 5352 8134
rect 5044 8123 5352 8132
rect 4804 7812 4856 7818
rect 4804 7754 4856 7760
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 5044 7100 5352 7109
rect 5044 7098 5050 7100
rect 5106 7098 5130 7100
rect 5186 7098 5210 7100
rect 5266 7098 5290 7100
rect 5346 7098 5352 7100
rect 5106 7046 5108 7098
rect 5288 7046 5290 7098
rect 5044 7044 5050 7046
rect 5106 7044 5130 7046
rect 5186 7044 5210 7046
rect 5266 7044 5290 7046
rect 5346 7044 5352 7046
rect 5044 7035 5352 7044
rect 4632 6886 4752 6914
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4356 6310 4476 6338
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4356 5914 4384 6190
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4448 5234 4476 6310
rect 4540 5914 4568 6734
rect 4724 6458 4752 6886
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 5044 6012 5352 6021
rect 5044 6010 5050 6012
rect 5106 6010 5130 6012
rect 5186 6010 5210 6012
rect 5266 6010 5290 6012
rect 5346 6010 5352 6012
rect 5106 5958 5108 6010
rect 5288 5958 5290 6010
rect 5044 5956 5050 5958
rect 5106 5956 5130 5958
rect 5186 5956 5210 5958
rect 5266 5956 5290 5958
rect 5346 5956 5352 5958
rect 5044 5947 5352 5956
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4448 5030 4476 5170
rect 4540 5098 4568 5850
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8772 5302 8800 5578
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 4528 5092 4580 5098
rect 4528 5034 4580 5040
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4448 4826 4476 4966
rect 5044 4924 5352 4933
rect 5044 4922 5050 4924
rect 5106 4922 5130 4924
rect 5186 4922 5210 4924
rect 5266 4922 5290 4924
rect 5346 4922 5352 4924
rect 5106 4870 5108 4922
rect 5288 4870 5290 4922
rect 5044 4868 5050 4870
rect 5106 4868 5130 4870
rect 5186 4868 5210 4870
rect 5266 4868 5290 4870
rect 5346 4868 5352 4870
rect 5044 4859 5352 4868
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 8312 4758 8340 5102
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8404 4622 8432 5238
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8496 4826 8524 5034
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8588 4826 8616 4966
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 5044 3836 5352 3845
rect 5044 3834 5050 3836
rect 5106 3834 5130 3836
rect 5186 3834 5210 3836
rect 5266 3834 5290 3836
rect 5346 3834 5352 3836
rect 5106 3782 5108 3834
rect 5288 3782 5290 3834
rect 5044 3780 5050 3782
rect 5106 3780 5130 3782
rect 5186 3780 5210 3782
rect 5266 3780 5290 3782
rect 5346 3780 5352 3782
rect 5044 3771 5352 3780
rect 6656 3602 6684 3878
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6012 3058 6040 3334
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 2596 2984 2648 2990
rect 4988 2984 5040 2990
rect 2596 2926 2648 2932
rect 4908 2932 4988 2938
rect 4908 2926 5040 2932
rect 1582 2816 1638 2825
rect 1582 2751 1638 2760
rect 1596 2514 1624 2751
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 848 2372 900 2378
rect 848 2314 900 2320
rect 860 800 888 2314
rect 2240 870 2360 898
rect 2240 800 2268 870
rect 846 0 902 800
rect 2226 0 2282 800
rect 2332 762 2360 870
rect 2516 762 2544 2518
rect 2608 2446 2636 2926
rect 4908 2910 5028 2926
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3804 1306 3832 2382
rect 4908 1578 4936 2910
rect 5044 2748 5352 2757
rect 5044 2746 5050 2748
rect 5106 2746 5130 2748
rect 5186 2746 5210 2748
rect 5266 2746 5290 2748
rect 5346 2746 5352 2748
rect 5106 2694 5108 2746
rect 5288 2694 5290 2746
rect 5044 2692 5050 2694
rect 5106 2692 5130 2694
rect 5186 2692 5210 2694
rect 5266 2692 5290 2694
rect 5346 2692 5352 2694
rect 5044 2683 5352 2692
rect 4908 1550 5028 1578
rect 3620 1278 3832 1306
rect 3620 800 3648 1278
rect 5000 800 5028 1550
rect 6380 870 6500 898
rect 6380 800 6408 870
rect 2332 734 2544 762
rect 3606 0 3662 800
rect 4986 0 5042 800
rect 6366 0 6422 800
rect 6472 762 6500 870
rect 6748 762 6776 4014
rect 7760 800 7788 4014
rect 7852 2514 7880 4082
rect 8680 3534 8708 4966
rect 8772 4826 8800 4966
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 7840 2508 7892 2514
rect 7840 2450 7892 2456
rect 8128 2446 8156 3334
rect 8312 3194 8340 3402
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8864 3074 8892 5714
rect 8956 3738 8984 12038
rect 9138 11996 9446 12005
rect 9138 11994 9144 11996
rect 9200 11994 9224 11996
rect 9280 11994 9304 11996
rect 9360 11994 9384 11996
rect 9440 11994 9446 11996
rect 9200 11942 9202 11994
rect 9382 11942 9384 11994
rect 9138 11940 9144 11942
rect 9200 11940 9224 11942
rect 9280 11940 9304 11942
rect 9360 11940 9384 11942
rect 9440 11940 9446 11942
rect 9138 11931 9446 11940
rect 9138 10908 9446 10917
rect 9138 10906 9144 10908
rect 9200 10906 9224 10908
rect 9280 10906 9304 10908
rect 9360 10906 9384 10908
rect 9440 10906 9446 10908
rect 9200 10854 9202 10906
rect 9382 10854 9384 10906
rect 9138 10852 9144 10854
rect 9200 10852 9224 10854
rect 9280 10852 9304 10854
rect 9360 10852 9384 10854
rect 9440 10852 9446 10854
rect 9138 10843 9446 10852
rect 9138 9820 9446 9829
rect 9138 9818 9144 9820
rect 9200 9818 9224 9820
rect 9280 9818 9304 9820
rect 9360 9818 9384 9820
rect 9440 9818 9446 9820
rect 9200 9766 9202 9818
rect 9382 9766 9384 9818
rect 9138 9764 9144 9766
rect 9200 9764 9224 9766
rect 9280 9764 9304 9766
rect 9360 9764 9384 9766
rect 9440 9764 9446 9766
rect 9138 9755 9446 9764
rect 9508 9178 9536 12174
rect 10336 10810 10364 17614
rect 13232 16892 13540 16901
rect 13232 16890 13238 16892
rect 13294 16890 13318 16892
rect 13374 16890 13398 16892
rect 13454 16890 13478 16892
rect 13534 16890 13540 16892
rect 13294 16838 13296 16890
rect 13476 16838 13478 16890
rect 13232 16836 13238 16838
rect 13294 16836 13318 16838
rect 13374 16836 13398 16838
rect 13454 16836 13478 16838
rect 13534 16836 13540 16838
rect 13232 16827 13540 16836
rect 13232 15804 13540 15813
rect 13232 15802 13238 15804
rect 13294 15802 13318 15804
rect 13374 15802 13398 15804
rect 13454 15802 13478 15804
rect 13534 15802 13540 15804
rect 13294 15750 13296 15802
rect 13476 15750 13478 15802
rect 13232 15748 13238 15750
rect 13294 15748 13318 15750
rect 13374 15748 13398 15750
rect 13454 15748 13478 15750
rect 13534 15748 13540 15750
rect 13232 15739 13540 15748
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10612 13462 10640 15438
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11624 14618 11652 14962
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 11830 11192 13126
rect 11440 12238 11468 14486
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 13190 12020 14214
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 12728 11762 12756 14894
rect 13232 14716 13540 14725
rect 13232 14714 13238 14716
rect 13294 14714 13318 14716
rect 13374 14714 13398 14716
rect 13454 14714 13478 14716
rect 13534 14714 13540 14716
rect 13294 14662 13296 14714
rect 13476 14662 13478 14714
rect 13232 14660 13238 14662
rect 13294 14660 13318 14662
rect 13374 14660 13398 14662
rect 13454 14660 13478 14662
rect 13534 14660 13540 14662
rect 13232 14651 13540 14660
rect 15948 13870 15976 24754
rect 16776 24750 16804 25774
rect 17326 25052 17634 25061
rect 17326 25050 17332 25052
rect 17388 25050 17412 25052
rect 17468 25050 17492 25052
rect 17548 25050 17572 25052
rect 17628 25050 17634 25052
rect 17388 24998 17390 25050
rect 17570 24998 17572 25050
rect 17326 24996 17332 24998
rect 17388 24996 17412 24998
rect 17468 24996 17492 24998
rect 17548 24996 17572 24998
rect 17628 24996 17634 24998
rect 17326 24987 17634 24996
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 17326 23964 17634 23973
rect 17326 23962 17332 23964
rect 17388 23962 17412 23964
rect 17468 23962 17492 23964
rect 17548 23962 17572 23964
rect 17628 23962 17634 23964
rect 17388 23910 17390 23962
rect 17570 23910 17572 23962
rect 17326 23908 17332 23910
rect 17388 23908 17412 23910
rect 17468 23908 17492 23910
rect 17548 23908 17572 23910
rect 17628 23908 17634 23910
rect 17326 23899 17634 23908
rect 18156 23322 18184 26318
rect 25514 26140 25822 26149
rect 25514 26138 25520 26140
rect 25576 26138 25600 26140
rect 25656 26138 25680 26140
rect 25736 26138 25760 26140
rect 25816 26138 25822 26140
rect 25576 26086 25578 26138
rect 25758 26086 25760 26138
rect 25514 26084 25520 26086
rect 25576 26084 25600 26086
rect 25656 26084 25680 26086
rect 25736 26084 25760 26086
rect 25816 26084 25822 26086
rect 25514 26075 25822 26084
rect 21420 25596 21728 25605
rect 21420 25594 21426 25596
rect 21482 25594 21506 25596
rect 21562 25594 21586 25596
rect 21642 25594 21666 25596
rect 21722 25594 21728 25596
rect 21482 25542 21484 25594
rect 21664 25542 21666 25594
rect 21420 25540 21426 25542
rect 21482 25540 21506 25542
rect 21562 25540 21586 25542
rect 21642 25540 21666 25542
rect 21722 25540 21728 25542
rect 21420 25531 21728 25540
rect 26976 25356 27028 25362
rect 26976 25298 27028 25304
rect 25514 25052 25822 25061
rect 25514 25050 25520 25052
rect 25576 25050 25600 25052
rect 25656 25050 25680 25052
rect 25736 25050 25760 25052
rect 25816 25050 25822 25052
rect 25576 24998 25578 25050
rect 25758 24998 25760 25050
rect 25514 24996 25520 24998
rect 25576 24996 25600 24998
rect 25656 24996 25680 24998
rect 25736 24996 25760 24998
rect 25816 24996 25822 24998
rect 25514 24987 25822 24996
rect 21420 24508 21728 24517
rect 21420 24506 21426 24508
rect 21482 24506 21506 24508
rect 21562 24506 21586 24508
rect 21642 24506 21666 24508
rect 21722 24506 21728 24508
rect 21482 24454 21484 24506
rect 21664 24454 21666 24506
rect 21420 24452 21426 24454
rect 21482 24452 21506 24454
rect 21562 24452 21586 24454
rect 21642 24452 21666 24454
rect 21722 24452 21728 24454
rect 21420 24443 21728 24452
rect 25514 23964 25822 23973
rect 25514 23962 25520 23964
rect 25576 23962 25600 23964
rect 25656 23962 25680 23964
rect 25736 23962 25760 23964
rect 25816 23962 25822 23964
rect 25576 23910 25578 23962
rect 25758 23910 25760 23962
rect 25514 23908 25520 23910
rect 25576 23908 25600 23910
rect 25656 23908 25680 23910
rect 25736 23908 25760 23910
rect 25816 23908 25822 23910
rect 25514 23899 25822 23908
rect 25412 23656 25464 23662
rect 25412 23598 25464 23604
rect 21420 23420 21728 23429
rect 21420 23418 21426 23420
rect 21482 23418 21506 23420
rect 21562 23418 21586 23420
rect 21642 23418 21666 23420
rect 21722 23418 21728 23420
rect 21482 23366 21484 23418
rect 21664 23366 21666 23418
rect 21420 23364 21426 23366
rect 21482 23364 21506 23366
rect 21562 23364 21586 23366
rect 21642 23364 21666 23366
rect 21722 23364 21728 23366
rect 21420 23355 21728 23364
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 17224 23112 17276 23118
rect 17224 23054 17276 23060
rect 17236 20058 17264 23054
rect 17326 22876 17634 22885
rect 17326 22874 17332 22876
rect 17388 22874 17412 22876
rect 17468 22874 17492 22876
rect 17548 22874 17572 22876
rect 17628 22874 17634 22876
rect 17388 22822 17390 22874
rect 17570 22822 17572 22874
rect 17326 22820 17332 22822
rect 17388 22820 17412 22822
rect 17468 22820 17492 22822
rect 17548 22820 17572 22822
rect 17628 22820 17634 22822
rect 17326 22811 17634 22820
rect 21420 22332 21728 22341
rect 21420 22330 21426 22332
rect 21482 22330 21506 22332
rect 21562 22330 21586 22332
rect 21642 22330 21666 22332
rect 21722 22330 21728 22332
rect 21482 22278 21484 22330
rect 21664 22278 21666 22330
rect 21420 22276 21426 22278
rect 21482 22276 21506 22278
rect 21562 22276 21586 22278
rect 21642 22276 21666 22278
rect 21722 22276 21728 22278
rect 21420 22267 21728 22276
rect 17326 21788 17634 21797
rect 17326 21786 17332 21788
rect 17388 21786 17412 21788
rect 17468 21786 17492 21788
rect 17548 21786 17572 21788
rect 17628 21786 17634 21788
rect 17388 21734 17390 21786
rect 17570 21734 17572 21786
rect 17326 21732 17332 21734
rect 17388 21732 17412 21734
rect 17468 21732 17492 21734
rect 17548 21732 17572 21734
rect 17628 21732 17634 21734
rect 17326 21723 17634 21732
rect 21420 21244 21728 21253
rect 21420 21242 21426 21244
rect 21482 21242 21506 21244
rect 21562 21242 21586 21244
rect 21642 21242 21666 21244
rect 21722 21242 21728 21244
rect 21482 21190 21484 21242
rect 21664 21190 21666 21242
rect 21420 21188 21426 21190
rect 21482 21188 21506 21190
rect 21562 21188 21586 21190
rect 21642 21188 21666 21190
rect 21722 21188 21728 21190
rect 21420 21179 21728 21188
rect 25424 21146 25452 23598
rect 25872 23520 25924 23526
rect 25872 23462 25924 23468
rect 25884 22982 25912 23462
rect 26988 23322 27016 25298
rect 27632 23866 27660 26794
rect 27816 26314 27844 26862
rect 28092 26450 28120 27338
rect 28368 27130 28396 27542
rect 28356 27124 28408 27130
rect 28356 27066 28408 27072
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 27804 26308 27856 26314
rect 27804 26250 27856 26256
rect 28552 25362 28580 31622
rect 29012 31482 29040 32302
rect 29608 32124 29916 32133
rect 29608 32122 29614 32124
rect 29670 32122 29694 32124
rect 29750 32122 29774 32124
rect 29830 32122 29854 32124
rect 29910 32122 29916 32124
rect 29670 32070 29672 32122
rect 29852 32070 29854 32122
rect 29608 32068 29614 32070
rect 29670 32068 29694 32070
rect 29750 32068 29774 32070
rect 29830 32068 29854 32070
rect 29910 32068 29916 32070
rect 29608 32059 29916 32068
rect 29092 31816 29144 31822
rect 29092 31758 29144 31764
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 29104 31346 29132 31758
rect 30196 31680 30248 31686
rect 30196 31622 30248 31628
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 29276 31340 29328 31346
rect 29276 31282 29328 31288
rect 29092 31136 29144 31142
rect 29092 31078 29144 31084
rect 28908 30660 28960 30666
rect 28908 30602 28960 30608
rect 28632 29572 28684 29578
rect 28632 29514 28684 29520
rect 28724 29572 28776 29578
rect 28724 29514 28776 29520
rect 28644 27470 28672 29514
rect 28736 28966 28764 29514
rect 28724 28960 28776 28966
rect 28724 28902 28776 28908
rect 28724 28552 28776 28558
rect 28724 28494 28776 28500
rect 28736 27470 28764 28494
rect 28920 27674 28948 30602
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 29012 29714 29040 30194
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 29104 29170 29132 31078
rect 29184 30184 29236 30190
rect 29184 30126 29236 30132
rect 29196 29170 29224 30126
rect 29288 30054 29316 31282
rect 29608 31036 29916 31045
rect 29608 31034 29614 31036
rect 29670 31034 29694 31036
rect 29750 31034 29774 31036
rect 29830 31034 29854 31036
rect 29910 31034 29916 31036
rect 29670 30982 29672 31034
rect 29852 30982 29854 31034
rect 29608 30980 29614 30982
rect 29670 30980 29694 30982
rect 29750 30980 29774 30982
rect 29830 30980 29854 30982
rect 29910 30980 29916 30982
rect 29608 30971 29916 30980
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 30104 30252 30156 30258
rect 30104 30194 30156 30200
rect 29276 30048 29328 30054
rect 29276 29990 29328 29996
rect 29368 30048 29420 30054
rect 29368 29990 29420 29996
rect 29380 29578 29408 29990
rect 29608 29948 29916 29957
rect 29608 29946 29614 29948
rect 29670 29946 29694 29948
rect 29750 29946 29774 29948
rect 29830 29946 29854 29948
rect 29910 29946 29916 29948
rect 29670 29894 29672 29946
rect 29852 29894 29854 29946
rect 29608 29892 29614 29894
rect 29670 29892 29694 29894
rect 29750 29892 29774 29894
rect 29830 29892 29854 29894
rect 29910 29892 29916 29894
rect 29608 29883 29916 29892
rect 29368 29572 29420 29578
rect 29368 29514 29420 29520
rect 29276 29504 29328 29510
rect 29276 29446 29328 29452
rect 29460 29504 29512 29510
rect 29460 29446 29512 29452
rect 29092 29164 29144 29170
rect 29092 29106 29144 29112
rect 29184 29164 29236 29170
rect 29184 29106 29236 29112
rect 29184 28008 29236 28014
rect 29184 27950 29236 27956
rect 28908 27668 28960 27674
rect 28908 27610 28960 27616
rect 28632 27464 28684 27470
rect 28632 27406 28684 27412
rect 28724 27464 28776 27470
rect 28724 27406 28776 27412
rect 29092 26920 29144 26926
rect 29092 26862 29144 26868
rect 29104 26518 29132 26862
rect 29092 26512 29144 26518
rect 29092 26454 29144 26460
rect 28816 26240 28868 26246
rect 28816 26182 28868 26188
rect 28828 25838 28856 26182
rect 28816 25832 28868 25838
rect 28816 25774 28868 25780
rect 29196 25498 29224 27950
rect 29288 27470 29316 29446
rect 29368 29028 29420 29034
rect 29368 28970 29420 28976
rect 29276 27464 29328 27470
rect 29276 27406 29328 27412
rect 29380 26586 29408 28970
rect 29472 28082 29500 29446
rect 29608 28860 29916 28869
rect 29608 28858 29614 28860
rect 29670 28858 29694 28860
rect 29750 28858 29774 28860
rect 29830 28858 29854 28860
rect 29910 28858 29916 28860
rect 29670 28806 29672 28858
rect 29852 28806 29854 28858
rect 29608 28804 29614 28806
rect 29670 28804 29694 28806
rect 29750 28804 29774 28806
rect 29830 28804 29854 28806
rect 29910 28804 29916 28806
rect 29608 28795 29916 28804
rect 29920 28416 29972 28422
rect 29920 28358 29972 28364
rect 29932 28082 29960 28358
rect 29460 28076 29512 28082
rect 29460 28018 29512 28024
rect 29920 28076 29972 28082
rect 29920 28018 29972 28024
rect 29608 27772 29916 27781
rect 29608 27770 29614 27772
rect 29670 27770 29694 27772
rect 29750 27770 29774 27772
rect 29830 27770 29854 27772
rect 29910 27770 29916 27772
rect 29670 27718 29672 27770
rect 29852 27718 29854 27770
rect 29608 27716 29614 27718
rect 29670 27716 29694 27718
rect 29750 27716 29774 27718
rect 29830 27716 29854 27718
rect 29910 27716 29916 27718
rect 29608 27707 29916 27716
rect 29552 27464 29604 27470
rect 29552 27406 29604 27412
rect 29564 26858 29592 27406
rect 30024 27130 30052 30194
rect 30116 28218 30144 30194
rect 30208 30054 30236 31622
rect 30196 30048 30248 30054
rect 30196 29990 30248 29996
rect 30288 29640 30340 29646
rect 30288 29582 30340 29588
rect 30196 29572 30248 29578
rect 30196 29514 30248 29520
rect 30104 28212 30156 28218
rect 30104 28154 30156 28160
rect 30104 27872 30156 27878
rect 30104 27814 30156 27820
rect 30012 27124 30064 27130
rect 30012 27066 30064 27072
rect 30116 26994 30144 27814
rect 30208 27130 30236 29514
rect 30300 27674 30328 29582
rect 30392 29102 30420 32302
rect 30472 30592 30524 30598
rect 30472 30534 30524 30540
rect 30380 29096 30432 29102
rect 30380 29038 30432 29044
rect 30288 27668 30340 27674
rect 30288 27610 30340 27616
rect 30484 27606 30512 30534
rect 30748 28960 30800 28966
rect 30748 28902 30800 28908
rect 30760 28626 30788 28902
rect 30852 28626 30880 34326
rect 32232 34326 32366 34354
rect 31298 33008 31354 33017
rect 31298 32943 31354 32952
rect 31024 32224 31076 32230
rect 31024 32166 31076 32172
rect 30932 31408 30984 31414
rect 30932 31350 30984 31356
rect 30944 30802 30972 31350
rect 30932 30796 30984 30802
rect 30932 30738 30984 30744
rect 30932 30184 30984 30190
rect 30932 30126 30984 30132
rect 30748 28620 30800 28626
rect 30748 28562 30800 28568
rect 30840 28620 30892 28626
rect 30840 28562 30892 28568
rect 30564 28552 30616 28558
rect 30564 28494 30616 28500
rect 30576 28218 30604 28494
rect 30564 28212 30616 28218
rect 30564 28154 30616 28160
rect 30472 27600 30524 27606
rect 30472 27542 30524 27548
rect 30196 27124 30248 27130
rect 30196 27066 30248 27072
rect 30944 26994 30972 30126
rect 31036 30122 31064 32166
rect 31116 30592 31168 30598
rect 31116 30534 31168 30540
rect 31024 30116 31076 30122
rect 31024 30058 31076 30064
rect 31128 29306 31156 30534
rect 31312 30326 31340 32943
rect 32128 32428 32180 32434
rect 32128 32370 32180 32376
rect 32140 31890 32168 32370
rect 32128 31884 32180 31890
rect 32128 31826 32180 31832
rect 31852 31680 31904 31686
rect 31852 31622 31904 31628
rect 31864 31414 31892 31622
rect 31852 31408 31904 31414
rect 31852 31350 31904 31356
rect 31576 31340 31628 31346
rect 31576 31282 31628 31288
rect 31484 31204 31536 31210
rect 31484 31146 31536 31152
rect 31392 30796 31444 30802
rect 31392 30738 31444 30744
rect 31300 30320 31352 30326
rect 31300 30262 31352 30268
rect 31404 29782 31432 30738
rect 31392 29776 31444 29782
rect 31392 29718 31444 29724
rect 31116 29300 31168 29306
rect 31116 29242 31168 29248
rect 31496 29186 31524 31146
rect 31404 29158 31524 29186
rect 31404 28014 31432 29158
rect 31484 29096 31536 29102
rect 31484 29038 31536 29044
rect 31496 28937 31524 29038
rect 31482 28928 31538 28937
rect 31482 28863 31538 28872
rect 31588 28762 31616 31282
rect 31852 31272 31904 31278
rect 31852 31214 31904 31220
rect 31576 28756 31628 28762
rect 31576 28698 31628 28704
rect 31864 28558 31892 31214
rect 32128 31136 32180 31142
rect 32128 31078 32180 31084
rect 32140 30666 32168 31078
rect 32036 30660 32088 30666
rect 32036 30602 32088 30608
rect 32128 30660 32180 30666
rect 32128 30602 32180 30608
rect 32048 30546 32076 30602
rect 32048 30518 32168 30546
rect 32140 30190 32168 30518
rect 32128 30184 32180 30190
rect 32128 30126 32180 30132
rect 32140 29578 32168 30126
rect 32128 29572 32180 29578
rect 32128 29514 32180 29520
rect 31944 29164 31996 29170
rect 31944 29106 31996 29112
rect 31956 28626 31984 29106
rect 32140 29102 32168 29514
rect 32128 29096 32180 29102
rect 32128 29038 32180 29044
rect 31944 28620 31996 28626
rect 31944 28562 31996 28568
rect 31852 28552 31904 28558
rect 31852 28494 31904 28500
rect 31944 28076 31996 28082
rect 31944 28018 31996 28024
rect 31392 28008 31444 28014
rect 31392 27950 31444 27956
rect 31484 28008 31536 28014
rect 31484 27950 31536 27956
rect 31668 28008 31720 28014
rect 31668 27950 31720 27956
rect 31496 27577 31524 27950
rect 31482 27568 31538 27577
rect 31482 27503 31538 27512
rect 30104 26988 30156 26994
rect 30104 26930 30156 26936
rect 30932 26988 30984 26994
rect 30932 26930 30984 26936
rect 29552 26852 29604 26858
rect 29552 26794 29604 26800
rect 29608 26684 29916 26693
rect 29608 26682 29614 26684
rect 29670 26682 29694 26684
rect 29750 26682 29774 26684
rect 29830 26682 29854 26684
rect 29910 26682 29916 26684
rect 29670 26630 29672 26682
rect 29852 26630 29854 26682
rect 29608 26628 29614 26630
rect 29670 26628 29694 26630
rect 29750 26628 29774 26630
rect 29830 26628 29854 26630
rect 29910 26628 29916 26630
rect 29608 26619 29916 26628
rect 29368 26580 29420 26586
rect 29368 26522 29420 26528
rect 30116 26518 30144 26930
rect 30104 26512 30156 26518
rect 30104 26454 30156 26460
rect 30748 26444 30800 26450
rect 30748 26386 30800 26392
rect 30196 26376 30248 26382
rect 30196 26318 30248 26324
rect 30208 26042 30236 26318
rect 30196 26036 30248 26042
rect 30196 25978 30248 25984
rect 30380 25968 30432 25974
rect 30380 25910 30432 25916
rect 29608 25596 29916 25605
rect 29608 25594 29614 25596
rect 29670 25594 29694 25596
rect 29750 25594 29774 25596
rect 29830 25594 29854 25596
rect 29910 25594 29916 25596
rect 29670 25542 29672 25594
rect 29852 25542 29854 25594
rect 29608 25540 29614 25542
rect 29670 25540 29694 25542
rect 29750 25540 29774 25542
rect 29830 25540 29854 25542
rect 29910 25540 29916 25542
rect 29608 25531 29916 25540
rect 29184 25492 29236 25498
rect 29184 25434 29236 25440
rect 28540 25356 28592 25362
rect 28540 25298 28592 25304
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 27620 23860 27672 23866
rect 27620 23802 27672 23808
rect 26976 23316 27028 23322
rect 26976 23258 27028 23264
rect 25872 22976 25924 22982
rect 25872 22918 25924 22924
rect 25514 22876 25822 22885
rect 25514 22874 25520 22876
rect 25576 22874 25600 22876
rect 25656 22874 25680 22876
rect 25736 22874 25760 22876
rect 25816 22874 25822 22876
rect 25576 22822 25578 22874
rect 25758 22822 25760 22874
rect 25514 22820 25520 22822
rect 25576 22820 25600 22822
rect 25656 22820 25680 22822
rect 25736 22820 25760 22822
rect 25816 22820 25822 22822
rect 25514 22811 25822 22820
rect 25514 21788 25822 21797
rect 25514 21786 25520 21788
rect 25576 21786 25600 21788
rect 25656 21786 25680 21788
rect 25736 21786 25760 21788
rect 25816 21786 25822 21788
rect 25576 21734 25578 21786
rect 25758 21734 25760 21786
rect 25514 21732 25520 21734
rect 25576 21732 25600 21734
rect 25656 21732 25680 21734
rect 25736 21732 25760 21734
rect 25816 21732 25822 21734
rect 25514 21723 25822 21732
rect 25412 21140 25464 21146
rect 25412 21082 25464 21088
rect 24768 20936 24820 20942
rect 24768 20878 24820 20884
rect 17326 20700 17634 20709
rect 17326 20698 17332 20700
rect 17388 20698 17412 20700
rect 17468 20698 17492 20700
rect 17548 20698 17572 20700
rect 17628 20698 17634 20700
rect 17388 20646 17390 20698
rect 17570 20646 17572 20698
rect 17326 20644 17332 20646
rect 17388 20644 17412 20646
rect 17468 20644 17492 20646
rect 17548 20644 17572 20646
rect 17628 20644 17634 20646
rect 17326 20635 17634 20644
rect 21420 20156 21728 20165
rect 21420 20154 21426 20156
rect 21482 20154 21506 20156
rect 21562 20154 21586 20156
rect 21642 20154 21666 20156
rect 21722 20154 21728 20156
rect 21482 20102 21484 20154
rect 21664 20102 21666 20154
rect 21420 20100 21426 20102
rect 21482 20100 21506 20102
rect 21562 20100 21586 20102
rect 21642 20100 21666 20102
rect 21722 20100 21728 20102
rect 21420 20091 21728 20100
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 17326 19612 17634 19621
rect 17326 19610 17332 19612
rect 17388 19610 17412 19612
rect 17468 19610 17492 19612
rect 17548 19610 17572 19612
rect 17628 19610 17634 19612
rect 17388 19558 17390 19610
rect 17570 19558 17572 19610
rect 17326 19556 17332 19558
rect 17388 19556 17412 19558
rect 17468 19556 17492 19558
rect 17548 19556 17572 19558
rect 17628 19556 17634 19558
rect 17326 19547 17634 19556
rect 18064 18970 18092 19722
rect 21420 19068 21728 19077
rect 21420 19066 21426 19068
rect 21482 19066 21506 19068
rect 21562 19066 21586 19068
rect 21642 19066 21666 19068
rect 21722 19066 21728 19068
rect 21482 19014 21484 19066
rect 21664 19014 21666 19066
rect 21420 19012 21426 19014
rect 21482 19012 21506 19014
rect 21562 19012 21586 19014
rect 21642 19012 21666 19014
rect 21722 19012 21728 19014
rect 21420 19003 21728 19012
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 19432 18896 19484 18902
rect 19432 18838 19484 18844
rect 17326 18524 17634 18533
rect 17326 18522 17332 18524
rect 17388 18522 17412 18524
rect 17468 18522 17492 18524
rect 17548 18522 17572 18524
rect 17628 18522 17634 18524
rect 17388 18470 17390 18522
rect 17570 18470 17572 18522
rect 17326 18468 17332 18470
rect 17388 18468 17412 18470
rect 17468 18468 17492 18470
rect 17548 18468 17572 18470
rect 17628 18468 17634 18470
rect 17326 18459 17634 18468
rect 19064 17604 19116 17610
rect 19064 17546 19116 17552
rect 19156 17604 19208 17610
rect 19156 17546 19208 17552
rect 17326 17436 17634 17445
rect 17326 17434 17332 17436
rect 17388 17434 17412 17436
rect 17468 17434 17492 17436
rect 17548 17434 17572 17436
rect 17628 17434 17634 17436
rect 17388 17382 17390 17434
rect 17570 17382 17572 17434
rect 17326 17380 17332 17382
rect 17388 17380 17412 17382
rect 17468 17380 17492 17382
rect 17548 17380 17572 17382
rect 17628 17380 17634 17382
rect 17326 17371 17634 17380
rect 17326 16348 17634 16357
rect 17326 16346 17332 16348
rect 17388 16346 17412 16348
rect 17468 16346 17492 16348
rect 17548 16346 17572 16348
rect 17628 16346 17634 16348
rect 17388 16294 17390 16346
rect 17570 16294 17572 16346
rect 17326 16292 17332 16294
rect 17388 16292 17412 16294
rect 17468 16292 17492 16294
rect 17548 16292 17572 16294
rect 17628 16292 17634 16294
rect 17326 16283 17634 16292
rect 17326 15260 17634 15269
rect 17326 15258 17332 15260
rect 17388 15258 17412 15260
rect 17468 15258 17492 15260
rect 17548 15258 17572 15260
rect 17628 15258 17634 15260
rect 17388 15206 17390 15258
rect 17570 15206 17572 15258
rect 17326 15204 17332 15206
rect 17388 15204 17412 15206
rect 17468 15204 17492 15206
rect 17548 15204 17572 15206
rect 17628 15204 17634 15206
rect 17326 15195 17634 15204
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18524 14618 18552 15030
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18616 14618 18644 14758
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 17326 14172 17634 14181
rect 17326 14170 17332 14172
rect 17388 14170 17412 14172
rect 17468 14170 17492 14172
rect 17548 14170 17572 14172
rect 17628 14170 17634 14172
rect 17388 14118 17390 14170
rect 17570 14118 17572 14170
rect 17326 14116 17332 14118
rect 17388 14116 17412 14118
rect 17468 14116 17492 14118
rect 17548 14116 17572 14118
rect 17628 14116 17634 14118
rect 17326 14107 17634 14116
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 13232 13628 13540 13637
rect 13232 13626 13238 13628
rect 13294 13626 13318 13628
rect 13374 13626 13398 13628
rect 13454 13626 13478 13628
rect 13534 13626 13540 13628
rect 13294 13574 13296 13626
rect 13476 13574 13478 13626
rect 13232 13572 13238 13574
rect 13294 13572 13318 13574
rect 13374 13572 13398 13574
rect 13454 13572 13478 13574
rect 13534 13572 13540 13574
rect 13232 13563 13540 13572
rect 13648 13190 13676 13806
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13232 12540 13540 12549
rect 13232 12538 13238 12540
rect 13294 12538 13318 12540
rect 13374 12538 13398 12540
rect 13454 12538 13478 12540
rect 13534 12538 13540 12540
rect 13294 12486 13296 12538
rect 13476 12486 13478 12538
rect 13232 12484 13238 12486
rect 13294 12484 13318 12486
rect 13374 12484 13398 12486
rect 13454 12484 13478 12486
rect 13534 12484 13540 12486
rect 13232 12475 13540 12484
rect 12716 11756 12768 11762
rect 12716 11698 12768 11704
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 12728 10606 12756 11698
rect 13232 11452 13540 11461
rect 13232 11450 13238 11452
rect 13294 11450 13318 11452
rect 13374 11450 13398 11452
rect 13454 11450 13478 11452
rect 13534 11450 13540 11452
rect 13294 11398 13296 11450
rect 13476 11398 13478 11450
rect 13232 11396 13238 11398
rect 13294 11396 13318 11398
rect 13374 11396 13398 11398
rect 13454 11396 13478 11398
rect 13534 11396 13540 11398
rect 13232 11387 13540 11396
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 12716 10600 12768 10606
rect 12716 10542 12768 10548
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9138 8732 9446 8741
rect 9138 8730 9144 8732
rect 9200 8730 9224 8732
rect 9280 8730 9304 8732
rect 9360 8730 9384 8732
rect 9440 8730 9446 8732
rect 9200 8678 9202 8730
rect 9382 8678 9384 8730
rect 9138 8676 9144 8678
rect 9200 8676 9224 8678
rect 9280 8676 9304 8678
rect 9360 8676 9384 8678
rect 9440 8676 9446 8678
rect 9138 8667 9446 8676
rect 9138 7644 9446 7653
rect 9138 7642 9144 7644
rect 9200 7642 9224 7644
rect 9280 7642 9304 7644
rect 9360 7642 9384 7644
rect 9440 7642 9446 7644
rect 9200 7590 9202 7642
rect 9382 7590 9384 7642
rect 9138 7588 9144 7590
rect 9200 7588 9224 7590
rect 9280 7588 9304 7590
rect 9360 7588 9384 7590
rect 9440 7588 9446 7590
rect 9138 7579 9446 7588
rect 9600 6914 9628 10542
rect 13232 10364 13540 10373
rect 13232 10362 13238 10364
rect 13294 10362 13318 10364
rect 13374 10362 13398 10364
rect 13454 10362 13478 10364
rect 13534 10362 13540 10364
rect 13294 10310 13296 10362
rect 13476 10310 13478 10362
rect 13232 10308 13238 10310
rect 13294 10308 13318 10310
rect 13374 10308 13398 10310
rect 13454 10308 13478 10310
rect 13534 10308 13540 10310
rect 13232 10299 13540 10308
rect 13232 9276 13540 9285
rect 13232 9274 13238 9276
rect 13294 9274 13318 9276
rect 13374 9274 13398 9276
rect 13454 9274 13478 9276
rect 13534 9274 13540 9276
rect 13294 9222 13296 9274
rect 13476 9222 13478 9274
rect 13232 9220 13238 9222
rect 13294 9220 13318 9222
rect 13374 9220 13398 9222
rect 13454 9220 13478 9222
rect 13534 9220 13540 9222
rect 13232 9211 13540 9220
rect 13232 8188 13540 8197
rect 13232 8186 13238 8188
rect 13294 8186 13318 8188
rect 13374 8186 13398 8188
rect 13454 8186 13478 8188
rect 13534 8186 13540 8188
rect 13294 8134 13296 8186
rect 13476 8134 13478 8186
rect 13232 8132 13238 8134
rect 13294 8132 13318 8134
rect 13374 8132 13398 8134
rect 13454 8132 13478 8134
rect 13534 8132 13540 8134
rect 13232 8123 13540 8132
rect 13232 7100 13540 7109
rect 13232 7098 13238 7100
rect 13294 7098 13318 7100
rect 13374 7098 13398 7100
rect 13454 7098 13478 7100
rect 13534 7098 13540 7100
rect 13294 7046 13296 7098
rect 13476 7046 13478 7098
rect 13232 7044 13238 7046
rect 13294 7044 13318 7046
rect 13374 7044 13398 7046
rect 13454 7044 13478 7046
rect 13534 7044 13540 7046
rect 13232 7035 13540 7044
rect 9508 6886 9628 6914
rect 9138 6556 9446 6565
rect 9138 6554 9144 6556
rect 9200 6554 9224 6556
rect 9280 6554 9304 6556
rect 9360 6554 9384 6556
rect 9440 6554 9446 6556
rect 9200 6502 9202 6554
rect 9382 6502 9384 6554
rect 9138 6500 9144 6502
rect 9200 6500 9224 6502
rect 9280 6500 9304 6502
rect 9360 6500 9384 6502
rect 9440 6500 9446 6502
rect 9138 6491 9446 6500
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9048 5166 9076 5510
rect 9138 5468 9446 5477
rect 9138 5466 9144 5468
rect 9200 5466 9224 5468
rect 9280 5466 9304 5468
rect 9360 5466 9384 5468
rect 9440 5466 9446 5468
rect 9200 5414 9202 5466
rect 9382 5414 9384 5466
rect 9138 5412 9144 5414
rect 9200 5412 9224 5414
rect 9280 5412 9304 5414
rect 9360 5412 9384 5414
rect 9440 5412 9446 5414
rect 9138 5403 9446 5412
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9508 4826 9536 6886
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9138 4380 9446 4389
rect 9138 4378 9144 4380
rect 9200 4378 9224 4380
rect 9280 4378 9304 4380
rect 9360 4378 9384 4380
rect 9440 4378 9446 4380
rect 9200 4326 9202 4378
rect 9382 4326 9384 4378
rect 9138 4324 9144 4326
rect 9200 4324 9224 4326
rect 9280 4324 9304 4326
rect 9360 4324 9384 4326
rect 9440 4324 9446 4326
rect 9138 4315 9446 4324
rect 9508 4282 9536 4762
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9508 3602 9536 4218
rect 9600 4146 9628 4422
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9138 3292 9446 3301
rect 9138 3290 9144 3292
rect 9200 3290 9224 3292
rect 9280 3290 9304 3292
rect 9360 3290 9384 3292
rect 9440 3290 9446 3292
rect 9200 3238 9202 3290
rect 9382 3238 9384 3290
rect 9138 3236 9144 3238
rect 9200 3236 9224 3238
rect 9280 3236 9304 3238
rect 9360 3236 9384 3238
rect 9440 3236 9446 3238
rect 9138 3227 9446 3236
rect 8772 3058 8892 3074
rect 9508 3058 9536 3538
rect 8760 3052 8892 3058
rect 8812 3046 8892 3052
rect 9496 3052 9548 3058
rect 8760 2994 8812 3000
rect 9496 2994 9548 3000
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 8116 2440 8168 2446
rect 9140 2394 9168 2790
rect 9784 2446 9812 5170
rect 9876 5030 9904 6122
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 10060 5370 10088 5646
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 3534 9904 4966
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10244 3466 10272 6054
rect 10428 5642 10456 6054
rect 13232 6012 13540 6021
rect 13232 6010 13238 6012
rect 13294 6010 13318 6012
rect 13374 6010 13398 6012
rect 13454 6010 13478 6012
rect 13534 6010 13540 6012
rect 13294 5958 13296 6010
rect 13476 5958 13478 6010
rect 13232 5956 13238 5958
rect 13294 5956 13318 5958
rect 13374 5956 13398 5958
rect 13454 5956 13478 5958
rect 13534 5956 13540 5958
rect 13232 5947 13540 5956
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10520 4826 10548 5102
rect 10704 4826 10732 5646
rect 11716 5370 11744 5782
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10796 4282 10824 5102
rect 12084 4826 12112 5102
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12360 4690 12388 5306
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 10784 4276 10836 4282
rect 10784 4218 10836 4224
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11348 3466 11376 3878
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 11440 3194 11468 4558
rect 11532 3738 11560 4626
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 9968 2514 9996 2994
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 8116 2382 8168 2388
rect 9048 2366 9168 2394
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9048 1578 9076 2366
rect 9138 2204 9446 2213
rect 9138 2202 9144 2204
rect 9200 2202 9224 2204
rect 9280 2202 9304 2204
rect 9360 2202 9384 2204
rect 9440 2202 9446 2204
rect 9200 2150 9202 2202
rect 9382 2150 9384 2202
rect 9138 2148 9144 2150
rect 9200 2148 9224 2150
rect 9280 2148 9304 2150
rect 9360 2148 9384 2150
rect 9440 2148 9446 2150
rect 9138 2139 9446 2148
rect 9048 1550 9168 1578
rect 9140 800 9168 1550
rect 10520 800 10548 2926
rect 11624 2514 11652 3334
rect 12452 2650 12480 5102
rect 12544 4282 12572 5510
rect 13648 5302 13676 13126
rect 17326 13084 17634 13093
rect 17326 13082 17332 13084
rect 17388 13082 17412 13084
rect 17468 13082 17492 13084
rect 17548 13082 17572 13084
rect 17628 13082 17634 13084
rect 17388 13030 17390 13082
rect 17570 13030 17572 13082
rect 17326 13028 17332 13030
rect 17388 13028 17412 13030
rect 17468 13028 17492 13030
rect 17548 13028 17572 13030
rect 17628 13028 17634 13030
rect 17326 13019 17634 13028
rect 17326 11996 17634 12005
rect 17326 11994 17332 11996
rect 17388 11994 17412 11996
rect 17468 11994 17492 11996
rect 17548 11994 17572 11996
rect 17628 11994 17634 11996
rect 17388 11942 17390 11994
rect 17570 11942 17572 11994
rect 17326 11940 17332 11942
rect 17388 11940 17412 11942
rect 17468 11940 17492 11942
rect 17548 11940 17572 11942
rect 17628 11940 17634 11942
rect 17326 11931 17634 11940
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 10130 15516 11494
rect 17326 10908 17634 10917
rect 17326 10906 17332 10908
rect 17388 10906 17412 10908
rect 17468 10906 17492 10908
rect 17548 10906 17572 10908
rect 17628 10906 17634 10908
rect 17388 10854 17390 10906
rect 17570 10854 17572 10906
rect 17326 10852 17332 10854
rect 17388 10852 17412 10854
rect 17468 10852 17492 10854
rect 17548 10852 17572 10854
rect 17628 10852 17634 10854
rect 17326 10843 17634 10852
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13740 5234 13768 5510
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13232 4924 13540 4933
rect 13232 4922 13238 4924
rect 13294 4922 13318 4924
rect 13374 4922 13398 4924
rect 13454 4922 13478 4924
rect 13534 4922 13540 4924
rect 13294 4870 13296 4922
rect 13476 4870 13478 4922
rect 13232 4868 13238 4870
rect 13294 4868 13318 4870
rect 13374 4868 13398 4870
rect 13454 4868 13478 4870
rect 13534 4868 13540 4870
rect 13232 4859 13540 4868
rect 13740 4826 13768 5170
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 13004 4146 13032 4422
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12624 4072 12676 4078
rect 12624 4014 12676 4020
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 11612 2508 11664 2514
rect 11612 2450 11664 2456
rect 12544 2446 12572 2926
rect 12636 2446 12664 4014
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3194 12940 3334
rect 13004 3194 13032 3470
rect 13096 3194 13124 4014
rect 13648 4010 13676 4422
rect 13832 4282 13860 4558
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13232 3836 13540 3845
rect 13232 3834 13238 3836
rect 13294 3834 13318 3836
rect 13374 3834 13398 3836
rect 13454 3834 13478 3836
rect 13534 3834 13540 3836
rect 13294 3782 13296 3834
rect 13476 3782 13478 3834
rect 13232 3780 13238 3782
rect 13294 3780 13318 3782
rect 13374 3780 13398 3782
rect 13454 3780 13478 3782
rect 13534 3780 13540 3782
rect 13232 3771 13540 3780
rect 13648 3602 13676 3946
rect 13924 3738 13952 9318
rect 15212 5914 15240 9454
rect 16960 7410 16988 9862
rect 17326 9820 17634 9829
rect 17326 9818 17332 9820
rect 17388 9818 17412 9820
rect 17468 9818 17492 9820
rect 17548 9818 17572 9820
rect 17628 9818 17634 9820
rect 17388 9766 17390 9818
rect 17570 9766 17572 9818
rect 17326 9764 17332 9766
rect 17388 9764 17412 9766
rect 17468 9764 17492 9766
rect 17548 9764 17572 9766
rect 17628 9764 17634 9766
rect 17326 9755 17634 9764
rect 18892 9518 18920 14486
rect 18880 9512 18932 9518
rect 18880 9454 18932 9460
rect 17326 8732 17634 8741
rect 17326 8730 17332 8732
rect 17388 8730 17412 8732
rect 17468 8730 17492 8732
rect 17548 8730 17572 8732
rect 17628 8730 17634 8732
rect 17388 8678 17390 8730
rect 17570 8678 17572 8730
rect 17326 8676 17332 8678
rect 17388 8676 17412 8678
rect 17468 8676 17492 8678
rect 17548 8676 17572 8678
rect 17628 8676 17634 8678
rect 17326 8667 17634 8676
rect 17326 7644 17634 7653
rect 17326 7642 17332 7644
rect 17388 7642 17412 7644
rect 17468 7642 17492 7644
rect 17548 7642 17572 7644
rect 17628 7642 17634 7644
rect 17388 7590 17390 7642
rect 17570 7590 17572 7642
rect 17326 7588 17332 7590
rect 17388 7588 17412 7590
rect 17468 7588 17492 7590
rect 17548 7588 17572 7590
rect 17628 7588 17634 7590
rect 17326 7579 17634 7588
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14108 3738 14136 4014
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 12900 3188 12952 3194
rect 12900 3130 12952 3136
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13232 2748 13540 2757
rect 13232 2746 13238 2748
rect 13294 2746 13318 2748
rect 13374 2746 13398 2748
rect 13454 2746 13478 2748
rect 13534 2746 13540 2748
rect 13294 2694 13296 2746
rect 13476 2694 13478 2746
rect 13232 2692 13238 2694
rect 13294 2692 13318 2694
rect 13374 2692 13398 2694
rect 13454 2692 13478 2694
rect 13534 2692 13540 2694
rect 13232 2683 13540 2692
rect 14384 2650 14412 4694
rect 15948 4622 15976 5238
rect 16776 5234 16804 7142
rect 17326 6556 17634 6565
rect 17326 6554 17332 6556
rect 17388 6554 17412 6556
rect 17468 6554 17492 6556
rect 17548 6554 17572 6556
rect 17628 6554 17634 6556
rect 17388 6502 17390 6554
rect 17570 6502 17572 6554
rect 17326 6500 17332 6502
rect 17388 6500 17412 6502
rect 17468 6500 17492 6502
rect 17548 6500 17572 6502
rect 17628 6500 17634 6502
rect 17326 6491 17634 6500
rect 17326 5468 17634 5477
rect 17326 5466 17332 5468
rect 17388 5466 17412 5468
rect 17468 5466 17492 5468
rect 17548 5466 17572 5468
rect 17628 5466 17634 5468
rect 17388 5414 17390 5466
rect 17570 5414 17572 5466
rect 17326 5412 17332 5414
rect 17388 5412 17412 5414
rect 17468 5412 17492 5414
rect 17548 5412 17572 5414
rect 17628 5412 17634 5414
rect 17326 5403 17634 5412
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 14476 3058 14504 4422
rect 15396 4146 15424 4422
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14660 2514 14688 3878
rect 15488 3398 15516 4422
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 16040 3194 16068 4014
rect 16592 3602 16620 5102
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 16672 4616 16724 4622
rect 16672 4558 16724 4564
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16684 3194 16712 4558
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16776 4146 16804 4422
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16868 3466 16896 4422
rect 17326 4380 17634 4389
rect 17326 4378 17332 4380
rect 17388 4378 17412 4380
rect 17468 4378 17492 4380
rect 17548 4378 17572 4380
rect 17628 4378 17634 4380
rect 17388 4326 17390 4378
rect 17570 4326 17572 4378
rect 17326 4324 17332 4326
rect 17388 4324 17412 4326
rect 17468 4324 17492 4326
rect 17548 4324 17572 4326
rect 17628 4324 17634 4326
rect 17326 4315 17634 4324
rect 18708 4146 18736 4694
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 14832 2984 14884 2990
rect 14832 2926 14884 2932
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 11900 800 11928 2382
rect 13280 800 13308 2450
rect 14844 1578 14872 2926
rect 16960 2514 16988 3334
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 16948 2508 17000 2514
rect 16948 2450 17000 2456
rect 14660 1550 14872 1578
rect 14660 800 14688 1550
rect 16040 800 16068 2450
rect 17052 2446 17080 4014
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 17326 3292 17634 3301
rect 17326 3290 17332 3292
rect 17388 3290 17412 3292
rect 17468 3290 17492 3292
rect 17548 3290 17572 3292
rect 17628 3290 17634 3292
rect 17388 3238 17390 3290
rect 17570 3238 17572 3290
rect 17326 3236 17332 3238
rect 17388 3236 17412 3238
rect 17468 3236 17492 3238
rect 17548 3236 17572 3238
rect 17628 3236 17634 3238
rect 17326 3227 17634 3236
rect 18156 3194 18184 3878
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17684 2984 17736 2990
rect 17684 2926 17736 2932
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 17328 2650 17356 2926
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17696 2446 17724 2926
rect 17880 2514 18000 2530
rect 17880 2508 18012 2514
rect 17880 2502 17960 2508
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17326 2204 17634 2213
rect 17326 2202 17332 2204
rect 17388 2202 17412 2204
rect 17468 2202 17492 2204
rect 17548 2202 17572 2204
rect 17628 2202 17634 2204
rect 17388 2150 17390 2202
rect 17570 2150 17572 2202
rect 17326 2148 17332 2150
rect 17388 2148 17412 2150
rect 17468 2148 17492 2150
rect 17548 2148 17572 2150
rect 17628 2148 17634 2150
rect 17326 2139 17634 2148
rect 17420 870 17540 898
rect 17420 800 17448 870
rect 6472 734 6776 762
rect 7746 0 7802 800
rect 9126 0 9182 800
rect 10506 0 10562 800
rect 11886 0 11942 800
rect 13266 0 13322 800
rect 14646 0 14702 800
rect 16026 0 16082 800
rect 17406 0 17462 800
rect 17512 762 17540 870
rect 17880 762 17908 2502
rect 17960 2450 18012 2456
rect 18800 800 18828 2926
rect 19076 2650 19104 17546
rect 19168 14618 19196 17546
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19352 11762 19380 14010
rect 19444 13326 19472 18838
rect 21420 17980 21728 17989
rect 21420 17978 21426 17980
rect 21482 17978 21506 17980
rect 21562 17978 21586 17980
rect 21642 17978 21666 17980
rect 21722 17978 21728 17980
rect 21482 17926 21484 17978
rect 21664 17926 21666 17978
rect 21420 17924 21426 17926
rect 21482 17924 21506 17926
rect 21562 17924 21586 17926
rect 21642 17924 21666 17926
rect 21722 17924 21728 17926
rect 21420 17915 21728 17924
rect 24780 17882 24808 20878
rect 25514 20700 25822 20709
rect 25514 20698 25520 20700
rect 25576 20698 25600 20700
rect 25656 20698 25680 20700
rect 25736 20698 25760 20700
rect 25816 20698 25822 20700
rect 25576 20646 25578 20698
rect 25758 20646 25760 20698
rect 25514 20644 25520 20646
rect 25576 20644 25600 20646
rect 25656 20644 25680 20646
rect 25736 20644 25760 20646
rect 25816 20644 25822 20646
rect 25514 20635 25822 20644
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25424 19378 25452 19654
rect 25514 19612 25822 19621
rect 25514 19610 25520 19612
rect 25576 19610 25600 19612
rect 25656 19610 25680 19612
rect 25736 19610 25760 19612
rect 25816 19610 25822 19612
rect 25576 19558 25578 19610
rect 25758 19558 25760 19610
rect 25514 19556 25520 19558
rect 25576 19556 25600 19558
rect 25656 19556 25680 19558
rect 25736 19556 25760 19558
rect 25816 19556 25822 19558
rect 25514 19547 25822 19556
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25516 18714 25544 19382
rect 25424 18686 25544 18714
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 21420 16892 21728 16901
rect 21420 16890 21426 16892
rect 21482 16890 21506 16892
rect 21562 16890 21586 16892
rect 21642 16890 21666 16892
rect 21722 16890 21728 16892
rect 21482 16838 21484 16890
rect 21664 16838 21666 16890
rect 21420 16836 21426 16838
rect 21482 16836 21506 16838
rect 21562 16836 21586 16838
rect 21642 16836 21666 16838
rect 21722 16836 21728 16838
rect 21420 16827 21728 16836
rect 21836 16794 21864 17818
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19536 14822 19564 16594
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20732 15026 20760 16526
rect 21420 15804 21728 15813
rect 21420 15802 21426 15804
rect 21482 15802 21506 15804
rect 21562 15802 21586 15804
rect 21642 15802 21666 15804
rect 21722 15802 21728 15804
rect 21482 15750 21484 15802
rect 21664 15750 21666 15802
rect 21420 15748 21426 15750
rect 21482 15748 21506 15750
rect 21562 15748 21586 15750
rect 21642 15748 21666 15750
rect 21722 15748 21728 15750
rect 21420 15739 21728 15748
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 19524 14816 19576 14822
rect 19524 14758 19576 14764
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19812 14074 19840 14758
rect 21420 14716 21728 14725
rect 21420 14714 21426 14716
rect 21482 14714 21506 14716
rect 21562 14714 21586 14716
rect 21642 14714 21666 14716
rect 21722 14714 21728 14716
rect 21482 14662 21484 14714
rect 21664 14662 21666 14714
rect 21420 14660 21426 14662
rect 21482 14660 21506 14662
rect 21562 14660 21586 14662
rect 21642 14660 21666 14662
rect 21722 14660 21728 14662
rect 21420 14651 21728 14660
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 21008 13938 21036 14214
rect 22020 13938 22048 17614
rect 24964 16522 24992 17614
rect 24952 16516 25004 16522
rect 24952 16458 25004 16464
rect 25424 15706 25452 18686
rect 25514 18524 25822 18533
rect 25514 18522 25520 18524
rect 25576 18522 25600 18524
rect 25656 18522 25680 18524
rect 25736 18522 25760 18524
rect 25816 18522 25822 18524
rect 25576 18470 25578 18522
rect 25758 18470 25760 18522
rect 25514 18468 25520 18470
rect 25576 18468 25600 18470
rect 25656 18468 25680 18470
rect 25736 18468 25760 18470
rect 25816 18468 25822 18470
rect 25514 18459 25822 18468
rect 25884 17610 25912 22918
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 26804 19514 26832 22510
rect 26988 19718 27016 23258
rect 28736 22778 28764 25230
rect 29608 24508 29916 24517
rect 29608 24506 29614 24508
rect 29670 24506 29694 24508
rect 29750 24506 29774 24508
rect 29830 24506 29854 24508
rect 29910 24506 29916 24508
rect 29670 24454 29672 24506
rect 29852 24454 29854 24506
rect 29608 24452 29614 24454
rect 29670 24452 29694 24454
rect 29750 24452 29774 24454
rect 29830 24452 29854 24454
rect 29910 24452 29916 24454
rect 29608 24443 29916 24452
rect 29608 23420 29916 23429
rect 29608 23418 29614 23420
rect 29670 23418 29694 23420
rect 29750 23418 29774 23420
rect 29830 23418 29854 23420
rect 29910 23418 29916 23420
rect 29670 23366 29672 23418
rect 29852 23366 29854 23418
rect 29608 23364 29614 23366
rect 29670 23364 29694 23366
rect 29750 23364 29774 23366
rect 29830 23364 29854 23366
rect 29910 23364 29916 23366
rect 29608 23355 29916 23364
rect 28724 22772 28776 22778
rect 28724 22714 28776 22720
rect 29608 22332 29916 22341
rect 29608 22330 29614 22332
rect 29670 22330 29694 22332
rect 29750 22330 29774 22332
rect 29830 22330 29854 22332
rect 29910 22330 29916 22332
rect 29670 22278 29672 22330
rect 29852 22278 29854 22330
rect 29608 22276 29614 22278
rect 29670 22276 29694 22278
rect 29750 22276 29774 22278
rect 29830 22276 29854 22278
rect 29910 22276 29916 22278
rect 29608 22267 29916 22276
rect 29608 21244 29916 21253
rect 29608 21242 29614 21244
rect 29670 21242 29694 21244
rect 29750 21242 29774 21244
rect 29830 21242 29854 21244
rect 29910 21242 29916 21244
rect 29670 21190 29672 21242
rect 29852 21190 29854 21242
rect 29608 21188 29614 21190
rect 29670 21188 29694 21190
rect 29750 21188 29774 21190
rect 29830 21188 29854 21190
rect 29910 21188 29916 21190
rect 29608 21179 29916 21188
rect 29608 20156 29916 20165
rect 29608 20154 29614 20156
rect 29670 20154 29694 20156
rect 29750 20154 29774 20156
rect 29830 20154 29854 20156
rect 29910 20154 29916 20156
rect 29670 20102 29672 20154
rect 29852 20102 29854 20154
rect 29608 20100 29614 20102
rect 29670 20100 29694 20102
rect 29750 20100 29774 20102
rect 29830 20100 29854 20102
rect 29910 20100 29916 20102
rect 29608 20091 29916 20100
rect 28540 19848 28592 19854
rect 28540 19790 28592 19796
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26988 19514 27016 19654
rect 26792 19508 26844 19514
rect 26792 19450 26844 19456
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 25872 17604 25924 17610
rect 25872 17546 25924 17552
rect 25514 17436 25822 17445
rect 25514 17434 25520 17436
rect 25576 17434 25600 17436
rect 25656 17434 25680 17436
rect 25736 17434 25760 17436
rect 25816 17434 25822 17436
rect 25576 17382 25578 17434
rect 25758 17382 25760 17434
rect 25514 17380 25520 17382
rect 25576 17380 25600 17382
rect 25656 17380 25680 17382
rect 25736 17380 25760 17382
rect 25816 17380 25822 17382
rect 25514 17371 25822 17380
rect 25514 16348 25822 16357
rect 25514 16346 25520 16348
rect 25576 16346 25600 16348
rect 25656 16346 25680 16348
rect 25736 16346 25760 16348
rect 25816 16346 25822 16348
rect 25576 16294 25578 16346
rect 25758 16294 25760 16346
rect 25514 16292 25520 16294
rect 25576 16292 25600 16294
rect 25656 16292 25680 16294
rect 25736 16292 25760 16294
rect 25816 16292 25822 16294
rect 25514 16283 25822 16292
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 24952 15632 25004 15638
rect 24952 15574 25004 15580
rect 24584 15428 24636 15434
rect 24584 15370 24636 15376
rect 24596 15162 24624 15370
rect 24584 15156 24636 15162
rect 24584 15098 24636 15104
rect 23480 14884 23532 14890
rect 23480 14826 23532 14832
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21420 13628 21728 13637
rect 21420 13626 21426 13628
rect 21482 13626 21506 13628
rect 21562 13626 21586 13628
rect 21642 13626 21666 13628
rect 21722 13626 21728 13628
rect 21482 13574 21484 13626
rect 21664 13574 21666 13626
rect 21420 13572 21426 13574
rect 21482 13572 21506 13574
rect 21562 13572 21586 13574
rect 21642 13572 21666 13574
rect 21722 13572 21728 13574
rect 21420 13563 21728 13572
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19720 9178 19748 13262
rect 20352 13184 20404 13190
rect 20352 13126 20404 13132
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19996 9042 20024 11494
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 19352 2446 19380 4966
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19536 3738 19564 4014
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 20364 3534 20392 13126
rect 23492 12986 23520 14826
rect 24400 14544 24452 14550
rect 24400 14486 24452 14492
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 21420 12540 21728 12549
rect 21420 12538 21426 12540
rect 21482 12538 21506 12540
rect 21562 12538 21586 12540
rect 21642 12538 21666 12540
rect 21722 12538 21728 12540
rect 21482 12486 21484 12538
rect 21664 12486 21666 12538
rect 21420 12484 21426 12486
rect 21482 12484 21506 12486
rect 21562 12484 21586 12486
rect 21642 12484 21666 12486
rect 21722 12484 21728 12486
rect 21420 12475 21728 12484
rect 23676 12434 23704 12582
rect 23676 12406 23980 12434
rect 21420 11452 21728 11461
rect 21420 11450 21426 11452
rect 21482 11450 21506 11452
rect 21562 11450 21586 11452
rect 21642 11450 21666 11452
rect 21722 11450 21728 11452
rect 21482 11398 21484 11450
rect 21664 11398 21666 11450
rect 21420 11396 21426 11398
rect 21482 11396 21506 11398
rect 21562 11396 21586 11398
rect 21642 11396 21666 11398
rect 21722 11396 21728 11398
rect 21420 11387 21728 11396
rect 21420 10364 21728 10373
rect 21420 10362 21426 10364
rect 21482 10362 21506 10364
rect 21562 10362 21586 10364
rect 21642 10362 21666 10364
rect 21722 10362 21728 10364
rect 21482 10310 21484 10362
rect 21664 10310 21666 10362
rect 21420 10308 21426 10310
rect 21482 10308 21506 10310
rect 21562 10308 21586 10310
rect 21642 10308 21666 10310
rect 21722 10308 21728 10310
rect 21420 10299 21728 10308
rect 23664 9376 23716 9382
rect 23664 9318 23716 9324
rect 21420 9276 21728 9285
rect 21420 9274 21426 9276
rect 21482 9274 21506 9276
rect 21562 9274 21586 9276
rect 21642 9274 21666 9276
rect 21722 9274 21728 9276
rect 21482 9222 21484 9274
rect 21664 9222 21666 9274
rect 21420 9220 21426 9222
rect 21482 9220 21506 9222
rect 21562 9220 21586 9222
rect 21642 9220 21666 9222
rect 21722 9220 21728 9222
rect 21420 9211 21728 9220
rect 21420 8188 21728 8197
rect 21420 8186 21426 8188
rect 21482 8186 21506 8188
rect 21562 8186 21586 8188
rect 21642 8186 21666 8188
rect 21722 8186 21728 8188
rect 21482 8134 21484 8186
rect 21664 8134 21666 8186
rect 21420 8132 21426 8134
rect 21482 8132 21506 8134
rect 21562 8132 21586 8134
rect 21642 8132 21666 8134
rect 21722 8132 21728 8134
rect 21420 8123 21728 8132
rect 21420 7100 21728 7109
rect 21420 7098 21426 7100
rect 21482 7098 21506 7100
rect 21562 7098 21586 7100
rect 21642 7098 21666 7100
rect 21722 7098 21728 7100
rect 21482 7046 21484 7098
rect 21664 7046 21666 7098
rect 21420 7044 21426 7046
rect 21482 7044 21506 7046
rect 21562 7044 21586 7046
rect 21642 7044 21666 7046
rect 21722 7044 21728 7046
rect 21420 7035 21728 7044
rect 21420 6012 21728 6021
rect 21420 6010 21426 6012
rect 21482 6010 21506 6012
rect 21562 6010 21586 6012
rect 21642 6010 21666 6012
rect 21722 6010 21728 6012
rect 21482 5958 21484 6010
rect 21664 5958 21666 6010
rect 21420 5956 21426 5958
rect 21482 5956 21506 5958
rect 21562 5956 21586 5958
rect 21642 5956 21666 5958
rect 21722 5956 21728 5958
rect 21420 5947 21728 5956
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 21420 4924 21728 4933
rect 21420 4922 21426 4924
rect 21482 4922 21506 4924
rect 21562 4922 21586 4924
rect 21642 4922 21666 4924
rect 21722 4922 21728 4924
rect 21482 4870 21484 4922
rect 21664 4870 21666 4922
rect 21420 4868 21426 4870
rect 21482 4868 21506 4870
rect 21562 4868 21586 4870
rect 21642 4868 21666 4870
rect 21722 4868 21728 4870
rect 21420 4859 21728 4868
rect 23400 4690 23428 5238
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 22744 4480 22796 4486
rect 22744 4422 22796 4428
rect 21420 3836 21728 3845
rect 21420 3834 21426 3836
rect 21482 3834 21506 3836
rect 21562 3834 21586 3836
rect 21642 3834 21666 3836
rect 21722 3834 21728 3836
rect 21482 3782 21484 3834
rect 21664 3782 21666 3834
rect 21420 3780 21426 3782
rect 21482 3780 21506 3782
rect 21562 3780 21586 3782
rect 21642 3780 21666 3782
rect 21722 3780 21728 3782
rect 21420 3771 21728 3780
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 21916 3460 21968 3466
rect 21916 3402 21968 3408
rect 19708 3052 19760 3058
rect 19708 2994 19760 3000
rect 19720 2514 19748 2994
rect 21824 2916 21876 2922
rect 21824 2858 21876 2864
rect 21420 2748 21728 2757
rect 21420 2746 21426 2748
rect 21482 2746 21506 2748
rect 21562 2746 21586 2748
rect 21642 2746 21666 2748
rect 21722 2746 21728 2748
rect 21482 2694 21484 2746
rect 21664 2694 21666 2746
rect 21420 2692 21426 2694
rect 21482 2692 21506 2694
rect 21562 2692 21586 2694
rect 21642 2692 21666 2694
rect 21722 2692 21728 2694
rect 21420 2683 21728 2692
rect 19708 2508 19760 2514
rect 19708 2450 19760 2456
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 21836 1578 21864 2858
rect 21928 2446 21956 3402
rect 22204 3194 22232 3538
rect 22756 3534 22784 4422
rect 23204 4072 23256 4078
rect 23204 4014 23256 4020
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 21560 1550 21864 1578
rect 20352 1420 20404 1426
rect 20352 1362 20404 1368
rect 20364 1170 20392 1362
rect 20180 1142 20392 1170
rect 20180 800 20208 1142
rect 21560 800 21588 1550
rect 22020 1426 22048 2450
rect 22008 1420 22060 1426
rect 22008 1362 22060 1368
rect 22940 800 22968 3470
rect 23216 3194 23244 4014
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23308 2514 23336 3878
rect 23400 3738 23428 3878
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23388 3460 23440 3466
rect 23388 3402 23440 3408
rect 23296 2508 23348 2514
rect 23296 2450 23348 2456
rect 23400 2310 23428 3402
rect 23676 3058 23704 9318
rect 23952 4729 23980 12406
rect 24412 12306 24440 14486
rect 24400 12300 24452 12306
rect 24400 12242 24452 12248
rect 24964 9586 24992 15574
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 25044 12096 25096 12102
rect 25044 12038 25096 12044
rect 25056 9586 25084 12038
rect 24952 9580 25004 9586
rect 24952 9522 25004 9528
rect 25044 9580 25096 9586
rect 25044 9522 25096 9528
rect 24964 5534 24992 9522
rect 25240 6458 25268 15370
rect 25514 15260 25822 15269
rect 25514 15258 25520 15260
rect 25576 15258 25600 15260
rect 25656 15258 25680 15260
rect 25736 15258 25760 15260
rect 25816 15258 25822 15260
rect 25576 15206 25578 15258
rect 25758 15206 25760 15258
rect 25514 15204 25520 15206
rect 25576 15204 25600 15206
rect 25656 15204 25680 15206
rect 25736 15204 25760 15206
rect 25816 15204 25822 15206
rect 25514 15195 25822 15204
rect 25514 14172 25822 14181
rect 25514 14170 25520 14172
rect 25576 14170 25600 14172
rect 25656 14170 25680 14172
rect 25736 14170 25760 14172
rect 25816 14170 25822 14172
rect 25576 14118 25578 14170
rect 25758 14118 25760 14170
rect 25514 14116 25520 14118
rect 25576 14116 25600 14118
rect 25656 14116 25680 14118
rect 25736 14116 25760 14118
rect 25816 14116 25822 14118
rect 25514 14107 25822 14116
rect 25514 13084 25822 13093
rect 25514 13082 25520 13084
rect 25576 13082 25600 13084
rect 25656 13082 25680 13084
rect 25736 13082 25760 13084
rect 25816 13082 25822 13084
rect 25576 13030 25578 13082
rect 25758 13030 25760 13082
rect 25514 13028 25520 13030
rect 25576 13028 25600 13030
rect 25656 13028 25680 13030
rect 25736 13028 25760 13030
rect 25816 13028 25822 13030
rect 25514 13019 25822 13028
rect 25514 11996 25822 12005
rect 25514 11994 25520 11996
rect 25576 11994 25600 11996
rect 25656 11994 25680 11996
rect 25736 11994 25760 11996
rect 25816 11994 25822 11996
rect 25576 11942 25578 11994
rect 25758 11942 25760 11994
rect 25514 11940 25520 11942
rect 25576 11940 25600 11942
rect 25656 11940 25680 11942
rect 25736 11940 25760 11942
rect 25816 11940 25822 11942
rect 25514 11931 25822 11940
rect 25514 10908 25822 10917
rect 25514 10906 25520 10908
rect 25576 10906 25600 10908
rect 25656 10906 25680 10908
rect 25736 10906 25760 10908
rect 25816 10906 25822 10908
rect 25576 10854 25578 10906
rect 25758 10854 25760 10906
rect 25514 10852 25520 10854
rect 25576 10852 25600 10854
rect 25656 10852 25680 10854
rect 25736 10852 25760 10854
rect 25816 10852 25822 10854
rect 25514 10843 25822 10852
rect 25884 10266 25912 17546
rect 28552 16454 28580 19790
rect 29608 19068 29916 19077
rect 29608 19066 29614 19068
rect 29670 19066 29694 19068
rect 29750 19066 29774 19068
rect 29830 19066 29854 19068
rect 29910 19066 29916 19068
rect 29670 19014 29672 19066
rect 29852 19014 29854 19066
rect 29608 19012 29614 19014
rect 29670 19012 29694 19014
rect 29750 19012 29774 19014
rect 29830 19012 29854 19014
rect 29910 19012 29916 19014
rect 29608 19003 29916 19012
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 29608 17980 29916 17989
rect 29608 17978 29614 17980
rect 29670 17978 29694 17980
rect 29750 17978 29774 17980
rect 29830 17978 29854 17980
rect 29910 17978 29916 17980
rect 29670 17926 29672 17978
rect 29852 17926 29854 17978
rect 29608 17924 29614 17926
rect 29670 17924 29694 17926
rect 29750 17924 29774 17926
rect 29830 17924 29854 17926
rect 29910 17924 29916 17926
rect 29608 17915 29916 17924
rect 30300 17746 30328 18634
rect 30392 18426 30420 25910
rect 30564 25832 30616 25838
rect 30564 25774 30616 25780
rect 30576 24818 30604 25774
rect 30564 24812 30616 24818
rect 30564 24754 30616 24760
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 30668 23662 30696 24550
rect 30760 24410 30788 26386
rect 31680 26382 31708 27950
rect 31956 27538 31984 28018
rect 32140 28014 32168 29038
rect 32128 28008 32180 28014
rect 32128 27950 32180 27956
rect 32232 27606 32260 34326
rect 32310 34200 32366 34326
rect 33428 34326 33930 34354
rect 33048 31816 33100 31822
rect 33048 31758 33100 31764
rect 33060 30938 33088 31758
rect 33048 30932 33100 30938
rect 33048 30874 33100 30880
rect 32954 30288 33010 30297
rect 32954 30223 33010 30232
rect 32968 29238 32996 30223
rect 32956 29232 33008 29238
rect 32956 29174 33008 29180
rect 32220 27600 32272 27606
rect 32220 27542 32272 27548
rect 31944 27532 31996 27538
rect 31944 27474 31996 27480
rect 32220 27464 32272 27470
rect 32220 27406 32272 27412
rect 32232 27130 32260 27406
rect 32220 27124 32272 27130
rect 32220 27066 32272 27072
rect 33428 27062 33456 34326
rect 33874 34200 33930 34326
rect 33702 32668 34010 32677
rect 33702 32666 33708 32668
rect 33764 32666 33788 32668
rect 33844 32666 33868 32668
rect 33924 32666 33948 32668
rect 34004 32666 34010 32668
rect 33764 32614 33766 32666
rect 33946 32614 33948 32666
rect 33702 32612 33708 32614
rect 33764 32612 33788 32614
rect 33844 32612 33868 32614
rect 33924 32612 33948 32614
rect 34004 32612 34010 32614
rect 33702 32603 34010 32612
rect 33702 31580 34010 31589
rect 33702 31578 33708 31580
rect 33764 31578 33788 31580
rect 33844 31578 33868 31580
rect 33924 31578 33948 31580
rect 34004 31578 34010 31580
rect 33764 31526 33766 31578
rect 33946 31526 33948 31578
rect 33702 31524 33708 31526
rect 33764 31524 33788 31526
rect 33844 31524 33868 31526
rect 33924 31524 33948 31526
rect 34004 31524 34010 31526
rect 33702 31515 34010 31524
rect 33702 30492 34010 30501
rect 33702 30490 33708 30492
rect 33764 30490 33788 30492
rect 33844 30490 33868 30492
rect 33924 30490 33948 30492
rect 34004 30490 34010 30492
rect 33764 30438 33766 30490
rect 33946 30438 33948 30490
rect 33702 30436 33708 30438
rect 33764 30436 33788 30438
rect 33844 30436 33868 30438
rect 33924 30436 33948 30438
rect 34004 30436 34010 30438
rect 33702 30427 34010 30436
rect 33508 30048 33560 30054
rect 33508 29990 33560 29996
rect 33520 28694 33548 29990
rect 33702 29404 34010 29413
rect 33702 29402 33708 29404
rect 33764 29402 33788 29404
rect 33844 29402 33868 29404
rect 33924 29402 33948 29404
rect 34004 29402 34010 29404
rect 33764 29350 33766 29402
rect 33946 29350 33948 29402
rect 33702 29348 33708 29350
rect 33764 29348 33788 29350
rect 33844 29348 33868 29350
rect 33924 29348 33948 29350
rect 34004 29348 34010 29350
rect 33702 29339 34010 29348
rect 33508 28688 33560 28694
rect 33508 28630 33560 28636
rect 33702 28316 34010 28325
rect 33702 28314 33708 28316
rect 33764 28314 33788 28316
rect 33844 28314 33868 28316
rect 33924 28314 33948 28316
rect 34004 28314 34010 28316
rect 33764 28262 33766 28314
rect 33946 28262 33948 28314
rect 33702 28260 33708 28262
rect 33764 28260 33788 28262
rect 33844 28260 33868 28262
rect 33924 28260 33948 28262
rect 34004 28260 34010 28262
rect 33702 28251 34010 28260
rect 33702 27228 34010 27237
rect 33702 27226 33708 27228
rect 33764 27226 33788 27228
rect 33844 27226 33868 27228
rect 33924 27226 33948 27228
rect 34004 27226 34010 27228
rect 33764 27174 33766 27226
rect 33946 27174 33948 27226
rect 33702 27172 33708 27174
rect 33764 27172 33788 27174
rect 33844 27172 33868 27174
rect 33924 27172 33948 27174
rect 34004 27172 34010 27174
rect 33702 27163 34010 27172
rect 33416 27056 33468 27062
rect 33416 26998 33468 27004
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 30932 26376 30984 26382
rect 30932 26318 30984 26324
rect 31668 26376 31720 26382
rect 31668 26318 31720 26324
rect 30840 26240 30892 26246
rect 30944 26234 30972 26318
rect 30892 26206 30972 26234
rect 30840 26182 30892 26188
rect 30852 25770 30880 26182
rect 31208 25832 31260 25838
rect 31208 25774 31260 25780
rect 31300 25832 31352 25838
rect 31300 25774 31352 25780
rect 30840 25764 30892 25770
rect 30840 25706 30892 25712
rect 31220 25498 31248 25774
rect 31208 25492 31260 25498
rect 31208 25434 31260 25440
rect 31116 25220 31168 25226
rect 31116 25162 31168 25168
rect 31128 24857 31156 25162
rect 31312 24954 31340 25774
rect 31576 25288 31628 25294
rect 31576 25230 31628 25236
rect 31300 24948 31352 24954
rect 31300 24890 31352 24896
rect 31114 24848 31170 24857
rect 31114 24783 31170 24792
rect 30748 24404 30800 24410
rect 30748 24346 30800 24352
rect 30656 23656 30708 23662
rect 30656 23598 30708 23604
rect 30760 23322 30788 24346
rect 31312 24342 31340 24890
rect 31588 24886 31616 25230
rect 31576 24880 31628 24886
rect 31576 24822 31628 24828
rect 31300 24336 31352 24342
rect 31300 24278 31352 24284
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31300 24064 31352 24070
rect 31300 24006 31352 24012
rect 31312 23798 31340 24006
rect 31404 23866 31432 24142
rect 31392 23860 31444 23866
rect 31392 23802 31444 23808
rect 31300 23792 31352 23798
rect 31300 23734 31352 23740
rect 31300 23520 31352 23526
rect 31300 23462 31352 23468
rect 30748 23316 30800 23322
rect 30748 23258 30800 23264
rect 30760 21622 30788 23258
rect 31312 23186 31340 23462
rect 31404 23254 31432 23802
rect 31680 23730 31708 26318
rect 32220 26240 32272 26246
rect 32220 26182 32272 26188
rect 32232 25906 32260 26182
rect 32324 25974 32352 26930
rect 33324 26920 33376 26926
rect 33324 26862 33376 26868
rect 33336 26353 33364 26862
rect 33322 26344 33378 26353
rect 33322 26279 33378 26288
rect 33048 26240 33100 26246
rect 33048 26182 33100 26188
rect 33060 26042 33088 26182
rect 33702 26140 34010 26149
rect 33702 26138 33708 26140
rect 33764 26138 33788 26140
rect 33844 26138 33868 26140
rect 33924 26138 33948 26140
rect 34004 26138 34010 26140
rect 33764 26086 33766 26138
rect 33946 26086 33948 26138
rect 33702 26084 33708 26086
rect 33764 26084 33788 26086
rect 33844 26084 33868 26086
rect 33924 26084 33948 26086
rect 34004 26084 34010 26086
rect 33702 26075 34010 26084
rect 33048 26036 33100 26042
rect 33048 25978 33100 25984
rect 32312 25968 32364 25974
rect 32312 25910 32364 25916
rect 32220 25900 32272 25906
rect 32220 25842 32272 25848
rect 31760 25696 31812 25702
rect 31760 25638 31812 25644
rect 31944 25696 31996 25702
rect 31944 25638 31996 25644
rect 31772 25294 31800 25638
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 31956 24818 31984 25638
rect 33702 25052 34010 25061
rect 33702 25050 33708 25052
rect 33764 25050 33788 25052
rect 33844 25050 33868 25052
rect 33924 25050 33948 25052
rect 34004 25050 34010 25052
rect 33764 24998 33766 25050
rect 33946 24998 33948 25050
rect 33702 24996 33708 24998
rect 33764 24996 33788 24998
rect 33844 24996 33868 24998
rect 33924 24996 33948 24998
rect 34004 24996 34010 24998
rect 33702 24987 34010 24996
rect 31944 24812 31996 24818
rect 31944 24754 31996 24760
rect 31852 24744 31904 24750
rect 31852 24686 31904 24692
rect 31864 23866 31892 24686
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32036 24064 32088 24070
rect 32036 24006 32088 24012
rect 31852 23860 31904 23866
rect 31852 23802 31904 23808
rect 31668 23724 31720 23730
rect 31668 23666 31720 23672
rect 31392 23248 31444 23254
rect 31392 23190 31444 23196
rect 31300 23180 31352 23186
rect 31300 23122 31352 23128
rect 31300 22976 31352 22982
rect 31300 22918 31352 22924
rect 31392 22976 31444 22982
rect 31392 22918 31444 22924
rect 31312 21962 31340 22918
rect 31404 22098 31432 22918
rect 31484 22568 31536 22574
rect 31484 22510 31536 22516
rect 31496 22137 31524 22510
rect 31482 22128 31538 22137
rect 31392 22092 31444 22098
rect 31482 22063 31538 22072
rect 31392 22034 31444 22040
rect 31300 21956 31352 21962
rect 31300 21898 31352 21904
rect 30748 21616 30800 21622
rect 30748 21558 30800 21564
rect 30760 20058 30788 21558
rect 31404 21418 31432 22034
rect 31680 22030 31708 23666
rect 32048 23474 32076 24006
rect 32048 23446 32260 23474
rect 32232 23118 32260 23446
rect 32324 23186 32352 24142
rect 33324 24132 33376 24138
rect 33324 24074 33376 24080
rect 33048 23520 33100 23526
rect 33048 23462 33100 23468
rect 33336 23474 33364 24074
rect 33702 23964 34010 23973
rect 33702 23962 33708 23964
rect 33764 23962 33788 23964
rect 33844 23962 33868 23964
rect 33924 23962 33948 23964
rect 34004 23962 34010 23964
rect 33764 23910 33766 23962
rect 33946 23910 33948 23962
rect 33702 23908 33708 23910
rect 33764 23908 33788 23910
rect 33844 23908 33868 23910
rect 33924 23908 33948 23910
rect 34004 23908 34010 23910
rect 33702 23899 34010 23908
rect 33782 23488 33838 23497
rect 32312 23180 32364 23186
rect 32312 23122 32364 23128
rect 32220 23112 32272 23118
rect 32220 23054 32272 23060
rect 32036 22636 32088 22642
rect 32036 22578 32088 22584
rect 32048 22234 32076 22578
rect 33060 22234 33088 23462
rect 33336 23446 33782 23474
rect 33782 23423 33838 23432
rect 33702 22876 34010 22885
rect 33702 22874 33708 22876
rect 33764 22874 33788 22876
rect 33844 22874 33868 22876
rect 33924 22874 33948 22876
rect 34004 22874 34010 22876
rect 33764 22822 33766 22874
rect 33946 22822 33948 22874
rect 33702 22820 33708 22822
rect 33764 22820 33788 22822
rect 33844 22820 33868 22822
rect 33924 22820 33948 22822
rect 34004 22820 34010 22822
rect 33702 22811 34010 22820
rect 32036 22228 32088 22234
rect 32036 22170 32088 22176
rect 33048 22228 33100 22234
rect 33048 22170 33100 22176
rect 31668 22024 31720 22030
rect 31668 21966 31720 21972
rect 31392 21412 31444 21418
rect 31392 21354 31444 21360
rect 31208 21344 31260 21350
rect 31208 21286 31260 21292
rect 31300 21344 31352 21350
rect 31300 21286 31352 21292
rect 31220 20942 31248 21286
rect 31312 21010 31340 21286
rect 31300 21004 31352 21010
rect 31300 20946 31352 20952
rect 31680 20942 31708 21966
rect 33702 21788 34010 21797
rect 33702 21786 33708 21788
rect 33764 21786 33788 21788
rect 33844 21786 33868 21788
rect 33924 21786 33948 21788
rect 34004 21786 34010 21788
rect 33764 21734 33766 21786
rect 33946 21734 33948 21786
rect 33702 21732 33708 21734
rect 33764 21732 33788 21734
rect 33844 21732 33868 21734
rect 33924 21732 33948 21734
rect 34004 21732 34010 21734
rect 33702 21723 34010 21732
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 31944 21480 31996 21486
rect 31944 21422 31996 21428
rect 31956 21146 31984 21422
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31668 20936 31720 20942
rect 31668 20878 31720 20884
rect 31576 20800 31628 20806
rect 31576 20742 31628 20748
rect 31588 20398 31616 20742
rect 31576 20392 31628 20398
rect 31576 20334 31628 20340
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 30760 18426 30788 19994
rect 31300 19304 31352 19310
rect 31300 19246 31352 19252
rect 31312 18426 31340 19246
rect 31680 18834 31708 20878
rect 32324 20534 32352 21490
rect 33324 21480 33376 21486
rect 33324 21422 33376 21428
rect 33336 20913 33364 21422
rect 33322 20904 33378 20913
rect 33322 20839 33378 20848
rect 33702 20700 34010 20709
rect 33702 20698 33708 20700
rect 33764 20698 33788 20700
rect 33844 20698 33868 20700
rect 33924 20698 33948 20700
rect 34004 20698 34010 20700
rect 33764 20646 33766 20698
rect 33946 20646 33948 20698
rect 33702 20644 33708 20646
rect 33764 20644 33788 20646
rect 33844 20644 33868 20646
rect 33924 20644 33948 20646
rect 34004 20644 34010 20646
rect 33702 20635 34010 20644
rect 32312 20528 32364 20534
rect 32312 20470 32364 20476
rect 31852 20392 31904 20398
rect 31852 20334 31904 20340
rect 31864 19990 31892 20334
rect 31852 19984 31904 19990
rect 31852 19926 31904 19932
rect 32588 19780 32640 19786
rect 32588 19722 32640 19728
rect 32036 19712 32088 19718
rect 32036 19654 32088 19660
rect 31944 19168 31996 19174
rect 31944 19110 31996 19116
rect 31668 18828 31720 18834
rect 31668 18770 31720 18776
rect 31576 18624 31628 18630
rect 31576 18566 31628 18572
rect 30380 18420 30432 18426
rect 30380 18362 30432 18368
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 31024 18420 31076 18426
rect 31024 18362 31076 18368
rect 31300 18420 31352 18426
rect 31300 18362 31352 18368
rect 30288 17740 30340 17746
rect 30288 17682 30340 17688
rect 30392 17678 30420 18362
rect 31036 17746 31064 18362
rect 31312 17814 31340 18362
rect 31588 18290 31616 18566
rect 31956 18290 31984 19110
rect 32048 18698 32076 19654
rect 32600 19378 32628 19722
rect 33702 19612 34010 19621
rect 33702 19610 33708 19612
rect 33764 19610 33788 19612
rect 33844 19610 33868 19612
rect 33924 19610 33948 19612
rect 34004 19610 34010 19612
rect 33764 19558 33766 19610
rect 33946 19558 33948 19610
rect 33702 19556 33708 19558
rect 33764 19556 33788 19558
rect 33844 19556 33868 19558
rect 33924 19556 33948 19558
rect 34004 19556 34010 19558
rect 33702 19547 34010 19556
rect 33322 19408 33378 19417
rect 32588 19372 32640 19378
rect 33322 19343 33324 19352
rect 32588 19314 32640 19320
rect 33376 19343 33378 19352
rect 33324 19314 33376 19320
rect 32036 18692 32088 18698
rect 32036 18634 32088 18640
rect 33702 18524 34010 18533
rect 33702 18522 33708 18524
rect 33764 18522 33788 18524
rect 33844 18522 33868 18524
rect 33924 18522 33948 18524
rect 34004 18522 34010 18524
rect 33764 18470 33766 18522
rect 33946 18470 33948 18522
rect 33702 18468 33708 18470
rect 33764 18468 33788 18470
rect 33844 18468 33868 18470
rect 33924 18468 33948 18470
rect 34004 18468 34010 18470
rect 33702 18459 34010 18468
rect 31576 18284 31628 18290
rect 31576 18226 31628 18232
rect 31944 18284 31996 18290
rect 31944 18226 31996 18232
rect 32496 18216 32548 18222
rect 32496 18158 32548 18164
rect 31300 17808 31352 17814
rect 31300 17750 31352 17756
rect 31024 17740 31076 17746
rect 31024 17682 31076 17688
rect 32508 17678 32536 18158
rect 33322 18048 33378 18057
rect 33322 17983 33378 17992
rect 33336 17746 33364 17983
rect 33324 17740 33376 17746
rect 33324 17682 33376 17688
rect 30380 17672 30432 17678
rect 30380 17614 30432 17620
rect 32036 17672 32088 17678
rect 32036 17614 32088 17620
rect 32496 17672 32548 17678
rect 32496 17614 32548 17620
rect 29608 16892 29916 16901
rect 29608 16890 29614 16892
rect 29670 16890 29694 16892
rect 29750 16890 29774 16892
rect 29830 16890 29854 16892
rect 29910 16890 29916 16892
rect 29670 16838 29672 16890
rect 29852 16838 29854 16890
rect 29608 16836 29614 16838
rect 29670 16836 29694 16838
rect 29750 16836 29774 16838
rect 29830 16836 29854 16838
rect 29910 16836 29916 16838
rect 29608 16827 29916 16836
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 30392 16250 30420 17614
rect 30748 17536 30800 17542
rect 30748 17478 30800 17484
rect 31392 17536 31444 17542
rect 31392 17478 31444 17484
rect 30760 17270 30788 17478
rect 30748 17264 30800 17270
rect 30748 17206 30800 17212
rect 31404 16658 31432 17478
rect 32048 17338 32076 17614
rect 33702 17436 34010 17445
rect 33702 17434 33708 17436
rect 33764 17434 33788 17436
rect 33844 17434 33868 17436
rect 33924 17434 33948 17436
rect 34004 17434 34010 17436
rect 33764 17382 33766 17434
rect 33946 17382 33948 17434
rect 33702 17380 33708 17382
rect 33764 17380 33788 17382
rect 33844 17380 33868 17382
rect 33924 17380 33948 17382
rect 34004 17380 34010 17382
rect 33702 17371 34010 17380
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 31484 17128 31536 17134
rect 31484 17070 31536 17076
rect 31668 17128 31720 17134
rect 31668 17070 31720 17076
rect 31496 16697 31524 17070
rect 31482 16688 31538 16697
rect 31392 16652 31444 16658
rect 31482 16623 31538 16632
rect 31392 16594 31444 16600
rect 31392 16448 31444 16454
rect 31392 16390 31444 16396
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 29608 15804 29916 15813
rect 29608 15802 29614 15804
rect 29670 15802 29694 15804
rect 29750 15802 29774 15804
rect 29830 15802 29854 15804
rect 29910 15802 29916 15804
rect 29670 15750 29672 15802
rect 29852 15750 29854 15802
rect 29608 15748 29614 15750
rect 29670 15748 29694 15750
rect 29750 15748 29774 15750
rect 29830 15748 29854 15750
rect 29910 15748 29916 15750
rect 29608 15739 29916 15748
rect 30288 15564 30340 15570
rect 30288 15506 30340 15512
rect 30300 14890 30328 15506
rect 30392 14958 30420 16186
rect 31404 16114 31432 16390
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31680 15502 31708 17070
rect 31956 16794 31984 17138
rect 31944 16788 31996 16794
rect 31944 16730 31996 16736
rect 32220 16584 32272 16590
rect 32220 16526 32272 16532
rect 32232 16250 32260 16526
rect 33702 16348 34010 16357
rect 33702 16346 33708 16348
rect 33764 16346 33788 16348
rect 33844 16346 33868 16348
rect 33924 16346 33948 16348
rect 34004 16346 34010 16348
rect 33764 16294 33766 16346
rect 33946 16294 33948 16346
rect 33702 16292 33708 16294
rect 33764 16292 33788 16294
rect 33844 16292 33868 16294
rect 33924 16292 33948 16294
rect 34004 16292 34010 16294
rect 33702 16283 34010 16292
rect 32220 16244 32272 16250
rect 32220 16186 32272 16192
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31772 15502 31800 15846
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 31668 15496 31720 15502
rect 31668 15438 31720 15444
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 30852 15162 30880 15438
rect 31576 15360 31628 15366
rect 31576 15302 31628 15308
rect 30840 15156 30892 15162
rect 30840 15098 30892 15104
rect 31588 15026 31616 15302
rect 31576 15020 31628 15026
rect 31576 14962 31628 14968
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 29608 14716 29916 14725
rect 29608 14714 29614 14716
rect 29670 14714 29694 14716
rect 29750 14714 29774 14716
rect 29830 14714 29854 14716
rect 29910 14714 29916 14716
rect 29670 14662 29672 14714
rect 29852 14662 29854 14714
rect 29608 14660 29614 14662
rect 29670 14660 29694 14662
rect 29750 14660 29774 14662
rect 29830 14660 29854 14662
rect 29910 14660 29916 14662
rect 29608 14651 29916 14660
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26528 10266 26556 13874
rect 30024 13870 30052 14758
rect 30576 14074 30604 14894
rect 31300 14816 31352 14822
rect 31300 14758 31352 14764
rect 31116 14340 31168 14346
rect 31116 14282 31168 14288
rect 31024 14272 31076 14278
rect 31024 14214 31076 14220
rect 30564 14068 30616 14074
rect 30564 14010 30616 14016
rect 31036 13870 31064 14214
rect 31128 13977 31156 14282
rect 31114 13968 31170 13977
rect 31114 13903 31170 13912
rect 31208 13932 31260 13938
rect 31208 13874 31260 13880
rect 30012 13864 30064 13870
rect 30012 13806 30064 13812
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 31024 13864 31076 13870
rect 31024 13806 31076 13812
rect 29608 13628 29916 13637
rect 29608 13626 29614 13628
rect 29670 13626 29694 13628
rect 29750 13626 29774 13628
rect 29830 13626 29854 13628
rect 29910 13626 29916 13628
rect 29670 13574 29672 13626
rect 29852 13574 29854 13626
rect 29608 13572 29614 13574
rect 29670 13572 29694 13574
rect 29750 13572 29774 13574
rect 29830 13572 29854 13574
rect 29910 13572 29916 13574
rect 29608 13563 29916 13572
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 26516 10260 26568 10266
rect 26516 10202 26568 10208
rect 25514 9820 25822 9829
rect 25514 9818 25520 9820
rect 25576 9818 25600 9820
rect 25656 9818 25680 9820
rect 25736 9818 25760 9820
rect 25816 9818 25822 9820
rect 25576 9766 25578 9818
rect 25758 9766 25760 9818
rect 25514 9764 25520 9766
rect 25576 9764 25600 9766
rect 25656 9764 25680 9766
rect 25736 9764 25760 9766
rect 25816 9764 25822 9766
rect 25514 9755 25822 9764
rect 25514 8732 25822 8741
rect 25514 8730 25520 8732
rect 25576 8730 25600 8732
rect 25656 8730 25680 8732
rect 25736 8730 25760 8732
rect 25816 8730 25822 8732
rect 25576 8678 25578 8730
rect 25758 8678 25760 8730
rect 25514 8676 25520 8678
rect 25576 8676 25600 8678
rect 25656 8676 25680 8678
rect 25736 8676 25760 8678
rect 25816 8676 25822 8678
rect 25514 8667 25822 8676
rect 25514 7644 25822 7653
rect 25514 7642 25520 7644
rect 25576 7642 25600 7644
rect 25656 7642 25680 7644
rect 25736 7642 25760 7644
rect 25816 7642 25822 7644
rect 25576 7590 25578 7642
rect 25758 7590 25760 7642
rect 25514 7588 25520 7590
rect 25576 7588 25600 7590
rect 25656 7588 25680 7590
rect 25736 7588 25760 7590
rect 25816 7588 25822 7590
rect 25514 7579 25822 7588
rect 26240 6928 26292 6934
rect 26240 6870 26292 6876
rect 25514 6556 25822 6565
rect 25514 6554 25520 6556
rect 25576 6554 25600 6556
rect 25656 6554 25680 6556
rect 25736 6554 25760 6556
rect 25816 6554 25822 6556
rect 25576 6502 25578 6554
rect 25758 6502 25760 6554
rect 25514 6500 25520 6502
rect 25576 6500 25600 6502
rect 25656 6500 25680 6502
rect 25736 6500 25760 6502
rect 25816 6500 25822 6502
rect 25514 6491 25822 6500
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25240 5846 25268 6394
rect 26148 5908 26200 5914
rect 26148 5850 26200 5856
rect 25228 5840 25280 5846
rect 25228 5782 25280 5788
rect 24964 5506 25084 5534
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24032 5024 24084 5030
rect 24032 4966 24084 4972
rect 24044 4826 24072 4966
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 23938 4720 23994 4729
rect 23938 4655 23994 4664
rect 24216 4480 24268 4486
rect 24216 4422 24268 4428
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24136 3194 24164 3334
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 24228 2446 24256 4422
rect 24320 3738 24348 5170
rect 24584 5160 24636 5166
rect 24584 5102 24636 5108
rect 24596 4826 24624 5102
rect 24584 4820 24636 4826
rect 24584 4762 24636 4768
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 24860 4548 24912 4554
rect 24860 4490 24912 4496
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 24412 3738 24440 4082
rect 24596 3738 24624 4082
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 24584 3732 24636 3738
rect 24584 3674 24636 3680
rect 24320 3618 24348 3674
rect 24320 3590 24716 3618
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 24216 2440 24268 2446
rect 24216 2382 24268 2388
rect 23388 2304 23440 2310
rect 23388 2246 23440 2252
rect 23860 2106 23888 2382
rect 23848 2100 23900 2106
rect 23848 2042 23900 2048
rect 24504 1714 24532 3334
rect 24688 2446 24716 3590
rect 24780 3534 24808 4014
rect 24872 3738 24900 4490
rect 24964 4282 24992 4558
rect 24952 4276 25004 4282
rect 24952 4218 25004 4224
rect 24860 3732 24912 3738
rect 24860 3674 24912 3680
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25056 2666 25084 5506
rect 25240 5302 25268 5782
rect 25514 5468 25822 5477
rect 25514 5466 25520 5468
rect 25576 5466 25600 5468
rect 25656 5466 25680 5468
rect 25736 5466 25760 5468
rect 25816 5466 25822 5468
rect 25576 5414 25578 5466
rect 25758 5414 25760 5466
rect 25514 5412 25520 5414
rect 25576 5412 25600 5414
rect 25656 5412 25680 5414
rect 25736 5412 25760 5414
rect 25816 5412 25822 5414
rect 25514 5403 25822 5412
rect 26056 5364 26108 5370
rect 26056 5306 26108 5312
rect 25228 5296 25280 5302
rect 26068 5273 26096 5306
rect 25228 5238 25280 5244
rect 26054 5264 26110 5273
rect 26054 5199 26110 5208
rect 25412 4616 25464 4622
rect 25412 4558 25464 4564
rect 25424 3738 25452 4558
rect 26056 4480 26108 4486
rect 26056 4422 26108 4428
rect 25514 4380 25822 4389
rect 25514 4378 25520 4380
rect 25576 4378 25600 4380
rect 25656 4378 25680 4380
rect 25736 4378 25760 4380
rect 25816 4378 25822 4380
rect 25576 4326 25578 4378
rect 25758 4326 25760 4378
rect 25514 4324 25520 4326
rect 25576 4324 25600 4326
rect 25656 4324 25680 4326
rect 25736 4324 25760 4326
rect 25816 4324 25822 4326
rect 25514 4315 25822 4324
rect 25412 3732 25464 3738
rect 25412 3674 25464 3680
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 24964 2638 25084 2666
rect 24964 2582 24992 2638
rect 25332 2582 25360 3470
rect 25514 3292 25822 3301
rect 25514 3290 25520 3292
rect 25576 3290 25600 3292
rect 25656 3290 25680 3292
rect 25736 3290 25760 3292
rect 25816 3290 25822 3292
rect 25576 3238 25578 3290
rect 25758 3238 25760 3290
rect 25514 3236 25520 3238
rect 25576 3236 25600 3238
rect 25656 3236 25680 3238
rect 25736 3236 25760 3238
rect 25816 3236 25822 3238
rect 25514 3227 25822 3236
rect 24952 2576 25004 2582
rect 24952 2518 25004 2524
rect 25320 2576 25372 2582
rect 25320 2518 25372 2524
rect 26068 2446 26096 4422
rect 26160 4060 26188 5850
rect 26252 5234 26280 6870
rect 26528 5914 26556 10202
rect 26988 9722 27016 12786
rect 29608 12540 29916 12549
rect 29608 12538 29614 12540
rect 29670 12538 29694 12540
rect 29750 12538 29774 12540
rect 29830 12538 29854 12540
rect 29910 12538 29916 12540
rect 29670 12486 29672 12538
rect 29852 12486 29854 12538
rect 29608 12484 29614 12486
rect 29670 12484 29694 12486
rect 29750 12484 29774 12486
rect 29830 12484 29854 12486
rect 29910 12484 29916 12486
rect 29608 12475 29916 12484
rect 30576 12442 30604 13806
rect 31220 13326 31248 13874
rect 31312 13870 31340 14758
rect 31680 14482 31708 15438
rect 32324 15094 32352 16050
rect 33324 16040 33376 16046
rect 33324 15982 33376 15988
rect 33336 15473 33364 15982
rect 33322 15464 33378 15473
rect 33322 15399 33378 15408
rect 33048 15360 33100 15366
rect 33048 15302 33100 15308
rect 32312 15088 32364 15094
rect 32312 15030 32364 15036
rect 33060 15026 33088 15302
rect 33702 15260 34010 15269
rect 33702 15258 33708 15260
rect 33764 15258 33788 15260
rect 33844 15258 33868 15260
rect 33924 15258 33948 15260
rect 34004 15258 34010 15260
rect 33764 15206 33766 15258
rect 33946 15206 33948 15258
rect 33702 15204 33708 15206
rect 33764 15204 33788 15206
rect 33844 15204 33868 15206
rect 33924 15204 33948 15206
rect 34004 15204 34010 15206
rect 33702 15195 34010 15204
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 31760 14884 31812 14890
rect 31760 14826 31812 14832
rect 31668 14476 31720 14482
rect 31668 14418 31720 14424
rect 31576 14408 31628 14414
rect 31576 14350 31628 14356
rect 31588 14006 31616 14350
rect 31576 14000 31628 14006
rect 31576 13942 31628 13948
rect 31300 13864 31352 13870
rect 31300 13806 31352 13812
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 30840 13184 30892 13190
rect 30840 13126 30892 13132
rect 30852 12850 30880 13126
rect 30944 12850 30972 13262
rect 31220 12986 31248 13262
rect 31576 13184 31628 13190
rect 31576 13126 31628 13132
rect 31208 12980 31260 12986
rect 31208 12922 31260 12928
rect 31588 12850 31616 13126
rect 30840 12844 30892 12850
rect 30840 12786 30892 12792
rect 30932 12844 30984 12850
rect 30932 12786 30984 12792
rect 31576 12844 31628 12850
rect 31576 12786 31628 12792
rect 30564 12436 30616 12442
rect 30564 12378 30616 12384
rect 29608 11452 29916 11461
rect 29608 11450 29614 11452
rect 29670 11450 29694 11452
rect 29750 11450 29774 11452
rect 29830 11450 29854 11452
rect 29910 11450 29916 11452
rect 29670 11398 29672 11450
rect 29852 11398 29854 11450
rect 29608 11396 29614 11398
rect 29670 11396 29694 11398
rect 29750 11396 29774 11398
rect 29830 11396 29854 11398
rect 29910 11396 29916 11398
rect 29608 11387 29916 11396
rect 30576 11354 30604 12378
rect 30944 12374 30972 12786
rect 30932 12368 30984 12374
rect 30932 12310 30984 12316
rect 31300 12096 31352 12102
rect 31300 12038 31352 12044
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31312 11830 31340 12038
rect 31300 11824 31352 11830
rect 31300 11766 31352 11772
rect 30564 11348 30616 11354
rect 30564 11290 30616 11296
rect 30576 10674 30604 11290
rect 31404 11218 31432 12038
rect 31680 11762 31708 14418
rect 31772 14414 31800 14826
rect 31760 14408 31812 14414
rect 31760 14350 31812 14356
rect 33702 14172 34010 14181
rect 33702 14170 33708 14172
rect 33764 14170 33788 14172
rect 33844 14170 33868 14172
rect 33924 14170 33948 14172
rect 34004 14170 34010 14172
rect 33764 14118 33766 14170
rect 33946 14118 33948 14170
rect 33702 14116 33708 14118
rect 33764 14116 33788 14118
rect 33844 14116 33868 14118
rect 33924 14116 33948 14118
rect 34004 14116 34010 14118
rect 33702 14107 34010 14116
rect 31760 13728 31812 13734
rect 31760 13670 31812 13676
rect 31772 13326 31800 13670
rect 31760 13320 31812 13326
rect 31760 13262 31812 13268
rect 33702 13084 34010 13093
rect 33702 13082 33708 13084
rect 33764 13082 33788 13084
rect 33844 13082 33868 13084
rect 33924 13082 33948 13084
rect 34004 13082 34010 13084
rect 33764 13030 33766 13082
rect 33946 13030 33948 13082
rect 33702 13028 33708 13030
rect 33764 13028 33788 13030
rect 33844 13028 33868 13030
rect 33924 13028 33948 13030
rect 34004 13028 34010 13030
rect 33702 13019 34010 13028
rect 32496 12776 32548 12782
rect 32496 12718 32548 12724
rect 32508 12238 32536 12718
rect 33322 12608 33378 12617
rect 33322 12543 33378 12552
rect 33336 12306 33364 12543
rect 33324 12300 33376 12306
rect 33324 12242 33376 12248
rect 32036 12232 32088 12238
rect 32036 12174 32088 12180
rect 32496 12232 32548 12238
rect 32496 12174 32548 12180
rect 32048 11898 32076 12174
rect 33702 11996 34010 12005
rect 33702 11994 33708 11996
rect 33764 11994 33788 11996
rect 33844 11994 33868 11996
rect 33924 11994 33948 11996
rect 34004 11994 34010 11996
rect 33764 11942 33766 11994
rect 33946 11942 33948 11994
rect 33702 11940 33708 11942
rect 33764 11940 33788 11942
rect 33844 11940 33868 11942
rect 33924 11940 33948 11942
rect 34004 11940 34010 11942
rect 33702 11931 34010 11940
rect 32036 11892 32088 11898
rect 32036 11834 32088 11840
rect 31668 11756 31720 11762
rect 31668 11698 31720 11704
rect 31944 11756 31996 11762
rect 31944 11698 31996 11704
rect 31484 11688 31536 11694
rect 31484 11630 31536 11636
rect 31496 11257 31524 11630
rect 31482 11248 31538 11257
rect 31392 11212 31444 11218
rect 31482 11183 31538 11192
rect 31392 11154 31444 11160
rect 31392 11008 31444 11014
rect 31392 10950 31444 10956
rect 31404 10674 31432 10950
rect 31680 10742 31708 11698
rect 31956 11354 31984 11698
rect 31944 11348 31996 11354
rect 31944 11290 31996 11296
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32232 10810 32260 11086
rect 33702 10908 34010 10917
rect 33702 10906 33708 10908
rect 33764 10906 33788 10908
rect 33844 10906 33868 10908
rect 33924 10906 33948 10908
rect 34004 10906 34010 10908
rect 33764 10854 33766 10906
rect 33946 10854 33948 10906
rect 33702 10852 33708 10854
rect 33764 10852 33788 10854
rect 33844 10852 33868 10854
rect 33924 10852 33948 10854
rect 34004 10852 34010 10854
rect 33702 10843 34010 10852
rect 32220 10804 32272 10810
rect 32220 10746 32272 10752
rect 31668 10736 31720 10742
rect 31668 10678 31720 10684
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 31392 10668 31444 10674
rect 31392 10610 31444 10616
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 27804 10464 27856 10470
rect 27804 10406 27856 10412
rect 27816 10062 27844 10406
rect 29608 10364 29916 10373
rect 29608 10362 29614 10364
rect 29670 10362 29694 10364
rect 29750 10362 29774 10364
rect 29830 10362 29854 10364
rect 29910 10362 29916 10364
rect 29670 10310 29672 10362
rect 29852 10310 29854 10362
rect 29608 10308 29614 10310
rect 29670 10308 29694 10310
rect 29750 10308 29774 10310
rect 29830 10308 29854 10310
rect 29910 10308 29916 10310
rect 29608 10299 29916 10308
rect 27804 10056 27856 10062
rect 27804 9998 27856 10004
rect 26976 9716 27028 9722
rect 26976 9658 27028 9664
rect 30024 9518 30052 10542
rect 31208 10464 31260 10470
rect 31208 10406 31260 10412
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30012 9512 30064 9518
rect 30012 9454 30064 9460
rect 30392 9450 30420 10066
rect 31220 10062 31248 10406
rect 31680 10130 31708 10678
rect 32312 10668 32364 10674
rect 32312 10610 32364 10616
rect 31668 10124 31720 10130
rect 31668 10066 31720 10072
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 30852 9722 30880 9998
rect 31576 9920 31628 9926
rect 31576 9862 31628 9868
rect 30840 9716 30892 9722
rect 30840 9658 30892 9664
rect 31588 9586 31616 9862
rect 31576 9580 31628 9586
rect 31576 9522 31628 9528
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 30380 9444 30432 9450
rect 30380 9386 30432 9392
rect 27620 9376 27672 9382
rect 27620 9318 27672 9324
rect 30472 9376 30524 9382
rect 30472 9318 30524 9324
rect 30564 9376 30616 9382
rect 30564 9318 30616 9324
rect 27252 7744 27304 7750
rect 27252 7686 27304 7692
rect 27264 6458 27292 7686
rect 27344 7336 27396 7342
rect 27344 7278 27396 7284
rect 27252 6452 27304 6458
rect 27252 6394 27304 6400
rect 27356 5914 27384 7278
rect 27528 7200 27580 7206
rect 27528 7142 27580 7148
rect 27540 6730 27568 7142
rect 27528 6724 27580 6730
rect 27528 6666 27580 6672
rect 26516 5908 26568 5914
rect 26516 5850 26568 5856
rect 27344 5908 27396 5914
rect 27344 5850 27396 5856
rect 27540 5817 27568 6666
rect 27632 6662 27660 9318
rect 29608 9276 29916 9285
rect 29608 9274 29614 9276
rect 29670 9274 29694 9276
rect 29750 9274 29774 9276
rect 29830 9274 29854 9276
rect 29910 9274 29916 9276
rect 29670 9222 29672 9274
rect 29852 9222 29854 9274
rect 29608 9220 29614 9222
rect 29670 9220 29694 9222
rect 29750 9220 29774 9222
rect 29830 9220 29854 9222
rect 29910 9220 29916 9222
rect 29608 9211 29916 9220
rect 30484 8974 30512 9318
rect 30472 8968 30524 8974
rect 30472 8910 30524 8916
rect 30104 8424 30156 8430
rect 30104 8366 30156 8372
rect 29000 8356 29052 8362
rect 29000 8298 29052 8304
rect 29012 7410 29040 8298
rect 29460 8288 29512 8294
rect 29460 8230 29512 8236
rect 29472 7818 29500 8230
rect 29608 8188 29916 8197
rect 29608 8186 29614 8188
rect 29670 8186 29694 8188
rect 29750 8186 29774 8188
rect 29830 8186 29854 8188
rect 29910 8186 29916 8188
rect 29670 8134 29672 8186
rect 29852 8134 29854 8186
rect 29608 8132 29614 8134
rect 29670 8132 29694 8134
rect 29750 8132 29774 8134
rect 29830 8132 29854 8134
rect 29910 8132 29916 8134
rect 29608 8123 29916 8132
rect 29828 7948 29880 7954
rect 29828 7890 29880 7896
rect 29460 7812 29512 7818
rect 29460 7754 29512 7760
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 28356 7200 28408 7206
rect 28356 7142 28408 7148
rect 29092 7200 29144 7206
rect 29092 7142 29144 7148
rect 28080 6860 28132 6866
rect 28080 6802 28132 6808
rect 27620 6656 27672 6662
rect 27620 6598 27672 6604
rect 27632 6390 27660 6598
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27632 5914 27660 6190
rect 27620 5908 27672 5914
rect 27620 5850 27672 5856
rect 26422 5808 26478 5817
rect 27526 5808 27582 5817
rect 26422 5743 26478 5752
rect 26792 5772 26844 5778
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26436 4826 26464 5743
rect 27526 5743 27582 5752
rect 26792 5714 26844 5720
rect 26700 5704 26752 5710
rect 26698 5672 26700 5681
rect 26752 5672 26754 5681
rect 26698 5607 26754 5616
rect 26804 5534 26832 5714
rect 26712 5506 26832 5534
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26424 4820 26476 4826
rect 26424 4762 26476 4768
rect 26516 4684 26568 4690
rect 26516 4626 26568 4632
rect 26332 4072 26384 4078
rect 26160 4032 26332 4060
rect 26332 4014 26384 4020
rect 26240 3936 26292 3942
rect 26240 3878 26292 3884
rect 26252 3534 26280 3878
rect 26344 3534 26372 4014
rect 26528 4010 26556 4626
rect 26516 4004 26568 4010
rect 26516 3946 26568 3952
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26332 3528 26384 3534
rect 26332 3470 26384 3476
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26344 3126 26372 3470
rect 26332 3120 26384 3126
rect 26332 3062 26384 3068
rect 26332 2984 26384 2990
rect 26332 2926 26384 2932
rect 26344 2582 26372 2926
rect 26436 2582 26464 3470
rect 26332 2576 26384 2582
rect 26332 2518 26384 2524
rect 26424 2576 26476 2582
rect 26424 2518 26476 2524
rect 26620 2446 26648 4966
rect 26712 2922 26740 5506
rect 27068 5296 27120 5302
rect 27068 5238 27120 5244
rect 26976 5160 27028 5166
rect 26976 5102 27028 5108
rect 26792 4820 26844 4826
rect 26792 4762 26844 4768
rect 26700 2916 26752 2922
rect 26700 2858 26752 2864
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 26056 2440 26108 2446
rect 26056 2382 26108 2388
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 26804 2378 26832 4762
rect 26884 4140 26936 4146
rect 26884 4082 26936 4088
rect 26896 2514 26924 4082
rect 26988 3194 27016 5102
rect 27080 3942 27108 5238
rect 27712 5024 27764 5030
rect 27712 4966 27764 4972
rect 27724 4690 27752 4966
rect 27712 4684 27764 4690
rect 27712 4626 27764 4632
rect 27528 4548 27580 4554
rect 27528 4490 27580 4496
rect 27896 4548 27948 4554
rect 27896 4490 27948 4496
rect 27344 4480 27396 4486
rect 27344 4422 27396 4428
rect 27160 4072 27212 4078
rect 27160 4014 27212 4020
rect 27068 3936 27120 3942
rect 27068 3878 27120 3884
rect 26976 3188 27028 3194
rect 26976 3130 27028 3136
rect 27080 3058 27108 3878
rect 27068 3052 27120 3058
rect 27068 2994 27120 3000
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 27172 2378 27200 4014
rect 27356 3738 27384 4422
rect 27344 3732 27396 3738
rect 27344 3674 27396 3680
rect 27540 2514 27568 4490
rect 27804 4480 27856 4486
rect 27804 4422 27856 4428
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 27632 2582 27660 3878
rect 27816 3058 27844 4422
rect 27908 4078 27936 4490
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 27908 3398 27936 4014
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 27804 3052 27856 3058
rect 27804 2994 27856 3000
rect 27620 2576 27672 2582
rect 27620 2518 27672 2524
rect 27528 2508 27580 2514
rect 27528 2450 27580 2456
rect 26792 2372 26844 2378
rect 26792 2314 26844 2320
rect 27160 2372 27212 2378
rect 27160 2314 27212 2320
rect 25514 2204 25822 2213
rect 25514 2202 25520 2204
rect 25576 2202 25600 2204
rect 25656 2202 25680 2204
rect 25736 2202 25760 2204
rect 25816 2202 25822 2204
rect 25576 2150 25578 2202
rect 25758 2150 25760 2202
rect 25514 2148 25520 2150
rect 25576 2148 25600 2150
rect 25656 2148 25680 2150
rect 25736 2148 25760 2150
rect 25816 2148 25822 2150
rect 25514 2139 25822 2148
rect 28092 2106 28120 6802
rect 28368 5778 28396 7142
rect 29104 6866 29132 7142
rect 29092 6860 29144 6866
rect 29092 6802 29144 6808
rect 29184 6792 29236 6798
rect 29184 6734 29236 6740
rect 28816 6248 28868 6254
rect 28816 6190 28868 6196
rect 28356 5772 28408 5778
rect 28356 5714 28408 5720
rect 28172 5704 28224 5710
rect 28172 5646 28224 5652
rect 28184 4282 28212 5646
rect 28828 5234 28856 6190
rect 29092 6112 29144 6118
rect 29092 6054 29144 6060
rect 29196 6066 29224 6734
rect 29104 5846 29132 6054
rect 29196 6038 29408 6066
rect 29092 5840 29144 5846
rect 29092 5782 29144 5788
rect 29276 5636 29328 5642
rect 29276 5578 29328 5584
rect 28908 5568 28960 5574
rect 28960 5516 29040 5534
rect 28908 5510 29040 5516
rect 28920 5506 29040 5510
rect 28816 5228 28868 5234
rect 28816 5170 28868 5176
rect 28724 5160 28776 5166
rect 28724 5102 28776 5108
rect 28172 4276 28224 4282
rect 28172 4218 28224 4224
rect 28736 4146 28764 5102
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 28632 2984 28684 2990
rect 28632 2926 28684 2932
rect 28368 2582 28396 2926
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 28540 2372 28592 2378
rect 28540 2314 28592 2320
rect 28080 2100 28132 2106
rect 28080 2042 28132 2048
rect 24320 1686 24532 1714
rect 24320 800 24348 1686
rect 27068 1556 27120 1562
rect 27068 1498 27120 1504
rect 25688 1488 25740 1494
rect 25688 1430 25740 1436
rect 25700 800 25728 1430
rect 27080 800 27108 1498
rect 28552 1170 28580 2314
rect 28644 1494 28672 2926
rect 28828 2922 28856 5170
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28816 2916 28868 2922
rect 28816 2858 28868 2864
rect 28920 2310 28948 4626
rect 29012 4146 29040 5506
rect 29092 5296 29144 5302
rect 29184 5296 29236 5302
rect 29092 5238 29144 5244
rect 29182 5264 29184 5273
rect 29236 5264 29238 5273
rect 29104 4826 29132 5238
rect 29182 5199 29238 5208
rect 29092 4820 29144 4826
rect 29092 4762 29144 4768
rect 29288 4282 29316 5578
rect 29380 4808 29408 6038
rect 29472 5778 29500 7754
rect 29840 7410 29868 7890
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 29608 7100 29916 7109
rect 29608 7098 29614 7100
rect 29670 7098 29694 7100
rect 29750 7098 29774 7100
rect 29830 7098 29854 7100
rect 29910 7098 29916 7100
rect 29670 7046 29672 7098
rect 29852 7046 29854 7098
rect 29608 7044 29614 7046
rect 29670 7044 29694 7046
rect 29750 7044 29774 7046
rect 29830 7044 29854 7046
rect 29910 7044 29916 7046
rect 29608 7035 29916 7044
rect 29608 6012 29916 6021
rect 29608 6010 29614 6012
rect 29670 6010 29694 6012
rect 29750 6010 29774 6012
rect 29830 6010 29854 6012
rect 29910 6010 29916 6012
rect 29670 5958 29672 6010
rect 29852 5958 29854 6010
rect 29608 5956 29614 5958
rect 29670 5956 29694 5958
rect 29750 5956 29774 5958
rect 29830 5956 29854 5958
rect 29910 5956 29916 5958
rect 29608 5947 29916 5956
rect 29460 5772 29512 5778
rect 29460 5714 29512 5720
rect 29920 5568 29972 5574
rect 29972 5516 30052 5534
rect 29920 5510 30052 5516
rect 29932 5506 30052 5510
rect 30024 5098 30052 5506
rect 30116 5370 30144 8366
rect 30576 8022 30604 9318
rect 31128 8634 31156 9454
rect 31680 9042 31708 10066
rect 32324 9654 32352 10610
rect 33324 10600 33376 10606
rect 33324 10542 33376 10548
rect 33048 9920 33100 9926
rect 33048 9862 33100 9868
rect 32312 9648 32364 9654
rect 32312 9590 32364 9596
rect 33060 9586 33088 9862
rect 33336 9625 33364 10542
rect 33702 9820 34010 9829
rect 33702 9818 33708 9820
rect 33764 9818 33788 9820
rect 33844 9818 33868 9820
rect 33924 9818 33948 9820
rect 34004 9818 34010 9820
rect 33764 9766 33766 9818
rect 33946 9766 33948 9818
rect 33702 9764 33708 9766
rect 33764 9764 33788 9766
rect 33844 9764 33868 9766
rect 33924 9764 33948 9766
rect 34004 9764 34010 9766
rect 33702 9755 34010 9764
rect 33322 9616 33378 9625
rect 33048 9580 33100 9586
rect 33322 9551 33378 9560
rect 33048 9522 33100 9528
rect 31668 9036 31720 9042
rect 31668 8978 31720 8984
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 31576 8968 31628 8974
rect 31576 8910 31628 8916
rect 31208 8832 31260 8838
rect 31208 8774 31260 8780
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 31220 8430 31248 8774
rect 31312 8537 31340 8910
rect 31588 8566 31616 8910
rect 31576 8560 31628 8566
rect 31298 8528 31354 8537
rect 31576 8502 31628 8508
rect 31298 8463 31354 8472
rect 31208 8424 31260 8430
rect 31208 8366 31260 8372
rect 31300 8424 31352 8430
rect 31300 8366 31352 8372
rect 31312 8022 31340 8366
rect 30564 8016 30616 8022
rect 30564 7958 30616 7964
rect 31300 8016 31352 8022
rect 31300 7958 31352 7964
rect 31680 7954 31708 8978
rect 33702 8732 34010 8741
rect 33702 8730 33708 8732
rect 33764 8730 33788 8732
rect 33844 8730 33868 8732
rect 33924 8730 33948 8732
rect 34004 8730 34010 8732
rect 33764 8678 33766 8730
rect 33946 8678 33948 8730
rect 33702 8676 33708 8678
rect 33764 8676 33788 8678
rect 33844 8676 33868 8678
rect 33924 8676 33948 8678
rect 34004 8676 34010 8678
rect 33702 8667 34010 8676
rect 32036 8084 32088 8090
rect 32036 8026 32088 8032
rect 31668 7948 31720 7954
rect 31668 7890 31720 7896
rect 31024 7404 31076 7410
rect 31024 7346 31076 7352
rect 31036 6798 31064 7346
rect 31208 7336 31260 7342
rect 31208 7278 31260 7284
rect 30564 6792 30616 6798
rect 30564 6734 30616 6740
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 30392 5534 30420 5782
rect 30484 5778 30512 6598
rect 30576 6390 30604 6734
rect 30760 6458 30788 6734
rect 30748 6452 30800 6458
rect 30748 6394 30800 6400
rect 30564 6384 30616 6390
rect 30564 6326 30616 6332
rect 30932 6316 30984 6322
rect 30932 6258 30984 6264
rect 30746 5808 30802 5817
rect 30472 5772 30524 5778
rect 30746 5743 30802 5752
rect 30472 5714 30524 5720
rect 30392 5506 30512 5534
rect 30104 5364 30156 5370
rect 30104 5306 30156 5312
rect 30104 5160 30156 5166
rect 30104 5102 30156 5108
rect 30012 5092 30064 5098
rect 30012 5034 30064 5040
rect 29608 4924 29916 4933
rect 29608 4922 29614 4924
rect 29670 4922 29694 4924
rect 29750 4922 29774 4924
rect 29830 4922 29854 4924
rect 29910 4922 29916 4924
rect 29670 4870 29672 4922
rect 29852 4870 29854 4922
rect 29608 4868 29614 4870
rect 29670 4868 29694 4870
rect 29750 4868 29774 4870
rect 29830 4868 29854 4870
rect 29910 4868 29916 4870
rect 29608 4859 29916 4868
rect 29380 4780 29776 4808
rect 29748 4622 29776 4780
rect 29552 4616 29604 4622
rect 29552 4558 29604 4564
rect 29736 4616 29788 4622
rect 29736 4558 29788 4564
rect 29276 4276 29328 4282
rect 29276 4218 29328 4224
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 29564 3942 29592 4558
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29608 3836 29916 3845
rect 29608 3834 29614 3836
rect 29670 3834 29694 3836
rect 29750 3834 29774 3836
rect 29830 3834 29854 3836
rect 29910 3834 29916 3836
rect 29670 3782 29672 3834
rect 29852 3782 29854 3834
rect 29608 3780 29614 3782
rect 29670 3780 29694 3782
rect 29750 3780 29774 3782
rect 29830 3780 29854 3782
rect 29910 3780 29916 3782
rect 29608 3771 29916 3780
rect 30024 3670 30052 5034
rect 30012 3664 30064 3670
rect 30012 3606 30064 3612
rect 29920 3528 29972 3534
rect 29920 3470 29972 3476
rect 29932 3058 29960 3470
rect 29920 3052 29972 3058
rect 29920 2994 29972 3000
rect 30012 2984 30064 2990
rect 30012 2926 30064 2932
rect 29608 2748 29916 2757
rect 29608 2746 29614 2748
rect 29670 2746 29694 2748
rect 29750 2746 29774 2748
rect 29830 2746 29854 2748
rect 29910 2746 29916 2748
rect 29670 2694 29672 2746
rect 29852 2694 29854 2746
rect 29608 2692 29614 2694
rect 29670 2692 29694 2694
rect 29750 2692 29774 2694
rect 29830 2692 29854 2694
rect 29910 2692 29916 2694
rect 29608 2683 29916 2692
rect 29552 2644 29604 2650
rect 29552 2586 29604 2592
rect 28908 2304 28960 2310
rect 28908 2246 28960 2252
rect 29564 1737 29592 2586
rect 30024 2514 30052 2926
rect 30012 2508 30064 2514
rect 30012 2450 30064 2456
rect 29550 1728 29606 1737
rect 29550 1663 29606 1672
rect 28632 1488 28684 1494
rect 28632 1430 28684 1436
rect 28460 1142 28580 1170
rect 28460 800 28488 1142
rect 29840 870 29960 898
rect 29840 800 29868 870
rect 17512 734 17908 762
rect 18786 0 18842 800
rect 20166 0 20222 800
rect 21546 0 21602 800
rect 22926 0 22982 800
rect 24306 0 24362 800
rect 25686 0 25742 800
rect 27066 0 27122 800
rect 28446 0 28502 800
rect 29826 0 29882 800
rect 29932 762 29960 870
rect 30116 762 30144 5102
rect 30196 4480 30248 4486
rect 30196 4422 30248 4428
rect 30208 3534 30236 4422
rect 30196 3528 30248 3534
rect 30196 3470 30248 3476
rect 30196 2984 30248 2990
rect 30196 2926 30248 2932
rect 30208 1562 30236 2926
rect 30484 2446 30512 5506
rect 30760 4826 30788 5743
rect 30748 4820 30800 4826
rect 30748 4762 30800 4768
rect 30944 4690 30972 6258
rect 31116 5704 31168 5710
rect 31116 5646 31168 5652
rect 30932 4684 30984 4690
rect 30932 4626 30984 4632
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 30852 3194 30880 4082
rect 31128 4078 31156 5646
rect 31116 4072 31168 4078
rect 31116 4014 31168 4020
rect 31116 3460 31168 3466
rect 31116 3402 31168 3408
rect 30840 3188 30892 3194
rect 30840 3130 30892 3136
rect 31128 2446 31156 3402
rect 30472 2440 30524 2446
rect 30472 2382 30524 2388
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 30196 1556 30248 1562
rect 30196 1498 30248 1504
rect 31220 800 31248 7278
rect 31680 6322 31708 7890
rect 32048 6390 32076 8026
rect 33702 7644 34010 7653
rect 33702 7642 33708 7644
rect 33764 7642 33788 7644
rect 33844 7642 33868 7644
rect 33924 7642 33948 7644
rect 34004 7642 34010 7644
rect 33764 7590 33766 7642
rect 33946 7590 33948 7642
rect 33702 7588 33708 7590
rect 33764 7588 33788 7590
rect 33844 7588 33868 7590
rect 33924 7588 33948 7590
rect 34004 7588 34010 7590
rect 33702 7579 34010 7588
rect 32496 7336 32548 7342
rect 32496 7278 32548 7284
rect 32508 6798 32536 7278
rect 33322 7168 33378 7177
rect 33322 7103 33378 7112
rect 33336 6866 33364 7103
rect 33324 6860 33376 6866
rect 33324 6802 33376 6808
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32588 6724 32640 6730
rect 32588 6666 32640 6672
rect 32036 6384 32088 6390
rect 32036 6326 32088 6332
rect 31668 6316 31720 6322
rect 31668 6258 31720 6264
rect 31944 6316 31996 6322
rect 31944 6258 31996 6264
rect 31484 6248 31536 6254
rect 31484 6190 31536 6196
rect 31496 5817 31524 6190
rect 31760 5908 31812 5914
rect 31760 5850 31812 5856
rect 31482 5808 31538 5817
rect 31482 5743 31538 5752
rect 31576 5636 31628 5642
rect 31576 5578 31628 5584
rect 31588 4593 31616 5578
rect 31574 4584 31630 4593
rect 31574 4519 31630 4528
rect 31668 4548 31720 4554
rect 31668 4490 31720 4496
rect 31680 4078 31708 4490
rect 31772 4214 31800 5850
rect 31956 5778 31984 6258
rect 32128 6248 32180 6254
rect 32128 6190 32180 6196
rect 31944 5772 31996 5778
rect 31944 5714 31996 5720
rect 32036 5704 32088 5710
rect 32036 5646 32088 5652
rect 31944 5228 31996 5234
rect 31944 5170 31996 5176
rect 31852 4548 31904 4554
rect 31852 4490 31904 4496
rect 31760 4208 31812 4214
rect 31760 4150 31812 4156
rect 31668 4072 31720 4078
rect 31668 4014 31720 4020
rect 31864 3738 31892 4490
rect 31852 3732 31904 3738
rect 31852 3674 31904 3680
rect 31956 3534 31984 5170
rect 32048 4690 32076 5646
rect 32140 5234 32168 6190
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32036 4684 32088 4690
rect 32036 4626 32088 4632
rect 32140 4146 32168 5170
rect 32218 4720 32274 4729
rect 32218 4655 32274 4664
rect 32232 4622 32260 4655
rect 32220 4616 32272 4622
rect 32220 4558 32272 4564
rect 32128 4140 32180 4146
rect 32128 4082 32180 4088
rect 31760 3528 31812 3534
rect 31760 3470 31812 3476
rect 31944 3528 31996 3534
rect 31944 3470 31996 3476
rect 31772 2650 31800 3470
rect 31852 3392 31904 3398
rect 31852 3334 31904 3340
rect 31864 3126 31892 3334
rect 31852 3120 31904 3126
rect 31852 3062 31904 3068
rect 32140 3058 32168 4082
rect 32600 3194 32628 6666
rect 33702 6556 34010 6565
rect 33702 6554 33708 6556
rect 33764 6554 33788 6556
rect 33844 6554 33868 6556
rect 33924 6554 33948 6556
rect 34004 6554 34010 6556
rect 33764 6502 33766 6554
rect 33946 6502 33948 6554
rect 33702 6500 33708 6502
rect 33764 6500 33788 6502
rect 33844 6500 33868 6502
rect 33924 6500 33948 6502
rect 34004 6500 34010 6502
rect 33702 6491 34010 6500
rect 34060 6112 34112 6118
rect 34060 6054 34112 6060
rect 32864 5704 32916 5710
rect 32864 5646 32916 5652
rect 33506 5672 33562 5681
rect 32876 3738 32904 5646
rect 33506 5607 33562 5616
rect 33520 5370 33548 5607
rect 33702 5468 34010 5477
rect 33702 5466 33708 5468
rect 33764 5466 33788 5468
rect 33844 5466 33868 5468
rect 33924 5466 33948 5468
rect 34004 5466 34010 5468
rect 33764 5414 33766 5466
rect 33946 5414 33948 5466
rect 33702 5412 33708 5414
rect 33764 5412 33788 5414
rect 33844 5412 33868 5414
rect 33924 5412 33948 5414
rect 34004 5412 34010 5414
rect 33702 5403 34010 5412
rect 33508 5364 33560 5370
rect 33508 5306 33560 5312
rect 33702 4380 34010 4389
rect 33702 4378 33708 4380
rect 33764 4378 33788 4380
rect 33844 4378 33868 4380
rect 33924 4378 33948 4380
rect 34004 4378 34010 4380
rect 33764 4326 33766 4378
rect 33946 4326 33948 4378
rect 33702 4324 33708 4326
rect 33764 4324 33788 4326
rect 33844 4324 33868 4326
rect 33924 4324 33948 4326
rect 34004 4324 34010 4326
rect 33702 4315 34010 4324
rect 32864 3732 32916 3738
rect 32864 3674 32916 3680
rect 33508 3392 33560 3398
rect 33508 3334 33560 3340
rect 32588 3188 32640 3194
rect 32588 3130 32640 3136
rect 33520 3097 33548 3334
rect 33702 3292 34010 3301
rect 33702 3290 33708 3292
rect 33764 3290 33788 3292
rect 33844 3290 33868 3292
rect 33924 3290 33948 3292
rect 34004 3290 34010 3292
rect 33764 3238 33766 3290
rect 33946 3238 33948 3290
rect 33702 3236 33708 3238
rect 33764 3236 33788 3238
rect 33844 3236 33868 3238
rect 33924 3236 33948 3238
rect 34004 3236 34010 3238
rect 33702 3227 34010 3236
rect 33506 3088 33562 3097
rect 32128 3052 32180 3058
rect 33506 3023 33562 3032
rect 32128 2994 32180 3000
rect 31760 2644 31812 2650
rect 31760 2586 31812 2592
rect 32588 2304 32640 2310
rect 32588 2246 32640 2252
rect 32600 800 32628 2246
rect 33702 2204 34010 2213
rect 33702 2202 33708 2204
rect 33764 2202 33788 2204
rect 33844 2202 33868 2204
rect 33924 2202 33948 2204
rect 34004 2202 34010 2204
rect 33764 2150 33766 2202
rect 33946 2150 33948 2202
rect 33702 2148 33708 2150
rect 33764 2148 33788 2150
rect 33844 2148 33868 2150
rect 33924 2148 33948 2150
rect 34004 2148 34010 2150
rect 33702 2139 34010 2148
rect 34072 1394 34100 6054
rect 33980 1366 34100 1394
rect 33980 800 34008 1366
rect 29932 734 30144 762
rect 31206 0 31262 800
rect 32586 0 32642 800
rect 33966 0 34022 800
<< via2 >>
rect 1398 30232 1454 30288
rect 5050 32122 5106 32124
rect 5130 32122 5186 32124
rect 5210 32122 5266 32124
rect 5290 32122 5346 32124
rect 5050 32070 5096 32122
rect 5096 32070 5106 32122
rect 5130 32070 5160 32122
rect 5160 32070 5172 32122
rect 5172 32070 5186 32122
rect 5210 32070 5224 32122
rect 5224 32070 5236 32122
rect 5236 32070 5266 32122
rect 5290 32070 5300 32122
rect 5300 32070 5346 32122
rect 5050 32068 5106 32070
rect 5130 32068 5186 32070
rect 5210 32068 5266 32070
rect 5290 32068 5346 32070
rect 4066 31592 4122 31648
rect 2778 27512 2834 27568
rect 1582 26152 1638 26208
rect 938 23432 994 23488
rect 3330 28872 3386 28928
rect 2778 24792 2834 24848
rect 5050 31034 5106 31036
rect 5130 31034 5186 31036
rect 5210 31034 5266 31036
rect 5290 31034 5346 31036
rect 5050 30982 5096 31034
rect 5096 30982 5106 31034
rect 5130 30982 5160 31034
rect 5160 30982 5172 31034
rect 5172 30982 5186 31034
rect 5210 30982 5224 31034
rect 5224 30982 5236 31034
rect 5236 30982 5266 31034
rect 5290 30982 5300 31034
rect 5300 30982 5346 31034
rect 5050 30980 5106 30982
rect 5130 30980 5186 30982
rect 5210 30980 5266 30982
rect 5290 30980 5346 30982
rect 5050 29946 5106 29948
rect 5130 29946 5186 29948
rect 5210 29946 5266 29948
rect 5290 29946 5346 29948
rect 5050 29894 5096 29946
rect 5096 29894 5106 29946
rect 5130 29894 5160 29946
rect 5160 29894 5172 29946
rect 5172 29894 5186 29946
rect 5210 29894 5224 29946
rect 5224 29894 5236 29946
rect 5236 29894 5266 29946
rect 5290 29894 5300 29946
rect 5300 29894 5346 29946
rect 5050 29892 5106 29894
rect 5130 29892 5186 29894
rect 5210 29892 5266 29894
rect 5290 29892 5346 29894
rect 5050 28858 5106 28860
rect 5130 28858 5186 28860
rect 5210 28858 5266 28860
rect 5290 28858 5346 28860
rect 5050 28806 5096 28858
rect 5096 28806 5106 28858
rect 5130 28806 5160 28858
rect 5160 28806 5172 28858
rect 5172 28806 5186 28858
rect 5210 28806 5224 28858
rect 5224 28806 5236 28858
rect 5236 28806 5266 28858
rect 5290 28806 5300 28858
rect 5300 28806 5346 28858
rect 5050 28804 5106 28806
rect 5130 28804 5186 28806
rect 5210 28804 5266 28806
rect 5290 28804 5346 28806
rect 5050 27770 5106 27772
rect 5130 27770 5186 27772
rect 5210 27770 5266 27772
rect 5290 27770 5346 27772
rect 5050 27718 5096 27770
rect 5096 27718 5106 27770
rect 5130 27718 5160 27770
rect 5160 27718 5172 27770
rect 5172 27718 5186 27770
rect 5210 27718 5224 27770
rect 5224 27718 5236 27770
rect 5236 27718 5266 27770
rect 5290 27718 5300 27770
rect 5300 27718 5346 27770
rect 5050 27716 5106 27718
rect 5130 27716 5186 27718
rect 5210 27716 5266 27718
rect 5290 27716 5346 27718
rect 9144 32666 9200 32668
rect 9224 32666 9280 32668
rect 9304 32666 9360 32668
rect 9384 32666 9440 32668
rect 9144 32614 9190 32666
rect 9190 32614 9200 32666
rect 9224 32614 9254 32666
rect 9254 32614 9266 32666
rect 9266 32614 9280 32666
rect 9304 32614 9318 32666
rect 9318 32614 9330 32666
rect 9330 32614 9360 32666
rect 9384 32614 9394 32666
rect 9394 32614 9440 32666
rect 9144 32612 9200 32614
rect 9224 32612 9280 32614
rect 9304 32612 9360 32614
rect 9384 32612 9440 32614
rect 9144 31578 9200 31580
rect 9224 31578 9280 31580
rect 9304 31578 9360 31580
rect 9384 31578 9440 31580
rect 9144 31526 9190 31578
rect 9190 31526 9200 31578
rect 9224 31526 9254 31578
rect 9254 31526 9266 31578
rect 9266 31526 9280 31578
rect 9304 31526 9318 31578
rect 9318 31526 9330 31578
rect 9330 31526 9360 31578
rect 9384 31526 9394 31578
rect 9394 31526 9440 31578
rect 9144 31524 9200 31526
rect 9224 31524 9280 31526
rect 9304 31524 9360 31526
rect 9384 31524 9440 31526
rect 9144 30490 9200 30492
rect 9224 30490 9280 30492
rect 9304 30490 9360 30492
rect 9384 30490 9440 30492
rect 9144 30438 9190 30490
rect 9190 30438 9200 30490
rect 9224 30438 9254 30490
rect 9254 30438 9266 30490
rect 9266 30438 9280 30490
rect 9304 30438 9318 30490
rect 9318 30438 9330 30490
rect 9330 30438 9360 30490
rect 9384 30438 9394 30490
rect 9394 30438 9440 30490
rect 9144 30436 9200 30438
rect 9224 30436 9280 30438
rect 9304 30436 9360 30438
rect 9384 30436 9440 30438
rect 13238 32122 13294 32124
rect 13318 32122 13374 32124
rect 13398 32122 13454 32124
rect 13478 32122 13534 32124
rect 13238 32070 13284 32122
rect 13284 32070 13294 32122
rect 13318 32070 13348 32122
rect 13348 32070 13360 32122
rect 13360 32070 13374 32122
rect 13398 32070 13412 32122
rect 13412 32070 13424 32122
rect 13424 32070 13454 32122
rect 13478 32070 13488 32122
rect 13488 32070 13534 32122
rect 13238 32068 13294 32070
rect 13318 32068 13374 32070
rect 13398 32068 13454 32070
rect 13478 32068 13534 32070
rect 13238 31034 13294 31036
rect 13318 31034 13374 31036
rect 13398 31034 13454 31036
rect 13478 31034 13534 31036
rect 13238 30982 13284 31034
rect 13284 30982 13294 31034
rect 13318 30982 13348 31034
rect 13348 30982 13360 31034
rect 13360 30982 13374 31034
rect 13398 30982 13412 31034
rect 13412 30982 13424 31034
rect 13424 30982 13454 31034
rect 13478 30982 13488 31034
rect 13488 30982 13534 31034
rect 13238 30980 13294 30982
rect 13318 30980 13374 30982
rect 13398 30980 13454 30982
rect 13478 30980 13534 30982
rect 5050 26682 5106 26684
rect 5130 26682 5186 26684
rect 5210 26682 5266 26684
rect 5290 26682 5346 26684
rect 5050 26630 5096 26682
rect 5096 26630 5106 26682
rect 5130 26630 5160 26682
rect 5160 26630 5172 26682
rect 5172 26630 5186 26682
rect 5210 26630 5224 26682
rect 5224 26630 5236 26682
rect 5236 26630 5266 26682
rect 5290 26630 5300 26682
rect 5300 26630 5346 26682
rect 5050 26628 5106 26630
rect 5130 26628 5186 26630
rect 5210 26628 5266 26630
rect 5290 26628 5346 26630
rect 5050 25594 5106 25596
rect 5130 25594 5186 25596
rect 5210 25594 5266 25596
rect 5290 25594 5346 25596
rect 5050 25542 5096 25594
rect 5096 25542 5106 25594
rect 5130 25542 5160 25594
rect 5160 25542 5172 25594
rect 5172 25542 5186 25594
rect 5210 25542 5224 25594
rect 5224 25542 5236 25594
rect 5236 25542 5266 25594
rect 5290 25542 5300 25594
rect 5300 25542 5346 25594
rect 5050 25540 5106 25542
rect 5130 25540 5186 25542
rect 5210 25540 5266 25542
rect 5290 25540 5346 25542
rect 1582 22344 1638 22400
rect 938 20712 994 20768
rect 938 19372 994 19408
rect 938 19352 940 19372
rect 940 19352 992 19372
rect 992 19352 994 19372
rect 1306 17992 1362 18048
rect 1582 16632 1638 16688
rect 1582 15272 1638 15328
rect 1306 13912 1362 13968
rect 1582 12416 1638 12472
rect 1306 11192 1362 11248
rect 1582 9696 1638 9752
rect 1582 8336 1638 8392
rect 1582 6976 1638 7032
rect 1306 5752 1362 5808
rect 1582 4120 1638 4176
rect 5050 24506 5106 24508
rect 5130 24506 5186 24508
rect 5210 24506 5266 24508
rect 5290 24506 5346 24508
rect 5050 24454 5096 24506
rect 5096 24454 5106 24506
rect 5130 24454 5160 24506
rect 5160 24454 5172 24506
rect 5172 24454 5186 24506
rect 5210 24454 5224 24506
rect 5224 24454 5236 24506
rect 5236 24454 5266 24506
rect 5290 24454 5300 24506
rect 5300 24454 5346 24506
rect 5050 24452 5106 24454
rect 5130 24452 5186 24454
rect 5210 24452 5266 24454
rect 5290 24452 5346 24454
rect 5050 23418 5106 23420
rect 5130 23418 5186 23420
rect 5210 23418 5266 23420
rect 5290 23418 5346 23420
rect 5050 23366 5096 23418
rect 5096 23366 5106 23418
rect 5130 23366 5160 23418
rect 5160 23366 5172 23418
rect 5172 23366 5186 23418
rect 5210 23366 5224 23418
rect 5224 23366 5236 23418
rect 5236 23366 5266 23418
rect 5290 23366 5300 23418
rect 5300 23366 5346 23418
rect 5050 23364 5106 23366
rect 5130 23364 5186 23366
rect 5210 23364 5266 23366
rect 5290 23364 5346 23366
rect 5050 22330 5106 22332
rect 5130 22330 5186 22332
rect 5210 22330 5266 22332
rect 5290 22330 5346 22332
rect 5050 22278 5096 22330
rect 5096 22278 5106 22330
rect 5130 22278 5160 22330
rect 5160 22278 5172 22330
rect 5172 22278 5186 22330
rect 5210 22278 5224 22330
rect 5224 22278 5236 22330
rect 5236 22278 5266 22330
rect 5290 22278 5300 22330
rect 5300 22278 5346 22330
rect 5050 22276 5106 22278
rect 5130 22276 5186 22278
rect 5210 22276 5266 22278
rect 5290 22276 5346 22278
rect 5050 21242 5106 21244
rect 5130 21242 5186 21244
rect 5210 21242 5266 21244
rect 5290 21242 5346 21244
rect 5050 21190 5096 21242
rect 5096 21190 5106 21242
rect 5130 21190 5160 21242
rect 5160 21190 5172 21242
rect 5172 21190 5186 21242
rect 5210 21190 5224 21242
rect 5224 21190 5236 21242
rect 5236 21190 5266 21242
rect 5290 21190 5300 21242
rect 5300 21190 5346 21242
rect 5050 21188 5106 21190
rect 5130 21188 5186 21190
rect 5210 21188 5266 21190
rect 5290 21188 5346 21190
rect 5050 20154 5106 20156
rect 5130 20154 5186 20156
rect 5210 20154 5266 20156
rect 5290 20154 5346 20156
rect 5050 20102 5096 20154
rect 5096 20102 5106 20154
rect 5130 20102 5160 20154
rect 5160 20102 5172 20154
rect 5172 20102 5186 20154
rect 5210 20102 5224 20154
rect 5224 20102 5236 20154
rect 5236 20102 5266 20154
rect 5290 20102 5300 20154
rect 5300 20102 5346 20154
rect 5050 20100 5106 20102
rect 5130 20100 5186 20102
rect 5210 20100 5266 20102
rect 5290 20100 5346 20102
rect 5050 19066 5106 19068
rect 5130 19066 5186 19068
rect 5210 19066 5266 19068
rect 5290 19066 5346 19068
rect 5050 19014 5096 19066
rect 5096 19014 5106 19066
rect 5130 19014 5160 19066
rect 5160 19014 5172 19066
rect 5172 19014 5186 19066
rect 5210 19014 5224 19066
rect 5224 19014 5236 19066
rect 5236 19014 5266 19066
rect 5290 19014 5300 19066
rect 5300 19014 5346 19066
rect 5050 19012 5106 19014
rect 5130 19012 5186 19014
rect 5210 19012 5266 19014
rect 5290 19012 5346 19014
rect 9144 29402 9200 29404
rect 9224 29402 9280 29404
rect 9304 29402 9360 29404
rect 9384 29402 9440 29404
rect 9144 29350 9190 29402
rect 9190 29350 9200 29402
rect 9224 29350 9254 29402
rect 9254 29350 9266 29402
rect 9266 29350 9280 29402
rect 9304 29350 9318 29402
rect 9318 29350 9330 29402
rect 9330 29350 9360 29402
rect 9384 29350 9394 29402
rect 9394 29350 9440 29402
rect 9144 29348 9200 29350
rect 9224 29348 9280 29350
rect 9304 29348 9360 29350
rect 9384 29348 9440 29350
rect 9144 28314 9200 28316
rect 9224 28314 9280 28316
rect 9304 28314 9360 28316
rect 9384 28314 9440 28316
rect 9144 28262 9190 28314
rect 9190 28262 9200 28314
rect 9224 28262 9254 28314
rect 9254 28262 9266 28314
rect 9266 28262 9280 28314
rect 9304 28262 9318 28314
rect 9318 28262 9330 28314
rect 9330 28262 9360 28314
rect 9384 28262 9394 28314
rect 9394 28262 9440 28314
rect 9144 28260 9200 28262
rect 9224 28260 9280 28262
rect 9304 28260 9360 28262
rect 9384 28260 9440 28262
rect 9144 27226 9200 27228
rect 9224 27226 9280 27228
rect 9304 27226 9360 27228
rect 9384 27226 9440 27228
rect 9144 27174 9190 27226
rect 9190 27174 9200 27226
rect 9224 27174 9254 27226
rect 9254 27174 9266 27226
rect 9266 27174 9280 27226
rect 9304 27174 9318 27226
rect 9318 27174 9330 27226
rect 9330 27174 9360 27226
rect 9384 27174 9394 27226
rect 9394 27174 9440 27226
rect 9144 27172 9200 27174
rect 9224 27172 9280 27174
rect 9304 27172 9360 27174
rect 9384 27172 9440 27174
rect 9144 26138 9200 26140
rect 9224 26138 9280 26140
rect 9304 26138 9360 26140
rect 9384 26138 9440 26140
rect 9144 26086 9190 26138
rect 9190 26086 9200 26138
rect 9224 26086 9254 26138
rect 9254 26086 9266 26138
rect 9266 26086 9280 26138
rect 9304 26086 9318 26138
rect 9318 26086 9330 26138
rect 9330 26086 9360 26138
rect 9384 26086 9394 26138
rect 9394 26086 9440 26138
rect 9144 26084 9200 26086
rect 9224 26084 9280 26086
rect 9304 26084 9360 26086
rect 9384 26084 9440 26086
rect 9144 25050 9200 25052
rect 9224 25050 9280 25052
rect 9304 25050 9360 25052
rect 9384 25050 9440 25052
rect 9144 24998 9190 25050
rect 9190 24998 9200 25050
rect 9224 24998 9254 25050
rect 9254 24998 9266 25050
rect 9266 24998 9280 25050
rect 9304 24998 9318 25050
rect 9318 24998 9330 25050
rect 9330 24998 9360 25050
rect 9384 24998 9394 25050
rect 9394 24998 9440 25050
rect 9144 24996 9200 24998
rect 9224 24996 9280 24998
rect 9304 24996 9360 24998
rect 9384 24996 9440 24998
rect 17332 32666 17388 32668
rect 17412 32666 17468 32668
rect 17492 32666 17548 32668
rect 17572 32666 17628 32668
rect 17332 32614 17378 32666
rect 17378 32614 17388 32666
rect 17412 32614 17442 32666
rect 17442 32614 17454 32666
rect 17454 32614 17468 32666
rect 17492 32614 17506 32666
rect 17506 32614 17518 32666
rect 17518 32614 17548 32666
rect 17572 32614 17582 32666
rect 17582 32614 17628 32666
rect 17332 32612 17388 32614
rect 17412 32612 17468 32614
rect 17492 32612 17548 32614
rect 17572 32612 17628 32614
rect 13238 29946 13294 29948
rect 13318 29946 13374 29948
rect 13398 29946 13454 29948
rect 13478 29946 13534 29948
rect 13238 29894 13284 29946
rect 13284 29894 13294 29946
rect 13318 29894 13348 29946
rect 13348 29894 13360 29946
rect 13360 29894 13374 29946
rect 13398 29894 13412 29946
rect 13412 29894 13424 29946
rect 13424 29894 13454 29946
rect 13478 29894 13488 29946
rect 13488 29894 13534 29946
rect 13238 29892 13294 29894
rect 13318 29892 13374 29894
rect 13398 29892 13454 29894
rect 13478 29892 13534 29894
rect 13238 28858 13294 28860
rect 13318 28858 13374 28860
rect 13398 28858 13454 28860
rect 13478 28858 13534 28860
rect 13238 28806 13284 28858
rect 13284 28806 13294 28858
rect 13318 28806 13348 28858
rect 13348 28806 13360 28858
rect 13360 28806 13374 28858
rect 13398 28806 13412 28858
rect 13412 28806 13424 28858
rect 13424 28806 13454 28858
rect 13478 28806 13488 28858
rect 13488 28806 13534 28858
rect 13238 28804 13294 28806
rect 13318 28804 13374 28806
rect 13398 28804 13454 28806
rect 13478 28804 13534 28806
rect 13238 27770 13294 27772
rect 13318 27770 13374 27772
rect 13398 27770 13454 27772
rect 13478 27770 13534 27772
rect 13238 27718 13284 27770
rect 13284 27718 13294 27770
rect 13318 27718 13348 27770
rect 13348 27718 13360 27770
rect 13360 27718 13374 27770
rect 13398 27718 13412 27770
rect 13412 27718 13424 27770
rect 13424 27718 13454 27770
rect 13478 27718 13488 27770
rect 13488 27718 13534 27770
rect 13238 27716 13294 27718
rect 13318 27716 13374 27718
rect 13398 27716 13454 27718
rect 13478 27716 13534 27718
rect 13238 26682 13294 26684
rect 13318 26682 13374 26684
rect 13398 26682 13454 26684
rect 13478 26682 13534 26684
rect 13238 26630 13284 26682
rect 13284 26630 13294 26682
rect 13318 26630 13348 26682
rect 13348 26630 13360 26682
rect 13360 26630 13374 26682
rect 13398 26630 13412 26682
rect 13412 26630 13424 26682
rect 13424 26630 13454 26682
rect 13478 26630 13488 26682
rect 13488 26630 13534 26682
rect 13238 26628 13294 26630
rect 13318 26628 13374 26630
rect 13398 26628 13454 26630
rect 13478 26628 13534 26630
rect 13238 25594 13294 25596
rect 13318 25594 13374 25596
rect 13398 25594 13454 25596
rect 13478 25594 13534 25596
rect 13238 25542 13284 25594
rect 13284 25542 13294 25594
rect 13318 25542 13348 25594
rect 13348 25542 13360 25594
rect 13360 25542 13374 25594
rect 13398 25542 13412 25594
rect 13412 25542 13424 25594
rect 13424 25542 13454 25594
rect 13478 25542 13488 25594
rect 13488 25542 13534 25594
rect 13238 25540 13294 25542
rect 13318 25540 13374 25542
rect 13398 25540 13454 25542
rect 13478 25540 13534 25542
rect 17332 31578 17388 31580
rect 17412 31578 17468 31580
rect 17492 31578 17548 31580
rect 17572 31578 17628 31580
rect 17332 31526 17378 31578
rect 17378 31526 17388 31578
rect 17412 31526 17442 31578
rect 17442 31526 17454 31578
rect 17454 31526 17468 31578
rect 17492 31526 17506 31578
rect 17506 31526 17518 31578
rect 17518 31526 17548 31578
rect 17572 31526 17582 31578
rect 17582 31526 17628 31578
rect 17332 31524 17388 31526
rect 17412 31524 17468 31526
rect 17492 31524 17548 31526
rect 17572 31524 17628 31526
rect 17332 30490 17388 30492
rect 17412 30490 17468 30492
rect 17492 30490 17548 30492
rect 17572 30490 17628 30492
rect 17332 30438 17378 30490
rect 17378 30438 17388 30490
rect 17412 30438 17442 30490
rect 17442 30438 17454 30490
rect 17454 30438 17468 30490
rect 17492 30438 17506 30490
rect 17506 30438 17518 30490
rect 17518 30438 17548 30490
rect 17572 30438 17582 30490
rect 17582 30438 17628 30490
rect 17332 30436 17388 30438
rect 17412 30436 17468 30438
rect 17492 30436 17548 30438
rect 17572 30436 17628 30438
rect 21426 32122 21482 32124
rect 21506 32122 21562 32124
rect 21586 32122 21642 32124
rect 21666 32122 21722 32124
rect 21426 32070 21472 32122
rect 21472 32070 21482 32122
rect 21506 32070 21536 32122
rect 21536 32070 21548 32122
rect 21548 32070 21562 32122
rect 21586 32070 21600 32122
rect 21600 32070 21612 32122
rect 21612 32070 21642 32122
rect 21666 32070 21676 32122
rect 21676 32070 21722 32122
rect 21426 32068 21482 32070
rect 21506 32068 21562 32070
rect 21586 32068 21642 32070
rect 21666 32068 21722 32070
rect 21426 31034 21482 31036
rect 21506 31034 21562 31036
rect 21586 31034 21642 31036
rect 21666 31034 21722 31036
rect 21426 30982 21472 31034
rect 21472 30982 21482 31034
rect 21506 30982 21536 31034
rect 21536 30982 21548 31034
rect 21548 30982 21562 31034
rect 21586 30982 21600 31034
rect 21600 30982 21612 31034
rect 21612 30982 21642 31034
rect 21666 30982 21676 31034
rect 21676 30982 21722 31034
rect 21426 30980 21482 30982
rect 21506 30980 21562 30982
rect 21586 30980 21642 30982
rect 21666 30980 21722 30982
rect 25520 32666 25576 32668
rect 25600 32666 25656 32668
rect 25680 32666 25736 32668
rect 25760 32666 25816 32668
rect 25520 32614 25566 32666
rect 25566 32614 25576 32666
rect 25600 32614 25630 32666
rect 25630 32614 25642 32666
rect 25642 32614 25656 32666
rect 25680 32614 25694 32666
rect 25694 32614 25706 32666
rect 25706 32614 25736 32666
rect 25760 32614 25770 32666
rect 25770 32614 25816 32666
rect 25520 32612 25576 32614
rect 25600 32612 25656 32614
rect 25680 32612 25736 32614
rect 25760 32612 25816 32614
rect 25520 31578 25576 31580
rect 25600 31578 25656 31580
rect 25680 31578 25736 31580
rect 25760 31578 25816 31580
rect 25520 31526 25566 31578
rect 25566 31526 25576 31578
rect 25600 31526 25630 31578
rect 25630 31526 25642 31578
rect 25642 31526 25656 31578
rect 25680 31526 25694 31578
rect 25694 31526 25706 31578
rect 25706 31526 25736 31578
rect 25760 31526 25770 31578
rect 25770 31526 25816 31578
rect 25520 31524 25576 31526
rect 25600 31524 25656 31526
rect 25680 31524 25736 31526
rect 25760 31524 25816 31526
rect 21426 29946 21482 29948
rect 21506 29946 21562 29948
rect 21586 29946 21642 29948
rect 21666 29946 21722 29948
rect 21426 29894 21472 29946
rect 21472 29894 21482 29946
rect 21506 29894 21536 29946
rect 21536 29894 21548 29946
rect 21548 29894 21562 29946
rect 21586 29894 21600 29946
rect 21600 29894 21612 29946
rect 21612 29894 21642 29946
rect 21666 29894 21676 29946
rect 21676 29894 21722 29946
rect 21426 29892 21482 29894
rect 21506 29892 21562 29894
rect 21586 29892 21642 29894
rect 21666 29892 21722 29894
rect 17332 29402 17388 29404
rect 17412 29402 17468 29404
rect 17492 29402 17548 29404
rect 17572 29402 17628 29404
rect 17332 29350 17378 29402
rect 17378 29350 17388 29402
rect 17412 29350 17442 29402
rect 17442 29350 17454 29402
rect 17454 29350 17468 29402
rect 17492 29350 17506 29402
rect 17506 29350 17518 29402
rect 17518 29350 17548 29402
rect 17572 29350 17582 29402
rect 17582 29350 17628 29402
rect 17332 29348 17388 29350
rect 17412 29348 17468 29350
rect 17492 29348 17548 29350
rect 17572 29348 17628 29350
rect 21426 28858 21482 28860
rect 21506 28858 21562 28860
rect 21586 28858 21642 28860
rect 21666 28858 21722 28860
rect 21426 28806 21472 28858
rect 21472 28806 21482 28858
rect 21506 28806 21536 28858
rect 21536 28806 21548 28858
rect 21548 28806 21562 28858
rect 21586 28806 21600 28858
rect 21600 28806 21612 28858
rect 21612 28806 21642 28858
rect 21666 28806 21676 28858
rect 21676 28806 21722 28858
rect 21426 28804 21482 28806
rect 21506 28804 21562 28806
rect 21586 28804 21642 28806
rect 21666 28804 21722 28806
rect 17332 28314 17388 28316
rect 17412 28314 17468 28316
rect 17492 28314 17548 28316
rect 17572 28314 17628 28316
rect 17332 28262 17378 28314
rect 17378 28262 17388 28314
rect 17412 28262 17442 28314
rect 17442 28262 17454 28314
rect 17454 28262 17468 28314
rect 17492 28262 17506 28314
rect 17506 28262 17518 28314
rect 17518 28262 17548 28314
rect 17572 28262 17582 28314
rect 17582 28262 17628 28314
rect 17332 28260 17388 28262
rect 17412 28260 17468 28262
rect 17492 28260 17548 28262
rect 17572 28260 17628 28262
rect 21426 27770 21482 27772
rect 21506 27770 21562 27772
rect 21586 27770 21642 27772
rect 21666 27770 21722 27772
rect 21426 27718 21472 27770
rect 21472 27718 21482 27770
rect 21506 27718 21536 27770
rect 21536 27718 21548 27770
rect 21548 27718 21562 27770
rect 21586 27718 21600 27770
rect 21600 27718 21612 27770
rect 21612 27718 21642 27770
rect 21666 27718 21676 27770
rect 21676 27718 21722 27770
rect 21426 27716 21482 27718
rect 21506 27716 21562 27718
rect 21586 27716 21642 27718
rect 21666 27716 21722 27718
rect 25520 30490 25576 30492
rect 25600 30490 25656 30492
rect 25680 30490 25736 30492
rect 25760 30490 25816 30492
rect 25520 30438 25566 30490
rect 25566 30438 25576 30490
rect 25600 30438 25630 30490
rect 25630 30438 25642 30490
rect 25642 30438 25656 30490
rect 25680 30438 25694 30490
rect 25694 30438 25706 30490
rect 25706 30438 25736 30490
rect 25760 30438 25770 30490
rect 25770 30438 25816 30490
rect 25520 30436 25576 30438
rect 25600 30436 25656 30438
rect 25680 30436 25736 30438
rect 25760 30436 25816 30438
rect 25520 29402 25576 29404
rect 25600 29402 25656 29404
rect 25680 29402 25736 29404
rect 25760 29402 25816 29404
rect 25520 29350 25566 29402
rect 25566 29350 25576 29402
rect 25600 29350 25630 29402
rect 25630 29350 25642 29402
rect 25642 29350 25656 29402
rect 25680 29350 25694 29402
rect 25694 29350 25706 29402
rect 25706 29350 25736 29402
rect 25760 29350 25770 29402
rect 25770 29350 25816 29402
rect 25520 29348 25576 29350
rect 25600 29348 25656 29350
rect 25680 29348 25736 29350
rect 25760 29348 25816 29350
rect 27434 31320 27490 31376
rect 25520 28314 25576 28316
rect 25600 28314 25656 28316
rect 25680 28314 25736 28316
rect 25760 28314 25816 28316
rect 25520 28262 25566 28314
rect 25566 28262 25576 28314
rect 25600 28262 25630 28314
rect 25630 28262 25642 28314
rect 25642 28262 25656 28314
rect 25680 28262 25694 28314
rect 25694 28262 25706 28314
rect 25706 28262 25736 28314
rect 25760 28262 25770 28314
rect 25770 28262 25816 28314
rect 25520 28260 25576 28262
rect 25600 28260 25656 28262
rect 25680 28260 25736 28262
rect 25760 28260 25816 28262
rect 17332 27226 17388 27228
rect 17412 27226 17468 27228
rect 17492 27226 17548 27228
rect 17572 27226 17628 27228
rect 17332 27174 17378 27226
rect 17378 27174 17388 27226
rect 17412 27174 17442 27226
rect 17442 27174 17454 27226
rect 17454 27174 17468 27226
rect 17492 27174 17506 27226
rect 17506 27174 17518 27226
rect 17518 27174 17548 27226
rect 17572 27174 17582 27226
rect 17582 27174 17628 27226
rect 17332 27172 17388 27174
rect 17412 27172 17468 27174
rect 17492 27172 17548 27174
rect 17572 27172 17628 27174
rect 25520 27226 25576 27228
rect 25600 27226 25656 27228
rect 25680 27226 25736 27228
rect 25760 27226 25816 27228
rect 25520 27174 25566 27226
rect 25566 27174 25576 27226
rect 25600 27174 25630 27226
rect 25630 27174 25642 27226
rect 25642 27174 25656 27226
rect 25680 27174 25694 27226
rect 25694 27174 25706 27226
rect 25706 27174 25736 27226
rect 25760 27174 25770 27226
rect 25770 27174 25816 27226
rect 25520 27172 25576 27174
rect 25600 27172 25656 27174
rect 25680 27172 25736 27174
rect 25760 27172 25816 27174
rect 21426 26682 21482 26684
rect 21506 26682 21562 26684
rect 21586 26682 21642 26684
rect 21666 26682 21722 26684
rect 21426 26630 21472 26682
rect 21472 26630 21482 26682
rect 21506 26630 21536 26682
rect 21536 26630 21548 26682
rect 21548 26630 21562 26682
rect 21586 26630 21600 26682
rect 21600 26630 21612 26682
rect 21612 26630 21642 26682
rect 21666 26630 21676 26682
rect 21676 26630 21722 26682
rect 21426 26628 21482 26630
rect 21506 26628 21562 26630
rect 21586 26628 21642 26630
rect 21666 26628 21722 26630
rect 17332 26138 17388 26140
rect 17412 26138 17468 26140
rect 17492 26138 17548 26140
rect 17572 26138 17628 26140
rect 17332 26086 17378 26138
rect 17378 26086 17388 26138
rect 17412 26086 17442 26138
rect 17442 26086 17454 26138
rect 17454 26086 17468 26138
rect 17492 26086 17506 26138
rect 17506 26086 17518 26138
rect 17518 26086 17548 26138
rect 17572 26086 17582 26138
rect 17582 26086 17628 26138
rect 17332 26084 17388 26086
rect 17412 26084 17468 26086
rect 17492 26084 17548 26086
rect 17572 26084 17628 26086
rect 9144 23962 9200 23964
rect 9224 23962 9280 23964
rect 9304 23962 9360 23964
rect 9384 23962 9440 23964
rect 9144 23910 9190 23962
rect 9190 23910 9200 23962
rect 9224 23910 9254 23962
rect 9254 23910 9266 23962
rect 9266 23910 9280 23962
rect 9304 23910 9318 23962
rect 9318 23910 9330 23962
rect 9330 23910 9360 23962
rect 9384 23910 9394 23962
rect 9394 23910 9440 23962
rect 9144 23908 9200 23910
rect 9224 23908 9280 23910
rect 9304 23908 9360 23910
rect 9384 23908 9440 23910
rect 13238 24506 13294 24508
rect 13318 24506 13374 24508
rect 13398 24506 13454 24508
rect 13478 24506 13534 24508
rect 13238 24454 13284 24506
rect 13284 24454 13294 24506
rect 13318 24454 13348 24506
rect 13348 24454 13360 24506
rect 13360 24454 13374 24506
rect 13398 24454 13412 24506
rect 13412 24454 13424 24506
rect 13424 24454 13454 24506
rect 13478 24454 13488 24506
rect 13488 24454 13534 24506
rect 13238 24452 13294 24454
rect 13318 24452 13374 24454
rect 13398 24452 13454 24454
rect 13478 24452 13534 24454
rect 9144 22874 9200 22876
rect 9224 22874 9280 22876
rect 9304 22874 9360 22876
rect 9384 22874 9440 22876
rect 9144 22822 9190 22874
rect 9190 22822 9200 22874
rect 9224 22822 9254 22874
rect 9254 22822 9266 22874
rect 9266 22822 9280 22874
rect 9304 22822 9318 22874
rect 9318 22822 9330 22874
rect 9330 22822 9360 22874
rect 9384 22822 9394 22874
rect 9394 22822 9440 22874
rect 9144 22820 9200 22822
rect 9224 22820 9280 22822
rect 9304 22820 9360 22822
rect 9384 22820 9440 22822
rect 9144 21786 9200 21788
rect 9224 21786 9280 21788
rect 9304 21786 9360 21788
rect 9384 21786 9440 21788
rect 9144 21734 9190 21786
rect 9190 21734 9200 21786
rect 9224 21734 9254 21786
rect 9254 21734 9266 21786
rect 9266 21734 9280 21786
rect 9304 21734 9318 21786
rect 9318 21734 9330 21786
rect 9330 21734 9360 21786
rect 9384 21734 9394 21786
rect 9394 21734 9440 21786
rect 9144 21732 9200 21734
rect 9224 21732 9280 21734
rect 9304 21732 9360 21734
rect 9384 21732 9440 21734
rect 13238 23418 13294 23420
rect 13318 23418 13374 23420
rect 13398 23418 13454 23420
rect 13478 23418 13534 23420
rect 13238 23366 13284 23418
rect 13284 23366 13294 23418
rect 13318 23366 13348 23418
rect 13348 23366 13360 23418
rect 13360 23366 13374 23418
rect 13398 23366 13412 23418
rect 13412 23366 13424 23418
rect 13424 23366 13454 23418
rect 13478 23366 13488 23418
rect 13488 23366 13534 23418
rect 13238 23364 13294 23366
rect 13318 23364 13374 23366
rect 13398 23364 13454 23366
rect 13478 23364 13534 23366
rect 13238 22330 13294 22332
rect 13318 22330 13374 22332
rect 13398 22330 13454 22332
rect 13478 22330 13534 22332
rect 13238 22278 13284 22330
rect 13284 22278 13294 22330
rect 13318 22278 13348 22330
rect 13348 22278 13360 22330
rect 13360 22278 13374 22330
rect 13398 22278 13412 22330
rect 13412 22278 13424 22330
rect 13424 22278 13454 22330
rect 13478 22278 13488 22330
rect 13488 22278 13534 22330
rect 13238 22276 13294 22278
rect 13318 22276 13374 22278
rect 13398 22276 13454 22278
rect 13478 22276 13534 22278
rect 13238 21242 13294 21244
rect 13318 21242 13374 21244
rect 13398 21242 13454 21244
rect 13478 21242 13534 21244
rect 13238 21190 13284 21242
rect 13284 21190 13294 21242
rect 13318 21190 13348 21242
rect 13348 21190 13360 21242
rect 13360 21190 13374 21242
rect 13398 21190 13412 21242
rect 13412 21190 13424 21242
rect 13424 21190 13454 21242
rect 13478 21190 13488 21242
rect 13488 21190 13534 21242
rect 13238 21188 13294 21190
rect 13318 21188 13374 21190
rect 13398 21188 13454 21190
rect 13478 21188 13534 21190
rect 9144 20698 9200 20700
rect 9224 20698 9280 20700
rect 9304 20698 9360 20700
rect 9384 20698 9440 20700
rect 9144 20646 9190 20698
rect 9190 20646 9200 20698
rect 9224 20646 9254 20698
rect 9254 20646 9266 20698
rect 9266 20646 9280 20698
rect 9304 20646 9318 20698
rect 9318 20646 9330 20698
rect 9330 20646 9360 20698
rect 9384 20646 9394 20698
rect 9394 20646 9440 20698
rect 9144 20644 9200 20646
rect 9224 20644 9280 20646
rect 9304 20644 9360 20646
rect 9384 20644 9440 20646
rect 9144 19610 9200 19612
rect 9224 19610 9280 19612
rect 9304 19610 9360 19612
rect 9384 19610 9440 19612
rect 9144 19558 9190 19610
rect 9190 19558 9200 19610
rect 9224 19558 9254 19610
rect 9254 19558 9266 19610
rect 9266 19558 9280 19610
rect 9304 19558 9318 19610
rect 9318 19558 9330 19610
rect 9330 19558 9360 19610
rect 9384 19558 9394 19610
rect 9394 19558 9440 19610
rect 9144 19556 9200 19558
rect 9224 19556 9280 19558
rect 9304 19556 9360 19558
rect 9384 19556 9440 19558
rect 9144 18522 9200 18524
rect 9224 18522 9280 18524
rect 9304 18522 9360 18524
rect 9384 18522 9440 18524
rect 9144 18470 9190 18522
rect 9190 18470 9200 18522
rect 9224 18470 9254 18522
rect 9254 18470 9266 18522
rect 9266 18470 9280 18522
rect 9304 18470 9318 18522
rect 9318 18470 9330 18522
rect 9330 18470 9360 18522
rect 9384 18470 9394 18522
rect 9394 18470 9440 18522
rect 9144 18468 9200 18470
rect 9224 18468 9280 18470
rect 9304 18468 9360 18470
rect 9384 18468 9440 18470
rect 5050 17978 5106 17980
rect 5130 17978 5186 17980
rect 5210 17978 5266 17980
rect 5290 17978 5346 17980
rect 5050 17926 5096 17978
rect 5096 17926 5106 17978
rect 5130 17926 5160 17978
rect 5160 17926 5172 17978
rect 5172 17926 5186 17978
rect 5210 17926 5224 17978
rect 5224 17926 5236 17978
rect 5236 17926 5266 17978
rect 5290 17926 5300 17978
rect 5300 17926 5346 17978
rect 5050 17924 5106 17926
rect 5130 17924 5186 17926
rect 5210 17924 5266 17926
rect 5290 17924 5346 17926
rect 13238 20154 13294 20156
rect 13318 20154 13374 20156
rect 13398 20154 13454 20156
rect 13478 20154 13534 20156
rect 13238 20102 13284 20154
rect 13284 20102 13294 20154
rect 13318 20102 13348 20154
rect 13348 20102 13360 20154
rect 13360 20102 13374 20154
rect 13398 20102 13412 20154
rect 13412 20102 13424 20154
rect 13424 20102 13454 20154
rect 13478 20102 13488 20154
rect 13488 20102 13534 20154
rect 13238 20100 13294 20102
rect 13318 20100 13374 20102
rect 13398 20100 13454 20102
rect 13478 20100 13534 20102
rect 13238 19066 13294 19068
rect 13318 19066 13374 19068
rect 13398 19066 13454 19068
rect 13478 19066 13534 19068
rect 13238 19014 13284 19066
rect 13284 19014 13294 19066
rect 13318 19014 13348 19066
rect 13348 19014 13360 19066
rect 13360 19014 13374 19066
rect 13398 19014 13412 19066
rect 13412 19014 13424 19066
rect 13424 19014 13454 19066
rect 13478 19014 13488 19066
rect 13488 19014 13534 19066
rect 13238 19012 13294 19014
rect 13318 19012 13374 19014
rect 13398 19012 13454 19014
rect 13478 19012 13534 19014
rect 13238 17978 13294 17980
rect 13318 17978 13374 17980
rect 13398 17978 13454 17980
rect 13478 17978 13534 17980
rect 13238 17926 13284 17978
rect 13284 17926 13294 17978
rect 13318 17926 13348 17978
rect 13348 17926 13360 17978
rect 13360 17926 13374 17978
rect 13398 17926 13412 17978
rect 13412 17926 13424 17978
rect 13424 17926 13454 17978
rect 13478 17926 13488 17978
rect 13488 17926 13534 17978
rect 13238 17924 13294 17926
rect 13318 17924 13374 17926
rect 13398 17924 13454 17926
rect 13478 17924 13534 17926
rect 9144 17434 9200 17436
rect 9224 17434 9280 17436
rect 9304 17434 9360 17436
rect 9384 17434 9440 17436
rect 9144 17382 9190 17434
rect 9190 17382 9200 17434
rect 9224 17382 9254 17434
rect 9254 17382 9266 17434
rect 9266 17382 9280 17434
rect 9304 17382 9318 17434
rect 9318 17382 9330 17434
rect 9330 17382 9360 17434
rect 9384 17382 9394 17434
rect 9394 17382 9440 17434
rect 9144 17380 9200 17382
rect 9224 17380 9280 17382
rect 9304 17380 9360 17382
rect 9384 17380 9440 17382
rect 5050 16890 5106 16892
rect 5130 16890 5186 16892
rect 5210 16890 5266 16892
rect 5290 16890 5346 16892
rect 5050 16838 5096 16890
rect 5096 16838 5106 16890
rect 5130 16838 5160 16890
rect 5160 16838 5172 16890
rect 5172 16838 5186 16890
rect 5210 16838 5224 16890
rect 5224 16838 5236 16890
rect 5236 16838 5266 16890
rect 5290 16838 5300 16890
rect 5300 16838 5346 16890
rect 5050 16836 5106 16838
rect 5130 16836 5186 16838
rect 5210 16836 5266 16838
rect 5290 16836 5346 16838
rect 5050 15802 5106 15804
rect 5130 15802 5186 15804
rect 5210 15802 5266 15804
rect 5290 15802 5346 15804
rect 5050 15750 5096 15802
rect 5096 15750 5106 15802
rect 5130 15750 5160 15802
rect 5160 15750 5172 15802
rect 5172 15750 5186 15802
rect 5210 15750 5224 15802
rect 5224 15750 5236 15802
rect 5236 15750 5266 15802
rect 5290 15750 5300 15802
rect 5300 15750 5346 15802
rect 5050 15748 5106 15750
rect 5130 15748 5186 15750
rect 5210 15748 5266 15750
rect 5290 15748 5346 15750
rect 9144 16346 9200 16348
rect 9224 16346 9280 16348
rect 9304 16346 9360 16348
rect 9384 16346 9440 16348
rect 9144 16294 9190 16346
rect 9190 16294 9200 16346
rect 9224 16294 9254 16346
rect 9254 16294 9266 16346
rect 9266 16294 9280 16346
rect 9304 16294 9318 16346
rect 9318 16294 9330 16346
rect 9330 16294 9360 16346
rect 9384 16294 9394 16346
rect 9394 16294 9440 16346
rect 9144 16292 9200 16294
rect 9224 16292 9280 16294
rect 9304 16292 9360 16294
rect 9384 16292 9440 16294
rect 9144 15258 9200 15260
rect 9224 15258 9280 15260
rect 9304 15258 9360 15260
rect 9384 15258 9440 15260
rect 9144 15206 9190 15258
rect 9190 15206 9200 15258
rect 9224 15206 9254 15258
rect 9254 15206 9266 15258
rect 9266 15206 9280 15258
rect 9304 15206 9318 15258
rect 9318 15206 9330 15258
rect 9330 15206 9360 15258
rect 9384 15206 9394 15258
rect 9394 15206 9440 15258
rect 9144 15204 9200 15206
rect 9224 15204 9280 15206
rect 9304 15204 9360 15206
rect 9384 15204 9440 15206
rect 5050 14714 5106 14716
rect 5130 14714 5186 14716
rect 5210 14714 5266 14716
rect 5290 14714 5346 14716
rect 5050 14662 5096 14714
rect 5096 14662 5106 14714
rect 5130 14662 5160 14714
rect 5160 14662 5172 14714
rect 5172 14662 5186 14714
rect 5210 14662 5224 14714
rect 5224 14662 5236 14714
rect 5236 14662 5266 14714
rect 5290 14662 5300 14714
rect 5300 14662 5346 14714
rect 5050 14660 5106 14662
rect 5130 14660 5186 14662
rect 5210 14660 5266 14662
rect 5290 14660 5346 14662
rect 5050 13626 5106 13628
rect 5130 13626 5186 13628
rect 5210 13626 5266 13628
rect 5290 13626 5346 13628
rect 5050 13574 5096 13626
rect 5096 13574 5106 13626
rect 5130 13574 5160 13626
rect 5160 13574 5172 13626
rect 5172 13574 5186 13626
rect 5210 13574 5224 13626
rect 5224 13574 5236 13626
rect 5236 13574 5266 13626
rect 5290 13574 5300 13626
rect 5300 13574 5346 13626
rect 5050 13572 5106 13574
rect 5130 13572 5186 13574
rect 5210 13572 5266 13574
rect 5290 13572 5346 13574
rect 5050 12538 5106 12540
rect 5130 12538 5186 12540
rect 5210 12538 5266 12540
rect 5290 12538 5346 12540
rect 5050 12486 5096 12538
rect 5096 12486 5106 12538
rect 5130 12486 5160 12538
rect 5160 12486 5172 12538
rect 5172 12486 5186 12538
rect 5210 12486 5224 12538
rect 5224 12486 5236 12538
rect 5236 12486 5266 12538
rect 5290 12486 5300 12538
rect 5300 12486 5346 12538
rect 5050 12484 5106 12486
rect 5130 12484 5186 12486
rect 5210 12484 5266 12486
rect 5290 12484 5346 12486
rect 9144 14170 9200 14172
rect 9224 14170 9280 14172
rect 9304 14170 9360 14172
rect 9384 14170 9440 14172
rect 9144 14118 9190 14170
rect 9190 14118 9200 14170
rect 9224 14118 9254 14170
rect 9254 14118 9266 14170
rect 9266 14118 9280 14170
rect 9304 14118 9318 14170
rect 9318 14118 9330 14170
rect 9330 14118 9360 14170
rect 9384 14118 9394 14170
rect 9394 14118 9440 14170
rect 9144 14116 9200 14118
rect 9224 14116 9280 14118
rect 9304 14116 9360 14118
rect 9384 14116 9440 14118
rect 9144 13082 9200 13084
rect 9224 13082 9280 13084
rect 9304 13082 9360 13084
rect 9384 13082 9440 13084
rect 9144 13030 9190 13082
rect 9190 13030 9200 13082
rect 9224 13030 9254 13082
rect 9254 13030 9266 13082
rect 9266 13030 9280 13082
rect 9304 13030 9318 13082
rect 9318 13030 9330 13082
rect 9330 13030 9360 13082
rect 9384 13030 9394 13082
rect 9394 13030 9440 13082
rect 9144 13028 9200 13030
rect 9224 13028 9280 13030
rect 9304 13028 9360 13030
rect 9384 13028 9440 13030
rect 5050 11450 5106 11452
rect 5130 11450 5186 11452
rect 5210 11450 5266 11452
rect 5290 11450 5346 11452
rect 5050 11398 5096 11450
rect 5096 11398 5106 11450
rect 5130 11398 5160 11450
rect 5160 11398 5172 11450
rect 5172 11398 5186 11450
rect 5210 11398 5224 11450
rect 5224 11398 5236 11450
rect 5236 11398 5266 11450
rect 5290 11398 5300 11450
rect 5300 11398 5346 11450
rect 5050 11396 5106 11398
rect 5130 11396 5186 11398
rect 5210 11396 5266 11398
rect 5290 11396 5346 11398
rect 5050 10362 5106 10364
rect 5130 10362 5186 10364
rect 5210 10362 5266 10364
rect 5290 10362 5346 10364
rect 5050 10310 5096 10362
rect 5096 10310 5106 10362
rect 5130 10310 5160 10362
rect 5160 10310 5172 10362
rect 5172 10310 5186 10362
rect 5210 10310 5224 10362
rect 5224 10310 5236 10362
rect 5236 10310 5266 10362
rect 5290 10310 5300 10362
rect 5300 10310 5346 10362
rect 5050 10308 5106 10310
rect 5130 10308 5186 10310
rect 5210 10308 5266 10310
rect 5290 10308 5346 10310
rect 5050 9274 5106 9276
rect 5130 9274 5186 9276
rect 5210 9274 5266 9276
rect 5290 9274 5346 9276
rect 5050 9222 5096 9274
rect 5096 9222 5106 9274
rect 5130 9222 5160 9274
rect 5160 9222 5172 9274
rect 5172 9222 5186 9274
rect 5210 9222 5224 9274
rect 5224 9222 5236 9274
rect 5236 9222 5266 9274
rect 5290 9222 5300 9274
rect 5300 9222 5346 9274
rect 5050 9220 5106 9222
rect 5130 9220 5186 9222
rect 5210 9220 5266 9222
rect 5290 9220 5346 9222
rect 5050 8186 5106 8188
rect 5130 8186 5186 8188
rect 5210 8186 5266 8188
rect 5290 8186 5346 8188
rect 5050 8134 5096 8186
rect 5096 8134 5106 8186
rect 5130 8134 5160 8186
rect 5160 8134 5172 8186
rect 5172 8134 5186 8186
rect 5210 8134 5224 8186
rect 5224 8134 5236 8186
rect 5236 8134 5266 8186
rect 5290 8134 5300 8186
rect 5300 8134 5346 8186
rect 5050 8132 5106 8134
rect 5130 8132 5186 8134
rect 5210 8132 5266 8134
rect 5290 8132 5346 8134
rect 5050 7098 5106 7100
rect 5130 7098 5186 7100
rect 5210 7098 5266 7100
rect 5290 7098 5346 7100
rect 5050 7046 5096 7098
rect 5096 7046 5106 7098
rect 5130 7046 5160 7098
rect 5160 7046 5172 7098
rect 5172 7046 5186 7098
rect 5210 7046 5224 7098
rect 5224 7046 5236 7098
rect 5236 7046 5266 7098
rect 5290 7046 5300 7098
rect 5300 7046 5346 7098
rect 5050 7044 5106 7046
rect 5130 7044 5186 7046
rect 5210 7044 5266 7046
rect 5290 7044 5346 7046
rect 5050 6010 5106 6012
rect 5130 6010 5186 6012
rect 5210 6010 5266 6012
rect 5290 6010 5346 6012
rect 5050 5958 5096 6010
rect 5096 5958 5106 6010
rect 5130 5958 5160 6010
rect 5160 5958 5172 6010
rect 5172 5958 5186 6010
rect 5210 5958 5224 6010
rect 5224 5958 5236 6010
rect 5236 5958 5266 6010
rect 5290 5958 5300 6010
rect 5300 5958 5346 6010
rect 5050 5956 5106 5958
rect 5130 5956 5186 5958
rect 5210 5956 5266 5958
rect 5290 5956 5346 5958
rect 5050 4922 5106 4924
rect 5130 4922 5186 4924
rect 5210 4922 5266 4924
rect 5290 4922 5346 4924
rect 5050 4870 5096 4922
rect 5096 4870 5106 4922
rect 5130 4870 5160 4922
rect 5160 4870 5172 4922
rect 5172 4870 5186 4922
rect 5210 4870 5224 4922
rect 5224 4870 5236 4922
rect 5236 4870 5266 4922
rect 5290 4870 5300 4922
rect 5300 4870 5346 4922
rect 5050 4868 5106 4870
rect 5130 4868 5186 4870
rect 5210 4868 5266 4870
rect 5290 4868 5346 4870
rect 5050 3834 5106 3836
rect 5130 3834 5186 3836
rect 5210 3834 5266 3836
rect 5290 3834 5346 3836
rect 5050 3782 5096 3834
rect 5096 3782 5106 3834
rect 5130 3782 5160 3834
rect 5160 3782 5172 3834
rect 5172 3782 5186 3834
rect 5210 3782 5224 3834
rect 5224 3782 5236 3834
rect 5236 3782 5266 3834
rect 5290 3782 5300 3834
rect 5300 3782 5346 3834
rect 5050 3780 5106 3782
rect 5130 3780 5186 3782
rect 5210 3780 5266 3782
rect 5290 3780 5346 3782
rect 1582 2760 1638 2816
rect 5050 2746 5106 2748
rect 5130 2746 5186 2748
rect 5210 2746 5266 2748
rect 5290 2746 5346 2748
rect 5050 2694 5096 2746
rect 5096 2694 5106 2746
rect 5130 2694 5160 2746
rect 5160 2694 5172 2746
rect 5172 2694 5186 2746
rect 5210 2694 5224 2746
rect 5224 2694 5236 2746
rect 5236 2694 5266 2746
rect 5290 2694 5300 2746
rect 5300 2694 5346 2746
rect 5050 2692 5106 2694
rect 5130 2692 5186 2694
rect 5210 2692 5266 2694
rect 5290 2692 5346 2694
rect 9144 11994 9200 11996
rect 9224 11994 9280 11996
rect 9304 11994 9360 11996
rect 9384 11994 9440 11996
rect 9144 11942 9190 11994
rect 9190 11942 9200 11994
rect 9224 11942 9254 11994
rect 9254 11942 9266 11994
rect 9266 11942 9280 11994
rect 9304 11942 9318 11994
rect 9318 11942 9330 11994
rect 9330 11942 9360 11994
rect 9384 11942 9394 11994
rect 9394 11942 9440 11994
rect 9144 11940 9200 11942
rect 9224 11940 9280 11942
rect 9304 11940 9360 11942
rect 9384 11940 9440 11942
rect 9144 10906 9200 10908
rect 9224 10906 9280 10908
rect 9304 10906 9360 10908
rect 9384 10906 9440 10908
rect 9144 10854 9190 10906
rect 9190 10854 9200 10906
rect 9224 10854 9254 10906
rect 9254 10854 9266 10906
rect 9266 10854 9280 10906
rect 9304 10854 9318 10906
rect 9318 10854 9330 10906
rect 9330 10854 9360 10906
rect 9384 10854 9394 10906
rect 9394 10854 9440 10906
rect 9144 10852 9200 10854
rect 9224 10852 9280 10854
rect 9304 10852 9360 10854
rect 9384 10852 9440 10854
rect 9144 9818 9200 9820
rect 9224 9818 9280 9820
rect 9304 9818 9360 9820
rect 9384 9818 9440 9820
rect 9144 9766 9190 9818
rect 9190 9766 9200 9818
rect 9224 9766 9254 9818
rect 9254 9766 9266 9818
rect 9266 9766 9280 9818
rect 9304 9766 9318 9818
rect 9318 9766 9330 9818
rect 9330 9766 9360 9818
rect 9384 9766 9394 9818
rect 9394 9766 9440 9818
rect 9144 9764 9200 9766
rect 9224 9764 9280 9766
rect 9304 9764 9360 9766
rect 9384 9764 9440 9766
rect 13238 16890 13294 16892
rect 13318 16890 13374 16892
rect 13398 16890 13454 16892
rect 13478 16890 13534 16892
rect 13238 16838 13284 16890
rect 13284 16838 13294 16890
rect 13318 16838 13348 16890
rect 13348 16838 13360 16890
rect 13360 16838 13374 16890
rect 13398 16838 13412 16890
rect 13412 16838 13424 16890
rect 13424 16838 13454 16890
rect 13478 16838 13488 16890
rect 13488 16838 13534 16890
rect 13238 16836 13294 16838
rect 13318 16836 13374 16838
rect 13398 16836 13454 16838
rect 13478 16836 13534 16838
rect 13238 15802 13294 15804
rect 13318 15802 13374 15804
rect 13398 15802 13454 15804
rect 13478 15802 13534 15804
rect 13238 15750 13284 15802
rect 13284 15750 13294 15802
rect 13318 15750 13348 15802
rect 13348 15750 13360 15802
rect 13360 15750 13374 15802
rect 13398 15750 13412 15802
rect 13412 15750 13424 15802
rect 13424 15750 13454 15802
rect 13478 15750 13488 15802
rect 13488 15750 13534 15802
rect 13238 15748 13294 15750
rect 13318 15748 13374 15750
rect 13398 15748 13454 15750
rect 13478 15748 13534 15750
rect 13238 14714 13294 14716
rect 13318 14714 13374 14716
rect 13398 14714 13454 14716
rect 13478 14714 13534 14716
rect 13238 14662 13284 14714
rect 13284 14662 13294 14714
rect 13318 14662 13348 14714
rect 13348 14662 13360 14714
rect 13360 14662 13374 14714
rect 13398 14662 13412 14714
rect 13412 14662 13424 14714
rect 13424 14662 13454 14714
rect 13478 14662 13488 14714
rect 13488 14662 13534 14714
rect 13238 14660 13294 14662
rect 13318 14660 13374 14662
rect 13398 14660 13454 14662
rect 13478 14660 13534 14662
rect 17332 25050 17388 25052
rect 17412 25050 17468 25052
rect 17492 25050 17548 25052
rect 17572 25050 17628 25052
rect 17332 24998 17378 25050
rect 17378 24998 17388 25050
rect 17412 24998 17442 25050
rect 17442 24998 17454 25050
rect 17454 24998 17468 25050
rect 17492 24998 17506 25050
rect 17506 24998 17518 25050
rect 17518 24998 17548 25050
rect 17572 24998 17582 25050
rect 17582 24998 17628 25050
rect 17332 24996 17388 24998
rect 17412 24996 17468 24998
rect 17492 24996 17548 24998
rect 17572 24996 17628 24998
rect 17332 23962 17388 23964
rect 17412 23962 17468 23964
rect 17492 23962 17548 23964
rect 17572 23962 17628 23964
rect 17332 23910 17378 23962
rect 17378 23910 17388 23962
rect 17412 23910 17442 23962
rect 17442 23910 17454 23962
rect 17454 23910 17468 23962
rect 17492 23910 17506 23962
rect 17506 23910 17518 23962
rect 17518 23910 17548 23962
rect 17572 23910 17582 23962
rect 17582 23910 17628 23962
rect 17332 23908 17388 23910
rect 17412 23908 17468 23910
rect 17492 23908 17548 23910
rect 17572 23908 17628 23910
rect 25520 26138 25576 26140
rect 25600 26138 25656 26140
rect 25680 26138 25736 26140
rect 25760 26138 25816 26140
rect 25520 26086 25566 26138
rect 25566 26086 25576 26138
rect 25600 26086 25630 26138
rect 25630 26086 25642 26138
rect 25642 26086 25656 26138
rect 25680 26086 25694 26138
rect 25694 26086 25706 26138
rect 25706 26086 25736 26138
rect 25760 26086 25770 26138
rect 25770 26086 25816 26138
rect 25520 26084 25576 26086
rect 25600 26084 25656 26086
rect 25680 26084 25736 26086
rect 25760 26084 25816 26086
rect 21426 25594 21482 25596
rect 21506 25594 21562 25596
rect 21586 25594 21642 25596
rect 21666 25594 21722 25596
rect 21426 25542 21472 25594
rect 21472 25542 21482 25594
rect 21506 25542 21536 25594
rect 21536 25542 21548 25594
rect 21548 25542 21562 25594
rect 21586 25542 21600 25594
rect 21600 25542 21612 25594
rect 21612 25542 21642 25594
rect 21666 25542 21676 25594
rect 21676 25542 21722 25594
rect 21426 25540 21482 25542
rect 21506 25540 21562 25542
rect 21586 25540 21642 25542
rect 21666 25540 21722 25542
rect 25520 25050 25576 25052
rect 25600 25050 25656 25052
rect 25680 25050 25736 25052
rect 25760 25050 25816 25052
rect 25520 24998 25566 25050
rect 25566 24998 25576 25050
rect 25600 24998 25630 25050
rect 25630 24998 25642 25050
rect 25642 24998 25656 25050
rect 25680 24998 25694 25050
rect 25694 24998 25706 25050
rect 25706 24998 25736 25050
rect 25760 24998 25770 25050
rect 25770 24998 25816 25050
rect 25520 24996 25576 24998
rect 25600 24996 25656 24998
rect 25680 24996 25736 24998
rect 25760 24996 25816 24998
rect 21426 24506 21482 24508
rect 21506 24506 21562 24508
rect 21586 24506 21642 24508
rect 21666 24506 21722 24508
rect 21426 24454 21472 24506
rect 21472 24454 21482 24506
rect 21506 24454 21536 24506
rect 21536 24454 21548 24506
rect 21548 24454 21562 24506
rect 21586 24454 21600 24506
rect 21600 24454 21612 24506
rect 21612 24454 21642 24506
rect 21666 24454 21676 24506
rect 21676 24454 21722 24506
rect 21426 24452 21482 24454
rect 21506 24452 21562 24454
rect 21586 24452 21642 24454
rect 21666 24452 21722 24454
rect 25520 23962 25576 23964
rect 25600 23962 25656 23964
rect 25680 23962 25736 23964
rect 25760 23962 25816 23964
rect 25520 23910 25566 23962
rect 25566 23910 25576 23962
rect 25600 23910 25630 23962
rect 25630 23910 25642 23962
rect 25642 23910 25656 23962
rect 25680 23910 25694 23962
rect 25694 23910 25706 23962
rect 25706 23910 25736 23962
rect 25760 23910 25770 23962
rect 25770 23910 25816 23962
rect 25520 23908 25576 23910
rect 25600 23908 25656 23910
rect 25680 23908 25736 23910
rect 25760 23908 25816 23910
rect 21426 23418 21482 23420
rect 21506 23418 21562 23420
rect 21586 23418 21642 23420
rect 21666 23418 21722 23420
rect 21426 23366 21472 23418
rect 21472 23366 21482 23418
rect 21506 23366 21536 23418
rect 21536 23366 21548 23418
rect 21548 23366 21562 23418
rect 21586 23366 21600 23418
rect 21600 23366 21612 23418
rect 21612 23366 21642 23418
rect 21666 23366 21676 23418
rect 21676 23366 21722 23418
rect 21426 23364 21482 23366
rect 21506 23364 21562 23366
rect 21586 23364 21642 23366
rect 21666 23364 21722 23366
rect 17332 22874 17388 22876
rect 17412 22874 17468 22876
rect 17492 22874 17548 22876
rect 17572 22874 17628 22876
rect 17332 22822 17378 22874
rect 17378 22822 17388 22874
rect 17412 22822 17442 22874
rect 17442 22822 17454 22874
rect 17454 22822 17468 22874
rect 17492 22822 17506 22874
rect 17506 22822 17518 22874
rect 17518 22822 17548 22874
rect 17572 22822 17582 22874
rect 17582 22822 17628 22874
rect 17332 22820 17388 22822
rect 17412 22820 17468 22822
rect 17492 22820 17548 22822
rect 17572 22820 17628 22822
rect 21426 22330 21482 22332
rect 21506 22330 21562 22332
rect 21586 22330 21642 22332
rect 21666 22330 21722 22332
rect 21426 22278 21472 22330
rect 21472 22278 21482 22330
rect 21506 22278 21536 22330
rect 21536 22278 21548 22330
rect 21548 22278 21562 22330
rect 21586 22278 21600 22330
rect 21600 22278 21612 22330
rect 21612 22278 21642 22330
rect 21666 22278 21676 22330
rect 21676 22278 21722 22330
rect 21426 22276 21482 22278
rect 21506 22276 21562 22278
rect 21586 22276 21642 22278
rect 21666 22276 21722 22278
rect 17332 21786 17388 21788
rect 17412 21786 17468 21788
rect 17492 21786 17548 21788
rect 17572 21786 17628 21788
rect 17332 21734 17378 21786
rect 17378 21734 17388 21786
rect 17412 21734 17442 21786
rect 17442 21734 17454 21786
rect 17454 21734 17468 21786
rect 17492 21734 17506 21786
rect 17506 21734 17518 21786
rect 17518 21734 17548 21786
rect 17572 21734 17582 21786
rect 17582 21734 17628 21786
rect 17332 21732 17388 21734
rect 17412 21732 17468 21734
rect 17492 21732 17548 21734
rect 17572 21732 17628 21734
rect 21426 21242 21482 21244
rect 21506 21242 21562 21244
rect 21586 21242 21642 21244
rect 21666 21242 21722 21244
rect 21426 21190 21472 21242
rect 21472 21190 21482 21242
rect 21506 21190 21536 21242
rect 21536 21190 21548 21242
rect 21548 21190 21562 21242
rect 21586 21190 21600 21242
rect 21600 21190 21612 21242
rect 21612 21190 21642 21242
rect 21666 21190 21676 21242
rect 21676 21190 21722 21242
rect 21426 21188 21482 21190
rect 21506 21188 21562 21190
rect 21586 21188 21642 21190
rect 21666 21188 21722 21190
rect 29614 32122 29670 32124
rect 29694 32122 29750 32124
rect 29774 32122 29830 32124
rect 29854 32122 29910 32124
rect 29614 32070 29660 32122
rect 29660 32070 29670 32122
rect 29694 32070 29724 32122
rect 29724 32070 29736 32122
rect 29736 32070 29750 32122
rect 29774 32070 29788 32122
rect 29788 32070 29800 32122
rect 29800 32070 29830 32122
rect 29854 32070 29864 32122
rect 29864 32070 29910 32122
rect 29614 32068 29670 32070
rect 29694 32068 29750 32070
rect 29774 32068 29830 32070
rect 29854 32068 29910 32070
rect 29614 31034 29670 31036
rect 29694 31034 29750 31036
rect 29774 31034 29830 31036
rect 29854 31034 29910 31036
rect 29614 30982 29660 31034
rect 29660 30982 29670 31034
rect 29694 30982 29724 31034
rect 29724 30982 29736 31034
rect 29736 30982 29750 31034
rect 29774 30982 29788 31034
rect 29788 30982 29800 31034
rect 29800 30982 29830 31034
rect 29854 30982 29864 31034
rect 29864 30982 29910 31034
rect 29614 30980 29670 30982
rect 29694 30980 29750 30982
rect 29774 30980 29830 30982
rect 29854 30980 29910 30982
rect 29614 29946 29670 29948
rect 29694 29946 29750 29948
rect 29774 29946 29830 29948
rect 29854 29946 29910 29948
rect 29614 29894 29660 29946
rect 29660 29894 29670 29946
rect 29694 29894 29724 29946
rect 29724 29894 29736 29946
rect 29736 29894 29750 29946
rect 29774 29894 29788 29946
rect 29788 29894 29800 29946
rect 29800 29894 29830 29946
rect 29854 29894 29864 29946
rect 29864 29894 29910 29946
rect 29614 29892 29670 29894
rect 29694 29892 29750 29894
rect 29774 29892 29830 29894
rect 29854 29892 29910 29894
rect 29614 28858 29670 28860
rect 29694 28858 29750 28860
rect 29774 28858 29830 28860
rect 29854 28858 29910 28860
rect 29614 28806 29660 28858
rect 29660 28806 29670 28858
rect 29694 28806 29724 28858
rect 29724 28806 29736 28858
rect 29736 28806 29750 28858
rect 29774 28806 29788 28858
rect 29788 28806 29800 28858
rect 29800 28806 29830 28858
rect 29854 28806 29864 28858
rect 29864 28806 29910 28858
rect 29614 28804 29670 28806
rect 29694 28804 29750 28806
rect 29774 28804 29830 28806
rect 29854 28804 29910 28806
rect 29614 27770 29670 27772
rect 29694 27770 29750 27772
rect 29774 27770 29830 27772
rect 29854 27770 29910 27772
rect 29614 27718 29660 27770
rect 29660 27718 29670 27770
rect 29694 27718 29724 27770
rect 29724 27718 29736 27770
rect 29736 27718 29750 27770
rect 29774 27718 29788 27770
rect 29788 27718 29800 27770
rect 29800 27718 29830 27770
rect 29854 27718 29864 27770
rect 29864 27718 29910 27770
rect 29614 27716 29670 27718
rect 29694 27716 29750 27718
rect 29774 27716 29830 27718
rect 29854 27716 29910 27718
rect 31298 32952 31354 33008
rect 31482 28872 31538 28928
rect 31482 27512 31538 27568
rect 29614 26682 29670 26684
rect 29694 26682 29750 26684
rect 29774 26682 29830 26684
rect 29854 26682 29910 26684
rect 29614 26630 29660 26682
rect 29660 26630 29670 26682
rect 29694 26630 29724 26682
rect 29724 26630 29736 26682
rect 29736 26630 29750 26682
rect 29774 26630 29788 26682
rect 29788 26630 29800 26682
rect 29800 26630 29830 26682
rect 29854 26630 29864 26682
rect 29864 26630 29910 26682
rect 29614 26628 29670 26630
rect 29694 26628 29750 26630
rect 29774 26628 29830 26630
rect 29854 26628 29910 26630
rect 29614 25594 29670 25596
rect 29694 25594 29750 25596
rect 29774 25594 29830 25596
rect 29854 25594 29910 25596
rect 29614 25542 29660 25594
rect 29660 25542 29670 25594
rect 29694 25542 29724 25594
rect 29724 25542 29736 25594
rect 29736 25542 29750 25594
rect 29774 25542 29788 25594
rect 29788 25542 29800 25594
rect 29800 25542 29830 25594
rect 29854 25542 29864 25594
rect 29864 25542 29910 25594
rect 29614 25540 29670 25542
rect 29694 25540 29750 25542
rect 29774 25540 29830 25542
rect 29854 25540 29910 25542
rect 25520 22874 25576 22876
rect 25600 22874 25656 22876
rect 25680 22874 25736 22876
rect 25760 22874 25816 22876
rect 25520 22822 25566 22874
rect 25566 22822 25576 22874
rect 25600 22822 25630 22874
rect 25630 22822 25642 22874
rect 25642 22822 25656 22874
rect 25680 22822 25694 22874
rect 25694 22822 25706 22874
rect 25706 22822 25736 22874
rect 25760 22822 25770 22874
rect 25770 22822 25816 22874
rect 25520 22820 25576 22822
rect 25600 22820 25656 22822
rect 25680 22820 25736 22822
rect 25760 22820 25816 22822
rect 25520 21786 25576 21788
rect 25600 21786 25656 21788
rect 25680 21786 25736 21788
rect 25760 21786 25816 21788
rect 25520 21734 25566 21786
rect 25566 21734 25576 21786
rect 25600 21734 25630 21786
rect 25630 21734 25642 21786
rect 25642 21734 25656 21786
rect 25680 21734 25694 21786
rect 25694 21734 25706 21786
rect 25706 21734 25736 21786
rect 25760 21734 25770 21786
rect 25770 21734 25816 21786
rect 25520 21732 25576 21734
rect 25600 21732 25656 21734
rect 25680 21732 25736 21734
rect 25760 21732 25816 21734
rect 17332 20698 17388 20700
rect 17412 20698 17468 20700
rect 17492 20698 17548 20700
rect 17572 20698 17628 20700
rect 17332 20646 17378 20698
rect 17378 20646 17388 20698
rect 17412 20646 17442 20698
rect 17442 20646 17454 20698
rect 17454 20646 17468 20698
rect 17492 20646 17506 20698
rect 17506 20646 17518 20698
rect 17518 20646 17548 20698
rect 17572 20646 17582 20698
rect 17582 20646 17628 20698
rect 17332 20644 17388 20646
rect 17412 20644 17468 20646
rect 17492 20644 17548 20646
rect 17572 20644 17628 20646
rect 21426 20154 21482 20156
rect 21506 20154 21562 20156
rect 21586 20154 21642 20156
rect 21666 20154 21722 20156
rect 21426 20102 21472 20154
rect 21472 20102 21482 20154
rect 21506 20102 21536 20154
rect 21536 20102 21548 20154
rect 21548 20102 21562 20154
rect 21586 20102 21600 20154
rect 21600 20102 21612 20154
rect 21612 20102 21642 20154
rect 21666 20102 21676 20154
rect 21676 20102 21722 20154
rect 21426 20100 21482 20102
rect 21506 20100 21562 20102
rect 21586 20100 21642 20102
rect 21666 20100 21722 20102
rect 17332 19610 17388 19612
rect 17412 19610 17468 19612
rect 17492 19610 17548 19612
rect 17572 19610 17628 19612
rect 17332 19558 17378 19610
rect 17378 19558 17388 19610
rect 17412 19558 17442 19610
rect 17442 19558 17454 19610
rect 17454 19558 17468 19610
rect 17492 19558 17506 19610
rect 17506 19558 17518 19610
rect 17518 19558 17548 19610
rect 17572 19558 17582 19610
rect 17582 19558 17628 19610
rect 17332 19556 17388 19558
rect 17412 19556 17468 19558
rect 17492 19556 17548 19558
rect 17572 19556 17628 19558
rect 21426 19066 21482 19068
rect 21506 19066 21562 19068
rect 21586 19066 21642 19068
rect 21666 19066 21722 19068
rect 21426 19014 21472 19066
rect 21472 19014 21482 19066
rect 21506 19014 21536 19066
rect 21536 19014 21548 19066
rect 21548 19014 21562 19066
rect 21586 19014 21600 19066
rect 21600 19014 21612 19066
rect 21612 19014 21642 19066
rect 21666 19014 21676 19066
rect 21676 19014 21722 19066
rect 21426 19012 21482 19014
rect 21506 19012 21562 19014
rect 21586 19012 21642 19014
rect 21666 19012 21722 19014
rect 17332 18522 17388 18524
rect 17412 18522 17468 18524
rect 17492 18522 17548 18524
rect 17572 18522 17628 18524
rect 17332 18470 17378 18522
rect 17378 18470 17388 18522
rect 17412 18470 17442 18522
rect 17442 18470 17454 18522
rect 17454 18470 17468 18522
rect 17492 18470 17506 18522
rect 17506 18470 17518 18522
rect 17518 18470 17548 18522
rect 17572 18470 17582 18522
rect 17582 18470 17628 18522
rect 17332 18468 17388 18470
rect 17412 18468 17468 18470
rect 17492 18468 17548 18470
rect 17572 18468 17628 18470
rect 17332 17434 17388 17436
rect 17412 17434 17468 17436
rect 17492 17434 17548 17436
rect 17572 17434 17628 17436
rect 17332 17382 17378 17434
rect 17378 17382 17388 17434
rect 17412 17382 17442 17434
rect 17442 17382 17454 17434
rect 17454 17382 17468 17434
rect 17492 17382 17506 17434
rect 17506 17382 17518 17434
rect 17518 17382 17548 17434
rect 17572 17382 17582 17434
rect 17582 17382 17628 17434
rect 17332 17380 17388 17382
rect 17412 17380 17468 17382
rect 17492 17380 17548 17382
rect 17572 17380 17628 17382
rect 17332 16346 17388 16348
rect 17412 16346 17468 16348
rect 17492 16346 17548 16348
rect 17572 16346 17628 16348
rect 17332 16294 17378 16346
rect 17378 16294 17388 16346
rect 17412 16294 17442 16346
rect 17442 16294 17454 16346
rect 17454 16294 17468 16346
rect 17492 16294 17506 16346
rect 17506 16294 17518 16346
rect 17518 16294 17548 16346
rect 17572 16294 17582 16346
rect 17582 16294 17628 16346
rect 17332 16292 17388 16294
rect 17412 16292 17468 16294
rect 17492 16292 17548 16294
rect 17572 16292 17628 16294
rect 17332 15258 17388 15260
rect 17412 15258 17468 15260
rect 17492 15258 17548 15260
rect 17572 15258 17628 15260
rect 17332 15206 17378 15258
rect 17378 15206 17388 15258
rect 17412 15206 17442 15258
rect 17442 15206 17454 15258
rect 17454 15206 17468 15258
rect 17492 15206 17506 15258
rect 17506 15206 17518 15258
rect 17518 15206 17548 15258
rect 17572 15206 17582 15258
rect 17582 15206 17628 15258
rect 17332 15204 17388 15206
rect 17412 15204 17468 15206
rect 17492 15204 17548 15206
rect 17572 15204 17628 15206
rect 17332 14170 17388 14172
rect 17412 14170 17468 14172
rect 17492 14170 17548 14172
rect 17572 14170 17628 14172
rect 17332 14118 17378 14170
rect 17378 14118 17388 14170
rect 17412 14118 17442 14170
rect 17442 14118 17454 14170
rect 17454 14118 17468 14170
rect 17492 14118 17506 14170
rect 17506 14118 17518 14170
rect 17518 14118 17548 14170
rect 17572 14118 17582 14170
rect 17582 14118 17628 14170
rect 17332 14116 17388 14118
rect 17412 14116 17468 14118
rect 17492 14116 17548 14118
rect 17572 14116 17628 14118
rect 13238 13626 13294 13628
rect 13318 13626 13374 13628
rect 13398 13626 13454 13628
rect 13478 13626 13534 13628
rect 13238 13574 13284 13626
rect 13284 13574 13294 13626
rect 13318 13574 13348 13626
rect 13348 13574 13360 13626
rect 13360 13574 13374 13626
rect 13398 13574 13412 13626
rect 13412 13574 13424 13626
rect 13424 13574 13454 13626
rect 13478 13574 13488 13626
rect 13488 13574 13534 13626
rect 13238 13572 13294 13574
rect 13318 13572 13374 13574
rect 13398 13572 13454 13574
rect 13478 13572 13534 13574
rect 13238 12538 13294 12540
rect 13318 12538 13374 12540
rect 13398 12538 13454 12540
rect 13478 12538 13534 12540
rect 13238 12486 13284 12538
rect 13284 12486 13294 12538
rect 13318 12486 13348 12538
rect 13348 12486 13360 12538
rect 13360 12486 13374 12538
rect 13398 12486 13412 12538
rect 13412 12486 13424 12538
rect 13424 12486 13454 12538
rect 13478 12486 13488 12538
rect 13488 12486 13534 12538
rect 13238 12484 13294 12486
rect 13318 12484 13374 12486
rect 13398 12484 13454 12486
rect 13478 12484 13534 12486
rect 13238 11450 13294 11452
rect 13318 11450 13374 11452
rect 13398 11450 13454 11452
rect 13478 11450 13534 11452
rect 13238 11398 13284 11450
rect 13284 11398 13294 11450
rect 13318 11398 13348 11450
rect 13348 11398 13360 11450
rect 13360 11398 13374 11450
rect 13398 11398 13412 11450
rect 13412 11398 13424 11450
rect 13424 11398 13454 11450
rect 13478 11398 13488 11450
rect 13488 11398 13534 11450
rect 13238 11396 13294 11398
rect 13318 11396 13374 11398
rect 13398 11396 13454 11398
rect 13478 11396 13534 11398
rect 9144 8730 9200 8732
rect 9224 8730 9280 8732
rect 9304 8730 9360 8732
rect 9384 8730 9440 8732
rect 9144 8678 9190 8730
rect 9190 8678 9200 8730
rect 9224 8678 9254 8730
rect 9254 8678 9266 8730
rect 9266 8678 9280 8730
rect 9304 8678 9318 8730
rect 9318 8678 9330 8730
rect 9330 8678 9360 8730
rect 9384 8678 9394 8730
rect 9394 8678 9440 8730
rect 9144 8676 9200 8678
rect 9224 8676 9280 8678
rect 9304 8676 9360 8678
rect 9384 8676 9440 8678
rect 9144 7642 9200 7644
rect 9224 7642 9280 7644
rect 9304 7642 9360 7644
rect 9384 7642 9440 7644
rect 9144 7590 9190 7642
rect 9190 7590 9200 7642
rect 9224 7590 9254 7642
rect 9254 7590 9266 7642
rect 9266 7590 9280 7642
rect 9304 7590 9318 7642
rect 9318 7590 9330 7642
rect 9330 7590 9360 7642
rect 9384 7590 9394 7642
rect 9394 7590 9440 7642
rect 9144 7588 9200 7590
rect 9224 7588 9280 7590
rect 9304 7588 9360 7590
rect 9384 7588 9440 7590
rect 13238 10362 13294 10364
rect 13318 10362 13374 10364
rect 13398 10362 13454 10364
rect 13478 10362 13534 10364
rect 13238 10310 13284 10362
rect 13284 10310 13294 10362
rect 13318 10310 13348 10362
rect 13348 10310 13360 10362
rect 13360 10310 13374 10362
rect 13398 10310 13412 10362
rect 13412 10310 13424 10362
rect 13424 10310 13454 10362
rect 13478 10310 13488 10362
rect 13488 10310 13534 10362
rect 13238 10308 13294 10310
rect 13318 10308 13374 10310
rect 13398 10308 13454 10310
rect 13478 10308 13534 10310
rect 13238 9274 13294 9276
rect 13318 9274 13374 9276
rect 13398 9274 13454 9276
rect 13478 9274 13534 9276
rect 13238 9222 13284 9274
rect 13284 9222 13294 9274
rect 13318 9222 13348 9274
rect 13348 9222 13360 9274
rect 13360 9222 13374 9274
rect 13398 9222 13412 9274
rect 13412 9222 13424 9274
rect 13424 9222 13454 9274
rect 13478 9222 13488 9274
rect 13488 9222 13534 9274
rect 13238 9220 13294 9222
rect 13318 9220 13374 9222
rect 13398 9220 13454 9222
rect 13478 9220 13534 9222
rect 13238 8186 13294 8188
rect 13318 8186 13374 8188
rect 13398 8186 13454 8188
rect 13478 8186 13534 8188
rect 13238 8134 13284 8186
rect 13284 8134 13294 8186
rect 13318 8134 13348 8186
rect 13348 8134 13360 8186
rect 13360 8134 13374 8186
rect 13398 8134 13412 8186
rect 13412 8134 13424 8186
rect 13424 8134 13454 8186
rect 13478 8134 13488 8186
rect 13488 8134 13534 8186
rect 13238 8132 13294 8134
rect 13318 8132 13374 8134
rect 13398 8132 13454 8134
rect 13478 8132 13534 8134
rect 13238 7098 13294 7100
rect 13318 7098 13374 7100
rect 13398 7098 13454 7100
rect 13478 7098 13534 7100
rect 13238 7046 13284 7098
rect 13284 7046 13294 7098
rect 13318 7046 13348 7098
rect 13348 7046 13360 7098
rect 13360 7046 13374 7098
rect 13398 7046 13412 7098
rect 13412 7046 13424 7098
rect 13424 7046 13454 7098
rect 13478 7046 13488 7098
rect 13488 7046 13534 7098
rect 13238 7044 13294 7046
rect 13318 7044 13374 7046
rect 13398 7044 13454 7046
rect 13478 7044 13534 7046
rect 9144 6554 9200 6556
rect 9224 6554 9280 6556
rect 9304 6554 9360 6556
rect 9384 6554 9440 6556
rect 9144 6502 9190 6554
rect 9190 6502 9200 6554
rect 9224 6502 9254 6554
rect 9254 6502 9266 6554
rect 9266 6502 9280 6554
rect 9304 6502 9318 6554
rect 9318 6502 9330 6554
rect 9330 6502 9360 6554
rect 9384 6502 9394 6554
rect 9394 6502 9440 6554
rect 9144 6500 9200 6502
rect 9224 6500 9280 6502
rect 9304 6500 9360 6502
rect 9384 6500 9440 6502
rect 9144 5466 9200 5468
rect 9224 5466 9280 5468
rect 9304 5466 9360 5468
rect 9384 5466 9440 5468
rect 9144 5414 9190 5466
rect 9190 5414 9200 5466
rect 9224 5414 9254 5466
rect 9254 5414 9266 5466
rect 9266 5414 9280 5466
rect 9304 5414 9318 5466
rect 9318 5414 9330 5466
rect 9330 5414 9360 5466
rect 9384 5414 9394 5466
rect 9394 5414 9440 5466
rect 9144 5412 9200 5414
rect 9224 5412 9280 5414
rect 9304 5412 9360 5414
rect 9384 5412 9440 5414
rect 9144 4378 9200 4380
rect 9224 4378 9280 4380
rect 9304 4378 9360 4380
rect 9384 4378 9440 4380
rect 9144 4326 9190 4378
rect 9190 4326 9200 4378
rect 9224 4326 9254 4378
rect 9254 4326 9266 4378
rect 9266 4326 9280 4378
rect 9304 4326 9318 4378
rect 9318 4326 9330 4378
rect 9330 4326 9360 4378
rect 9384 4326 9394 4378
rect 9394 4326 9440 4378
rect 9144 4324 9200 4326
rect 9224 4324 9280 4326
rect 9304 4324 9360 4326
rect 9384 4324 9440 4326
rect 9144 3290 9200 3292
rect 9224 3290 9280 3292
rect 9304 3290 9360 3292
rect 9384 3290 9440 3292
rect 9144 3238 9190 3290
rect 9190 3238 9200 3290
rect 9224 3238 9254 3290
rect 9254 3238 9266 3290
rect 9266 3238 9280 3290
rect 9304 3238 9318 3290
rect 9318 3238 9330 3290
rect 9330 3238 9360 3290
rect 9384 3238 9394 3290
rect 9394 3238 9440 3290
rect 9144 3236 9200 3238
rect 9224 3236 9280 3238
rect 9304 3236 9360 3238
rect 9384 3236 9440 3238
rect 13238 6010 13294 6012
rect 13318 6010 13374 6012
rect 13398 6010 13454 6012
rect 13478 6010 13534 6012
rect 13238 5958 13284 6010
rect 13284 5958 13294 6010
rect 13318 5958 13348 6010
rect 13348 5958 13360 6010
rect 13360 5958 13374 6010
rect 13398 5958 13412 6010
rect 13412 5958 13424 6010
rect 13424 5958 13454 6010
rect 13478 5958 13488 6010
rect 13488 5958 13534 6010
rect 13238 5956 13294 5958
rect 13318 5956 13374 5958
rect 13398 5956 13454 5958
rect 13478 5956 13534 5958
rect 9144 2202 9200 2204
rect 9224 2202 9280 2204
rect 9304 2202 9360 2204
rect 9384 2202 9440 2204
rect 9144 2150 9190 2202
rect 9190 2150 9200 2202
rect 9224 2150 9254 2202
rect 9254 2150 9266 2202
rect 9266 2150 9280 2202
rect 9304 2150 9318 2202
rect 9318 2150 9330 2202
rect 9330 2150 9360 2202
rect 9384 2150 9394 2202
rect 9394 2150 9440 2202
rect 9144 2148 9200 2150
rect 9224 2148 9280 2150
rect 9304 2148 9360 2150
rect 9384 2148 9440 2150
rect 17332 13082 17388 13084
rect 17412 13082 17468 13084
rect 17492 13082 17548 13084
rect 17572 13082 17628 13084
rect 17332 13030 17378 13082
rect 17378 13030 17388 13082
rect 17412 13030 17442 13082
rect 17442 13030 17454 13082
rect 17454 13030 17468 13082
rect 17492 13030 17506 13082
rect 17506 13030 17518 13082
rect 17518 13030 17548 13082
rect 17572 13030 17582 13082
rect 17582 13030 17628 13082
rect 17332 13028 17388 13030
rect 17412 13028 17468 13030
rect 17492 13028 17548 13030
rect 17572 13028 17628 13030
rect 17332 11994 17388 11996
rect 17412 11994 17468 11996
rect 17492 11994 17548 11996
rect 17572 11994 17628 11996
rect 17332 11942 17378 11994
rect 17378 11942 17388 11994
rect 17412 11942 17442 11994
rect 17442 11942 17454 11994
rect 17454 11942 17468 11994
rect 17492 11942 17506 11994
rect 17506 11942 17518 11994
rect 17518 11942 17548 11994
rect 17572 11942 17582 11994
rect 17582 11942 17628 11994
rect 17332 11940 17388 11942
rect 17412 11940 17468 11942
rect 17492 11940 17548 11942
rect 17572 11940 17628 11942
rect 17332 10906 17388 10908
rect 17412 10906 17468 10908
rect 17492 10906 17548 10908
rect 17572 10906 17628 10908
rect 17332 10854 17378 10906
rect 17378 10854 17388 10906
rect 17412 10854 17442 10906
rect 17442 10854 17454 10906
rect 17454 10854 17468 10906
rect 17492 10854 17506 10906
rect 17506 10854 17518 10906
rect 17518 10854 17548 10906
rect 17572 10854 17582 10906
rect 17582 10854 17628 10906
rect 17332 10852 17388 10854
rect 17412 10852 17468 10854
rect 17492 10852 17548 10854
rect 17572 10852 17628 10854
rect 13238 4922 13294 4924
rect 13318 4922 13374 4924
rect 13398 4922 13454 4924
rect 13478 4922 13534 4924
rect 13238 4870 13284 4922
rect 13284 4870 13294 4922
rect 13318 4870 13348 4922
rect 13348 4870 13360 4922
rect 13360 4870 13374 4922
rect 13398 4870 13412 4922
rect 13412 4870 13424 4922
rect 13424 4870 13454 4922
rect 13478 4870 13488 4922
rect 13488 4870 13534 4922
rect 13238 4868 13294 4870
rect 13318 4868 13374 4870
rect 13398 4868 13454 4870
rect 13478 4868 13534 4870
rect 13238 3834 13294 3836
rect 13318 3834 13374 3836
rect 13398 3834 13454 3836
rect 13478 3834 13534 3836
rect 13238 3782 13284 3834
rect 13284 3782 13294 3834
rect 13318 3782 13348 3834
rect 13348 3782 13360 3834
rect 13360 3782 13374 3834
rect 13398 3782 13412 3834
rect 13412 3782 13424 3834
rect 13424 3782 13454 3834
rect 13478 3782 13488 3834
rect 13488 3782 13534 3834
rect 13238 3780 13294 3782
rect 13318 3780 13374 3782
rect 13398 3780 13454 3782
rect 13478 3780 13534 3782
rect 17332 9818 17388 9820
rect 17412 9818 17468 9820
rect 17492 9818 17548 9820
rect 17572 9818 17628 9820
rect 17332 9766 17378 9818
rect 17378 9766 17388 9818
rect 17412 9766 17442 9818
rect 17442 9766 17454 9818
rect 17454 9766 17468 9818
rect 17492 9766 17506 9818
rect 17506 9766 17518 9818
rect 17518 9766 17548 9818
rect 17572 9766 17582 9818
rect 17582 9766 17628 9818
rect 17332 9764 17388 9766
rect 17412 9764 17468 9766
rect 17492 9764 17548 9766
rect 17572 9764 17628 9766
rect 17332 8730 17388 8732
rect 17412 8730 17468 8732
rect 17492 8730 17548 8732
rect 17572 8730 17628 8732
rect 17332 8678 17378 8730
rect 17378 8678 17388 8730
rect 17412 8678 17442 8730
rect 17442 8678 17454 8730
rect 17454 8678 17468 8730
rect 17492 8678 17506 8730
rect 17506 8678 17518 8730
rect 17518 8678 17548 8730
rect 17572 8678 17582 8730
rect 17582 8678 17628 8730
rect 17332 8676 17388 8678
rect 17412 8676 17468 8678
rect 17492 8676 17548 8678
rect 17572 8676 17628 8678
rect 17332 7642 17388 7644
rect 17412 7642 17468 7644
rect 17492 7642 17548 7644
rect 17572 7642 17628 7644
rect 17332 7590 17378 7642
rect 17378 7590 17388 7642
rect 17412 7590 17442 7642
rect 17442 7590 17454 7642
rect 17454 7590 17468 7642
rect 17492 7590 17506 7642
rect 17506 7590 17518 7642
rect 17518 7590 17548 7642
rect 17572 7590 17582 7642
rect 17582 7590 17628 7642
rect 17332 7588 17388 7590
rect 17412 7588 17468 7590
rect 17492 7588 17548 7590
rect 17572 7588 17628 7590
rect 13238 2746 13294 2748
rect 13318 2746 13374 2748
rect 13398 2746 13454 2748
rect 13478 2746 13534 2748
rect 13238 2694 13284 2746
rect 13284 2694 13294 2746
rect 13318 2694 13348 2746
rect 13348 2694 13360 2746
rect 13360 2694 13374 2746
rect 13398 2694 13412 2746
rect 13412 2694 13424 2746
rect 13424 2694 13454 2746
rect 13478 2694 13488 2746
rect 13488 2694 13534 2746
rect 13238 2692 13294 2694
rect 13318 2692 13374 2694
rect 13398 2692 13454 2694
rect 13478 2692 13534 2694
rect 17332 6554 17388 6556
rect 17412 6554 17468 6556
rect 17492 6554 17548 6556
rect 17572 6554 17628 6556
rect 17332 6502 17378 6554
rect 17378 6502 17388 6554
rect 17412 6502 17442 6554
rect 17442 6502 17454 6554
rect 17454 6502 17468 6554
rect 17492 6502 17506 6554
rect 17506 6502 17518 6554
rect 17518 6502 17548 6554
rect 17572 6502 17582 6554
rect 17582 6502 17628 6554
rect 17332 6500 17388 6502
rect 17412 6500 17468 6502
rect 17492 6500 17548 6502
rect 17572 6500 17628 6502
rect 17332 5466 17388 5468
rect 17412 5466 17468 5468
rect 17492 5466 17548 5468
rect 17572 5466 17628 5468
rect 17332 5414 17378 5466
rect 17378 5414 17388 5466
rect 17412 5414 17442 5466
rect 17442 5414 17454 5466
rect 17454 5414 17468 5466
rect 17492 5414 17506 5466
rect 17506 5414 17518 5466
rect 17518 5414 17548 5466
rect 17572 5414 17582 5466
rect 17582 5414 17628 5466
rect 17332 5412 17388 5414
rect 17412 5412 17468 5414
rect 17492 5412 17548 5414
rect 17572 5412 17628 5414
rect 17332 4378 17388 4380
rect 17412 4378 17468 4380
rect 17492 4378 17548 4380
rect 17572 4378 17628 4380
rect 17332 4326 17378 4378
rect 17378 4326 17388 4378
rect 17412 4326 17442 4378
rect 17442 4326 17454 4378
rect 17454 4326 17468 4378
rect 17492 4326 17506 4378
rect 17506 4326 17518 4378
rect 17518 4326 17548 4378
rect 17572 4326 17582 4378
rect 17582 4326 17628 4378
rect 17332 4324 17388 4326
rect 17412 4324 17468 4326
rect 17492 4324 17548 4326
rect 17572 4324 17628 4326
rect 17332 3290 17388 3292
rect 17412 3290 17468 3292
rect 17492 3290 17548 3292
rect 17572 3290 17628 3292
rect 17332 3238 17378 3290
rect 17378 3238 17388 3290
rect 17412 3238 17442 3290
rect 17442 3238 17454 3290
rect 17454 3238 17468 3290
rect 17492 3238 17506 3290
rect 17506 3238 17518 3290
rect 17518 3238 17548 3290
rect 17572 3238 17582 3290
rect 17582 3238 17628 3290
rect 17332 3236 17388 3238
rect 17412 3236 17468 3238
rect 17492 3236 17548 3238
rect 17572 3236 17628 3238
rect 17332 2202 17388 2204
rect 17412 2202 17468 2204
rect 17492 2202 17548 2204
rect 17572 2202 17628 2204
rect 17332 2150 17378 2202
rect 17378 2150 17388 2202
rect 17412 2150 17442 2202
rect 17442 2150 17454 2202
rect 17454 2150 17468 2202
rect 17492 2150 17506 2202
rect 17506 2150 17518 2202
rect 17518 2150 17548 2202
rect 17572 2150 17582 2202
rect 17582 2150 17628 2202
rect 17332 2148 17388 2150
rect 17412 2148 17468 2150
rect 17492 2148 17548 2150
rect 17572 2148 17628 2150
rect 21426 17978 21482 17980
rect 21506 17978 21562 17980
rect 21586 17978 21642 17980
rect 21666 17978 21722 17980
rect 21426 17926 21472 17978
rect 21472 17926 21482 17978
rect 21506 17926 21536 17978
rect 21536 17926 21548 17978
rect 21548 17926 21562 17978
rect 21586 17926 21600 17978
rect 21600 17926 21612 17978
rect 21612 17926 21642 17978
rect 21666 17926 21676 17978
rect 21676 17926 21722 17978
rect 21426 17924 21482 17926
rect 21506 17924 21562 17926
rect 21586 17924 21642 17926
rect 21666 17924 21722 17926
rect 25520 20698 25576 20700
rect 25600 20698 25656 20700
rect 25680 20698 25736 20700
rect 25760 20698 25816 20700
rect 25520 20646 25566 20698
rect 25566 20646 25576 20698
rect 25600 20646 25630 20698
rect 25630 20646 25642 20698
rect 25642 20646 25656 20698
rect 25680 20646 25694 20698
rect 25694 20646 25706 20698
rect 25706 20646 25736 20698
rect 25760 20646 25770 20698
rect 25770 20646 25816 20698
rect 25520 20644 25576 20646
rect 25600 20644 25656 20646
rect 25680 20644 25736 20646
rect 25760 20644 25816 20646
rect 25520 19610 25576 19612
rect 25600 19610 25656 19612
rect 25680 19610 25736 19612
rect 25760 19610 25816 19612
rect 25520 19558 25566 19610
rect 25566 19558 25576 19610
rect 25600 19558 25630 19610
rect 25630 19558 25642 19610
rect 25642 19558 25656 19610
rect 25680 19558 25694 19610
rect 25694 19558 25706 19610
rect 25706 19558 25736 19610
rect 25760 19558 25770 19610
rect 25770 19558 25816 19610
rect 25520 19556 25576 19558
rect 25600 19556 25656 19558
rect 25680 19556 25736 19558
rect 25760 19556 25816 19558
rect 21426 16890 21482 16892
rect 21506 16890 21562 16892
rect 21586 16890 21642 16892
rect 21666 16890 21722 16892
rect 21426 16838 21472 16890
rect 21472 16838 21482 16890
rect 21506 16838 21536 16890
rect 21536 16838 21548 16890
rect 21548 16838 21562 16890
rect 21586 16838 21600 16890
rect 21600 16838 21612 16890
rect 21612 16838 21642 16890
rect 21666 16838 21676 16890
rect 21676 16838 21722 16890
rect 21426 16836 21482 16838
rect 21506 16836 21562 16838
rect 21586 16836 21642 16838
rect 21666 16836 21722 16838
rect 21426 15802 21482 15804
rect 21506 15802 21562 15804
rect 21586 15802 21642 15804
rect 21666 15802 21722 15804
rect 21426 15750 21472 15802
rect 21472 15750 21482 15802
rect 21506 15750 21536 15802
rect 21536 15750 21548 15802
rect 21548 15750 21562 15802
rect 21586 15750 21600 15802
rect 21600 15750 21612 15802
rect 21612 15750 21642 15802
rect 21666 15750 21676 15802
rect 21676 15750 21722 15802
rect 21426 15748 21482 15750
rect 21506 15748 21562 15750
rect 21586 15748 21642 15750
rect 21666 15748 21722 15750
rect 21426 14714 21482 14716
rect 21506 14714 21562 14716
rect 21586 14714 21642 14716
rect 21666 14714 21722 14716
rect 21426 14662 21472 14714
rect 21472 14662 21482 14714
rect 21506 14662 21536 14714
rect 21536 14662 21548 14714
rect 21548 14662 21562 14714
rect 21586 14662 21600 14714
rect 21600 14662 21612 14714
rect 21612 14662 21642 14714
rect 21666 14662 21676 14714
rect 21676 14662 21722 14714
rect 21426 14660 21482 14662
rect 21506 14660 21562 14662
rect 21586 14660 21642 14662
rect 21666 14660 21722 14662
rect 25520 18522 25576 18524
rect 25600 18522 25656 18524
rect 25680 18522 25736 18524
rect 25760 18522 25816 18524
rect 25520 18470 25566 18522
rect 25566 18470 25576 18522
rect 25600 18470 25630 18522
rect 25630 18470 25642 18522
rect 25642 18470 25656 18522
rect 25680 18470 25694 18522
rect 25694 18470 25706 18522
rect 25706 18470 25736 18522
rect 25760 18470 25770 18522
rect 25770 18470 25816 18522
rect 25520 18468 25576 18470
rect 25600 18468 25656 18470
rect 25680 18468 25736 18470
rect 25760 18468 25816 18470
rect 29614 24506 29670 24508
rect 29694 24506 29750 24508
rect 29774 24506 29830 24508
rect 29854 24506 29910 24508
rect 29614 24454 29660 24506
rect 29660 24454 29670 24506
rect 29694 24454 29724 24506
rect 29724 24454 29736 24506
rect 29736 24454 29750 24506
rect 29774 24454 29788 24506
rect 29788 24454 29800 24506
rect 29800 24454 29830 24506
rect 29854 24454 29864 24506
rect 29864 24454 29910 24506
rect 29614 24452 29670 24454
rect 29694 24452 29750 24454
rect 29774 24452 29830 24454
rect 29854 24452 29910 24454
rect 29614 23418 29670 23420
rect 29694 23418 29750 23420
rect 29774 23418 29830 23420
rect 29854 23418 29910 23420
rect 29614 23366 29660 23418
rect 29660 23366 29670 23418
rect 29694 23366 29724 23418
rect 29724 23366 29736 23418
rect 29736 23366 29750 23418
rect 29774 23366 29788 23418
rect 29788 23366 29800 23418
rect 29800 23366 29830 23418
rect 29854 23366 29864 23418
rect 29864 23366 29910 23418
rect 29614 23364 29670 23366
rect 29694 23364 29750 23366
rect 29774 23364 29830 23366
rect 29854 23364 29910 23366
rect 29614 22330 29670 22332
rect 29694 22330 29750 22332
rect 29774 22330 29830 22332
rect 29854 22330 29910 22332
rect 29614 22278 29660 22330
rect 29660 22278 29670 22330
rect 29694 22278 29724 22330
rect 29724 22278 29736 22330
rect 29736 22278 29750 22330
rect 29774 22278 29788 22330
rect 29788 22278 29800 22330
rect 29800 22278 29830 22330
rect 29854 22278 29864 22330
rect 29864 22278 29910 22330
rect 29614 22276 29670 22278
rect 29694 22276 29750 22278
rect 29774 22276 29830 22278
rect 29854 22276 29910 22278
rect 29614 21242 29670 21244
rect 29694 21242 29750 21244
rect 29774 21242 29830 21244
rect 29854 21242 29910 21244
rect 29614 21190 29660 21242
rect 29660 21190 29670 21242
rect 29694 21190 29724 21242
rect 29724 21190 29736 21242
rect 29736 21190 29750 21242
rect 29774 21190 29788 21242
rect 29788 21190 29800 21242
rect 29800 21190 29830 21242
rect 29854 21190 29864 21242
rect 29864 21190 29910 21242
rect 29614 21188 29670 21190
rect 29694 21188 29750 21190
rect 29774 21188 29830 21190
rect 29854 21188 29910 21190
rect 29614 20154 29670 20156
rect 29694 20154 29750 20156
rect 29774 20154 29830 20156
rect 29854 20154 29910 20156
rect 29614 20102 29660 20154
rect 29660 20102 29670 20154
rect 29694 20102 29724 20154
rect 29724 20102 29736 20154
rect 29736 20102 29750 20154
rect 29774 20102 29788 20154
rect 29788 20102 29800 20154
rect 29800 20102 29830 20154
rect 29854 20102 29864 20154
rect 29864 20102 29910 20154
rect 29614 20100 29670 20102
rect 29694 20100 29750 20102
rect 29774 20100 29830 20102
rect 29854 20100 29910 20102
rect 25520 17434 25576 17436
rect 25600 17434 25656 17436
rect 25680 17434 25736 17436
rect 25760 17434 25816 17436
rect 25520 17382 25566 17434
rect 25566 17382 25576 17434
rect 25600 17382 25630 17434
rect 25630 17382 25642 17434
rect 25642 17382 25656 17434
rect 25680 17382 25694 17434
rect 25694 17382 25706 17434
rect 25706 17382 25736 17434
rect 25760 17382 25770 17434
rect 25770 17382 25816 17434
rect 25520 17380 25576 17382
rect 25600 17380 25656 17382
rect 25680 17380 25736 17382
rect 25760 17380 25816 17382
rect 25520 16346 25576 16348
rect 25600 16346 25656 16348
rect 25680 16346 25736 16348
rect 25760 16346 25816 16348
rect 25520 16294 25566 16346
rect 25566 16294 25576 16346
rect 25600 16294 25630 16346
rect 25630 16294 25642 16346
rect 25642 16294 25656 16346
rect 25680 16294 25694 16346
rect 25694 16294 25706 16346
rect 25706 16294 25736 16346
rect 25760 16294 25770 16346
rect 25770 16294 25816 16346
rect 25520 16292 25576 16294
rect 25600 16292 25656 16294
rect 25680 16292 25736 16294
rect 25760 16292 25816 16294
rect 21426 13626 21482 13628
rect 21506 13626 21562 13628
rect 21586 13626 21642 13628
rect 21666 13626 21722 13628
rect 21426 13574 21472 13626
rect 21472 13574 21482 13626
rect 21506 13574 21536 13626
rect 21536 13574 21548 13626
rect 21548 13574 21562 13626
rect 21586 13574 21600 13626
rect 21600 13574 21612 13626
rect 21612 13574 21642 13626
rect 21666 13574 21676 13626
rect 21676 13574 21722 13626
rect 21426 13572 21482 13574
rect 21506 13572 21562 13574
rect 21586 13572 21642 13574
rect 21666 13572 21722 13574
rect 21426 12538 21482 12540
rect 21506 12538 21562 12540
rect 21586 12538 21642 12540
rect 21666 12538 21722 12540
rect 21426 12486 21472 12538
rect 21472 12486 21482 12538
rect 21506 12486 21536 12538
rect 21536 12486 21548 12538
rect 21548 12486 21562 12538
rect 21586 12486 21600 12538
rect 21600 12486 21612 12538
rect 21612 12486 21642 12538
rect 21666 12486 21676 12538
rect 21676 12486 21722 12538
rect 21426 12484 21482 12486
rect 21506 12484 21562 12486
rect 21586 12484 21642 12486
rect 21666 12484 21722 12486
rect 21426 11450 21482 11452
rect 21506 11450 21562 11452
rect 21586 11450 21642 11452
rect 21666 11450 21722 11452
rect 21426 11398 21472 11450
rect 21472 11398 21482 11450
rect 21506 11398 21536 11450
rect 21536 11398 21548 11450
rect 21548 11398 21562 11450
rect 21586 11398 21600 11450
rect 21600 11398 21612 11450
rect 21612 11398 21642 11450
rect 21666 11398 21676 11450
rect 21676 11398 21722 11450
rect 21426 11396 21482 11398
rect 21506 11396 21562 11398
rect 21586 11396 21642 11398
rect 21666 11396 21722 11398
rect 21426 10362 21482 10364
rect 21506 10362 21562 10364
rect 21586 10362 21642 10364
rect 21666 10362 21722 10364
rect 21426 10310 21472 10362
rect 21472 10310 21482 10362
rect 21506 10310 21536 10362
rect 21536 10310 21548 10362
rect 21548 10310 21562 10362
rect 21586 10310 21600 10362
rect 21600 10310 21612 10362
rect 21612 10310 21642 10362
rect 21666 10310 21676 10362
rect 21676 10310 21722 10362
rect 21426 10308 21482 10310
rect 21506 10308 21562 10310
rect 21586 10308 21642 10310
rect 21666 10308 21722 10310
rect 21426 9274 21482 9276
rect 21506 9274 21562 9276
rect 21586 9274 21642 9276
rect 21666 9274 21722 9276
rect 21426 9222 21472 9274
rect 21472 9222 21482 9274
rect 21506 9222 21536 9274
rect 21536 9222 21548 9274
rect 21548 9222 21562 9274
rect 21586 9222 21600 9274
rect 21600 9222 21612 9274
rect 21612 9222 21642 9274
rect 21666 9222 21676 9274
rect 21676 9222 21722 9274
rect 21426 9220 21482 9222
rect 21506 9220 21562 9222
rect 21586 9220 21642 9222
rect 21666 9220 21722 9222
rect 21426 8186 21482 8188
rect 21506 8186 21562 8188
rect 21586 8186 21642 8188
rect 21666 8186 21722 8188
rect 21426 8134 21472 8186
rect 21472 8134 21482 8186
rect 21506 8134 21536 8186
rect 21536 8134 21548 8186
rect 21548 8134 21562 8186
rect 21586 8134 21600 8186
rect 21600 8134 21612 8186
rect 21612 8134 21642 8186
rect 21666 8134 21676 8186
rect 21676 8134 21722 8186
rect 21426 8132 21482 8134
rect 21506 8132 21562 8134
rect 21586 8132 21642 8134
rect 21666 8132 21722 8134
rect 21426 7098 21482 7100
rect 21506 7098 21562 7100
rect 21586 7098 21642 7100
rect 21666 7098 21722 7100
rect 21426 7046 21472 7098
rect 21472 7046 21482 7098
rect 21506 7046 21536 7098
rect 21536 7046 21548 7098
rect 21548 7046 21562 7098
rect 21586 7046 21600 7098
rect 21600 7046 21612 7098
rect 21612 7046 21642 7098
rect 21666 7046 21676 7098
rect 21676 7046 21722 7098
rect 21426 7044 21482 7046
rect 21506 7044 21562 7046
rect 21586 7044 21642 7046
rect 21666 7044 21722 7046
rect 21426 6010 21482 6012
rect 21506 6010 21562 6012
rect 21586 6010 21642 6012
rect 21666 6010 21722 6012
rect 21426 5958 21472 6010
rect 21472 5958 21482 6010
rect 21506 5958 21536 6010
rect 21536 5958 21548 6010
rect 21548 5958 21562 6010
rect 21586 5958 21600 6010
rect 21600 5958 21612 6010
rect 21612 5958 21642 6010
rect 21666 5958 21676 6010
rect 21676 5958 21722 6010
rect 21426 5956 21482 5958
rect 21506 5956 21562 5958
rect 21586 5956 21642 5958
rect 21666 5956 21722 5958
rect 21426 4922 21482 4924
rect 21506 4922 21562 4924
rect 21586 4922 21642 4924
rect 21666 4922 21722 4924
rect 21426 4870 21472 4922
rect 21472 4870 21482 4922
rect 21506 4870 21536 4922
rect 21536 4870 21548 4922
rect 21548 4870 21562 4922
rect 21586 4870 21600 4922
rect 21600 4870 21612 4922
rect 21612 4870 21642 4922
rect 21666 4870 21676 4922
rect 21676 4870 21722 4922
rect 21426 4868 21482 4870
rect 21506 4868 21562 4870
rect 21586 4868 21642 4870
rect 21666 4868 21722 4870
rect 21426 3834 21482 3836
rect 21506 3834 21562 3836
rect 21586 3834 21642 3836
rect 21666 3834 21722 3836
rect 21426 3782 21472 3834
rect 21472 3782 21482 3834
rect 21506 3782 21536 3834
rect 21536 3782 21548 3834
rect 21548 3782 21562 3834
rect 21586 3782 21600 3834
rect 21600 3782 21612 3834
rect 21612 3782 21642 3834
rect 21666 3782 21676 3834
rect 21676 3782 21722 3834
rect 21426 3780 21482 3782
rect 21506 3780 21562 3782
rect 21586 3780 21642 3782
rect 21666 3780 21722 3782
rect 21426 2746 21482 2748
rect 21506 2746 21562 2748
rect 21586 2746 21642 2748
rect 21666 2746 21722 2748
rect 21426 2694 21472 2746
rect 21472 2694 21482 2746
rect 21506 2694 21536 2746
rect 21536 2694 21548 2746
rect 21548 2694 21562 2746
rect 21586 2694 21600 2746
rect 21600 2694 21612 2746
rect 21612 2694 21642 2746
rect 21666 2694 21676 2746
rect 21676 2694 21722 2746
rect 21426 2692 21482 2694
rect 21506 2692 21562 2694
rect 21586 2692 21642 2694
rect 21666 2692 21722 2694
rect 25520 15258 25576 15260
rect 25600 15258 25656 15260
rect 25680 15258 25736 15260
rect 25760 15258 25816 15260
rect 25520 15206 25566 15258
rect 25566 15206 25576 15258
rect 25600 15206 25630 15258
rect 25630 15206 25642 15258
rect 25642 15206 25656 15258
rect 25680 15206 25694 15258
rect 25694 15206 25706 15258
rect 25706 15206 25736 15258
rect 25760 15206 25770 15258
rect 25770 15206 25816 15258
rect 25520 15204 25576 15206
rect 25600 15204 25656 15206
rect 25680 15204 25736 15206
rect 25760 15204 25816 15206
rect 25520 14170 25576 14172
rect 25600 14170 25656 14172
rect 25680 14170 25736 14172
rect 25760 14170 25816 14172
rect 25520 14118 25566 14170
rect 25566 14118 25576 14170
rect 25600 14118 25630 14170
rect 25630 14118 25642 14170
rect 25642 14118 25656 14170
rect 25680 14118 25694 14170
rect 25694 14118 25706 14170
rect 25706 14118 25736 14170
rect 25760 14118 25770 14170
rect 25770 14118 25816 14170
rect 25520 14116 25576 14118
rect 25600 14116 25656 14118
rect 25680 14116 25736 14118
rect 25760 14116 25816 14118
rect 25520 13082 25576 13084
rect 25600 13082 25656 13084
rect 25680 13082 25736 13084
rect 25760 13082 25816 13084
rect 25520 13030 25566 13082
rect 25566 13030 25576 13082
rect 25600 13030 25630 13082
rect 25630 13030 25642 13082
rect 25642 13030 25656 13082
rect 25680 13030 25694 13082
rect 25694 13030 25706 13082
rect 25706 13030 25736 13082
rect 25760 13030 25770 13082
rect 25770 13030 25816 13082
rect 25520 13028 25576 13030
rect 25600 13028 25656 13030
rect 25680 13028 25736 13030
rect 25760 13028 25816 13030
rect 25520 11994 25576 11996
rect 25600 11994 25656 11996
rect 25680 11994 25736 11996
rect 25760 11994 25816 11996
rect 25520 11942 25566 11994
rect 25566 11942 25576 11994
rect 25600 11942 25630 11994
rect 25630 11942 25642 11994
rect 25642 11942 25656 11994
rect 25680 11942 25694 11994
rect 25694 11942 25706 11994
rect 25706 11942 25736 11994
rect 25760 11942 25770 11994
rect 25770 11942 25816 11994
rect 25520 11940 25576 11942
rect 25600 11940 25656 11942
rect 25680 11940 25736 11942
rect 25760 11940 25816 11942
rect 25520 10906 25576 10908
rect 25600 10906 25656 10908
rect 25680 10906 25736 10908
rect 25760 10906 25816 10908
rect 25520 10854 25566 10906
rect 25566 10854 25576 10906
rect 25600 10854 25630 10906
rect 25630 10854 25642 10906
rect 25642 10854 25656 10906
rect 25680 10854 25694 10906
rect 25694 10854 25706 10906
rect 25706 10854 25736 10906
rect 25760 10854 25770 10906
rect 25770 10854 25816 10906
rect 25520 10852 25576 10854
rect 25600 10852 25656 10854
rect 25680 10852 25736 10854
rect 25760 10852 25816 10854
rect 29614 19066 29670 19068
rect 29694 19066 29750 19068
rect 29774 19066 29830 19068
rect 29854 19066 29910 19068
rect 29614 19014 29660 19066
rect 29660 19014 29670 19066
rect 29694 19014 29724 19066
rect 29724 19014 29736 19066
rect 29736 19014 29750 19066
rect 29774 19014 29788 19066
rect 29788 19014 29800 19066
rect 29800 19014 29830 19066
rect 29854 19014 29864 19066
rect 29864 19014 29910 19066
rect 29614 19012 29670 19014
rect 29694 19012 29750 19014
rect 29774 19012 29830 19014
rect 29854 19012 29910 19014
rect 29614 17978 29670 17980
rect 29694 17978 29750 17980
rect 29774 17978 29830 17980
rect 29854 17978 29910 17980
rect 29614 17926 29660 17978
rect 29660 17926 29670 17978
rect 29694 17926 29724 17978
rect 29724 17926 29736 17978
rect 29736 17926 29750 17978
rect 29774 17926 29788 17978
rect 29788 17926 29800 17978
rect 29800 17926 29830 17978
rect 29854 17926 29864 17978
rect 29864 17926 29910 17978
rect 29614 17924 29670 17926
rect 29694 17924 29750 17926
rect 29774 17924 29830 17926
rect 29854 17924 29910 17926
rect 32954 30232 33010 30288
rect 33708 32666 33764 32668
rect 33788 32666 33844 32668
rect 33868 32666 33924 32668
rect 33948 32666 34004 32668
rect 33708 32614 33754 32666
rect 33754 32614 33764 32666
rect 33788 32614 33818 32666
rect 33818 32614 33830 32666
rect 33830 32614 33844 32666
rect 33868 32614 33882 32666
rect 33882 32614 33894 32666
rect 33894 32614 33924 32666
rect 33948 32614 33958 32666
rect 33958 32614 34004 32666
rect 33708 32612 33764 32614
rect 33788 32612 33844 32614
rect 33868 32612 33924 32614
rect 33948 32612 34004 32614
rect 33708 31578 33764 31580
rect 33788 31578 33844 31580
rect 33868 31578 33924 31580
rect 33948 31578 34004 31580
rect 33708 31526 33754 31578
rect 33754 31526 33764 31578
rect 33788 31526 33818 31578
rect 33818 31526 33830 31578
rect 33830 31526 33844 31578
rect 33868 31526 33882 31578
rect 33882 31526 33894 31578
rect 33894 31526 33924 31578
rect 33948 31526 33958 31578
rect 33958 31526 34004 31578
rect 33708 31524 33764 31526
rect 33788 31524 33844 31526
rect 33868 31524 33924 31526
rect 33948 31524 34004 31526
rect 33708 30490 33764 30492
rect 33788 30490 33844 30492
rect 33868 30490 33924 30492
rect 33948 30490 34004 30492
rect 33708 30438 33754 30490
rect 33754 30438 33764 30490
rect 33788 30438 33818 30490
rect 33818 30438 33830 30490
rect 33830 30438 33844 30490
rect 33868 30438 33882 30490
rect 33882 30438 33894 30490
rect 33894 30438 33924 30490
rect 33948 30438 33958 30490
rect 33958 30438 34004 30490
rect 33708 30436 33764 30438
rect 33788 30436 33844 30438
rect 33868 30436 33924 30438
rect 33948 30436 34004 30438
rect 33708 29402 33764 29404
rect 33788 29402 33844 29404
rect 33868 29402 33924 29404
rect 33948 29402 34004 29404
rect 33708 29350 33754 29402
rect 33754 29350 33764 29402
rect 33788 29350 33818 29402
rect 33818 29350 33830 29402
rect 33830 29350 33844 29402
rect 33868 29350 33882 29402
rect 33882 29350 33894 29402
rect 33894 29350 33924 29402
rect 33948 29350 33958 29402
rect 33958 29350 34004 29402
rect 33708 29348 33764 29350
rect 33788 29348 33844 29350
rect 33868 29348 33924 29350
rect 33948 29348 34004 29350
rect 33708 28314 33764 28316
rect 33788 28314 33844 28316
rect 33868 28314 33924 28316
rect 33948 28314 34004 28316
rect 33708 28262 33754 28314
rect 33754 28262 33764 28314
rect 33788 28262 33818 28314
rect 33818 28262 33830 28314
rect 33830 28262 33844 28314
rect 33868 28262 33882 28314
rect 33882 28262 33894 28314
rect 33894 28262 33924 28314
rect 33948 28262 33958 28314
rect 33958 28262 34004 28314
rect 33708 28260 33764 28262
rect 33788 28260 33844 28262
rect 33868 28260 33924 28262
rect 33948 28260 34004 28262
rect 33708 27226 33764 27228
rect 33788 27226 33844 27228
rect 33868 27226 33924 27228
rect 33948 27226 34004 27228
rect 33708 27174 33754 27226
rect 33754 27174 33764 27226
rect 33788 27174 33818 27226
rect 33818 27174 33830 27226
rect 33830 27174 33844 27226
rect 33868 27174 33882 27226
rect 33882 27174 33894 27226
rect 33894 27174 33924 27226
rect 33948 27174 33958 27226
rect 33958 27174 34004 27226
rect 33708 27172 33764 27174
rect 33788 27172 33844 27174
rect 33868 27172 33924 27174
rect 33948 27172 34004 27174
rect 31114 24792 31170 24848
rect 33322 26288 33378 26344
rect 33708 26138 33764 26140
rect 33788 26138 33844 26140
rect 33868 26138 33924 26140
rect 33948 26138 34004 26140
rect 33708 26086 33754 26138
rect 33754 26086 33764 26138
rect 33788 26086 33818 26138
rect 33818 26086 33830 26138
rect 33830 26086 33844 26138
rect 33868 26086 33882 26138
rect 33882 26086 33894 26138
rect 33894 26086 33924 26138
rect 33948 26086 33958 26138
rect 33958 26086 34004 26138
rect 33708 26084 33764 26086
rect 33788 26084 33844 26086
rect 33868 26084 33924 26086
rect 33948 26084 34004 26086
rect 33708 25050 33764 25052
rect 33788 25050 33844 25052
rect 33868 25050 33924 25052
rect 33948 25050 34004 25052
rect 33708 24998 33754 25050
rect 33754 24998 33764 25050
rect 33788 24998 33818 25050
rect 33818 24998 33830 25050
rect 33830 24998 33844 25050
rect 33868 24998 33882 25050
rect 33882 24998 33894 25050
rect 33894 24998 33924 25050
rect 33948 24998 33958 25050
rect 33958 24998 34004 25050
rect 33708 24996 33764 24998
rect 33788 24996 33844 24998
rect 33868 24996 33924 24998
rect 33948 24996 34004 24998
rect 31482 22072 31538 22128
rect 33708 23962 33764 23964
rect 33788 23962 33844 23964
rect 33868 23962 33924 23964
rect 33948 23962 34004 23964
rect 33708 23910 33754 23962
rect 33754 23910 33764 23962
rect 33788 23910 33818 23962
rect 33818 23910 33830 23962
rect 33830 23910 33844 23962
rect 33868 23910 33882 23962
rect 33882 23910 33894 23962
rect 33894 23910 33924 23962
rect 33948 23910 33958 23962
rect 33958 23910 34004 23962
rect 33708 23908 33764 23910
rect 33788 23908 33844 23910
rect 33868 23908 33924 23910
rect 33948 23908 34004 23910
rect 33782 23432 33838 23488
rect 33708 22874 33764 22876
rect 33788 22874 33844 22876
rect 33868 22874 33924 22876
rect 33948 22874 34004 22876
rect 33708 22822 33754 22874
rect 33754 22822 33764 22874
rect 33788 22822 33818 22874
rect 33818 22822 33830 22874
rect 33830 22822 33844 22874
rect 33868 22822 33882 22874
rect 33882 22822 33894 22874
rect 33894 22822 33924 22874
rect 33948 22822 33958 22874
rect 33958 22822 34004 22874
rect 33708 22820 33764 22822
rect 33788 22820 33844 22822
rect 33868 22820 33924 22822
rect 33948 22820 34004 22822
rect 33708 21786 33764 21788
rect 33788 21786 33844 21788
rect 33868 21786 33924 21788
rect 33948 21786 34004 21788
rect 33708 21734 33754 21786
rect 33754 21734 33764 21786
rect 33788 21734 33818 21786
rect 33818 21734 33830 21786
rect 33830 21734 33844 21786
rect 33868 21734 33882 21786
rect 33882 21734 33894 21786
rect 33894 21734 33924 21786
rect 33948 21734 33958 21786
rect 33958 21734 34004 21786
rect 33708 21732 33764 21734
rect 33788 21732 33844 21734
rect 33868 21732 33924 21734
rect 33948 21732 34004 21734
rect 33322 20848 33378 20904
rect 33708 20698 33764 20700
rect 33788 20698 33844 20700
rect 33868 20698 33924 20700
rect 33948 20698 34004 20700
rect 33708 20646 33754 20698
rect 33754 20646 33764 20698
rect 33788 20646 33818 20698
rect 33818 20646 33830 20698
rect 33830 20646 33844 20698
rect 33868 20646 33882 20698
rect 33882 20646 33894 20698
rect 33894 20646 33924 20698
rect 33948 20646 33958 20698
rect 33958 20646 34004 20698
rect 33708 20644 33764 20646
rect 33788 20644 33844 20646
rect 33868 20644 33924 20646
rect 33948 20644 34004 20646
rect 33708 19610 33764 19612
rect 33788 19610 33844 19612
rect 33868 19610 33924 19612
rect 33948 19610 34004 19612
rect 33708 19558 33754 19610
rect 33754 19558 33764 19610
rect 33788 19558 33818 19610
rect 33818 19558 33830 19610
rect 33830 19558 33844 19610
rect 33868 19558 33882 19610
rect 33882 19558 33894 19610
rect 33894 19558 33924 19610
rect 33948 19558 33958 19610
rect 33958 19558 34004 19610
rect 33708 19556 33764 19558
rect 33788 19556 33844 19558
rect 33868 19556 33924 19558
rect 33948 19556 34004 19558
rect 33322 19372 33378 19408
rect 33322 19352 33324 19372
rect 33324 19352 33376 19372
rect 33376 19352 33378 19372
rect 33708 18522 33764 18524
rect 33788 18522 33844 18524
rect 33868 18522 33924 18524
rect 33948 18522 34004 18524
rect 33708 18470 33754 18522
rect 33754 18470 33764 18522
rect 33788 18470 33818 18522
rect 33818 18470 33830 18522
rect 33830 18470 33844 18522
rect 33868 18470 33882 18522
rect 33882 18470 33894 18522
rect 33894 18470 33924 18522
rect 33948 18470 33958 18522
rect 33958 18470 34004 18522
rect 33708 18468 33764 18470
rect 33788 18468 33844 18470
rect 33868 18468 33924 18470
rect 33948 18468 34004 18470
rect 33322 17992 33378 18048
rect 29614 16890 29670 16892
rect 29694 16890 29750 16892
rect 29774 16890 29830 16892
rect 29854 16890 29910 16892
rect 29614 16838 29660 16890
rect 29660 16838 29670 16890
rect 29694 16838 29724 16890
rect 29724 16838 29736 16890
rect 29736 16838 29750 16890
rect 29774 16838 29788 16890
rect 29788 16838 29800 16890
rect 29800 16838 29830 16890
rect 29854 16838 29864 16890
rect 29864 16838 29910 16890
rect 29614 16836 29670 16838
rect 29694 16836 29750 16838
rect 29774 16836 29830 16838
rect 29854 16836 29910 16838
rect 33708 17434 33764 17436
rect 33788 17434 33844 17436
rect 33868 17434 33924 17436
rect 33948 17434 34004 17436
rect 33708 17382 33754 17434
rect 33754 17382 33764 17434
rect 33788 17382 33818 17434
rect 33818 17382 33830 17434
rect 33830 17382 33844 17434
rect 33868 17382 33882 17434
rect 33882 17382 33894 17434
rect 33894 17382 33924 17434
rect 33948 17382 33958 17434
rect 33958 17382 34004 17434
rect 33708 17380 33764 17382
rect 33788 17380 33844 17382
rect 33868 17380 33924 17382
rect 33948 17380 34004 17382
rect 31482 16632 31538 16688
rect 29614 15802 29670 15804
rect 29694 15802 29750 15804
rect 29774 15802 29830 15804
rect 29854 15802 29910 15804
rect 29614 15750 29660 15802
rect 29660 15750 29670 15802
rect 29694 15750 29724 15802
rect 29724 15750 29736 15802
rect 29736 15750 29750 15802
rect 29774 15750 29788 15802
rect 29788 15750 29800 15802
rect 29800 15750 29830 15802
rect 29854 15750 29864 15802
rect 29864 15750 29910 15802
rect 29614 15748 29670 15750
rect 29694 15748 29750 15750
rect 29774 15748 29830 15750
rect 29854 15748 29910 15750
rect 33708 16346 33764 16348
rect 33788 16346 33844 16348
rect 33868 16346 33924 16348
rect 33948 16346 34004 16348
rect 33708 16294 33754 16346
rect 33754 16294 33764 16346
rect 33788 16294 33818 16346
rect 33818 16294 33830 16346
rect 33830 16294 33844 16346
rect 33868 16294 33882 16346
rect 33882 16294 33894 16346
rect 33894 16294 33924 16346
rect 33948 16294 33958 16346
rect 33958 16294 34004 16346
rect 33708 16292 33764 16294
rect 33788 16292 33844 16294
rect 33868 16292 33924 16294
rect 33948 16292 34004 16294
rect 29614 14714 29670 14716
rect 29694 14714 29750 14716
rect 29774 14714 29830 14716
rect 29854 14714 29910 14716
rect 29614 14662 29660 14714
rect 29660 14662 29670 14714
rect 29694 14662 29724 14714
rect 29724 14662 29736 14714
rect 29736 14662 29750 14714
rect 29774 14662 29788 14714
rect 29788 14662 29800 14714
rect 29800 14662 29830 14714
rect 29854 14662 29864 14714
rect 29864 14662 29910 14714
rect 29614 14660 29670 14662
rect 29694 14660 29750 14662
rect 29774 14660 29830 14662
rect 29854 14660 29910 14662
rect 31114 13912 31170 13968
rect 29614 13626 29670 13628
rect 29694 13626 29750 13628
rect 29774 13626 29830 13628
rect 29854 13626 29910 13628
rect 29614 13574 29660 13626
rect 29660 13574 29670 13626
rect 29694 13574 29724 13626
rect 29724 13574 29736 13626
rect 29736 13574 29750 13626
rect 29774 13574 29788 13626
rect 29788 13574 29800 13626
rect 29800 13574 29830 13626
rect 29854 13574 29864 13626
rect 29864 13574 29910 13626
rect 29614 13572 29670 13574
rect 29694 13572 29750 13574
rect 29774 13572 29830 13574
rect 29854 13572 29910 13574
rect 25520 9818 25576 9820
rect 25600 9818 25656 9820
rect 25680 9818 25736 9820
rect 25760 9818 25816 9820
rect 25520 9766 25566 9818
rect 25566 9766 25576 9818
rect 25600 9766 25630 9818
rect 25630 9766 25642 9818
rect 25642 9766 25656 9818
rect 25680 9766 25694 9818
rect 25694 9766 25706 9818
rect 25706 9766 25736 9818
rect 25760 9766 25770 9818
rect 25770 9766 25816 9818
rect 25520 9764 25576 9766
rect 25600 9764 25656 9766
rect 25680 9764 25736 9766
rect 25760 9764 25816 9766
rect 25520 8730 25576 8732
rect 25600 8730 25656 8732
rect 25680 8730 25736 8732
rect 25760 8730 25816 8732
rect 25520 8678 25566 8730
rect 25566 8678 25576 8730
rect 25600 8678 25630 8730
rect 25630 8678 25642 8730
rect 25642 8678 25656 8730
rect 25680 8678 25694 8730
rect 25694 8678 25706 8730
rect 25706 8678 25736 8730
rect 25760 8678 25770 8730
rect 25770 8678 25816 8730
rect 25520 8676 25576 8678
rect 25600 8676 25656 8678
rect 25680 8676 25736 8678
rect 25760 8676 25816 8678
rect 25520 7642 25576 7644
rect 25600 7642 25656 7644
rect 25680 7642 25736 7644
rect 25760 7642 25816 7644
rect 25520 7590 25566 7642
rect 25566 7590 25576 7642
rect 25600 7590 25630 7642
rect 25630 7590 25642 7642
rect 25642 7590 25656 7642
rect 25680 7590 25694 7642
rect 25694 7590 25706 7642
rect 25706 7590 25736 7642
rect 25760 7590 25770 7642
rect 25770 7590 25816 7642
rect 25520 7588 25576 7590
rect 25600 7588 25656 7590
rect 25680 7588 25736 7590
rect 25760 7588 25816 7590
rect 25520 6554 25576 6556
rect 25600 6554 25656 6556
rect 25680 6554 25736 6556
rect 25760 6554 25816 6556
rect 25520 6502 25566 6554
rect 25566 6502 25576 6554
rect 25600 6502 25630 6554
rect 25630 6502 25642 6554
rect 25642 6502 25656 6554
rect 25680 6502 25694 6554
rect 25694 6502 25706 6554
rect 25706 6502 25736 6554
rect 25760 6502 25770 6554
rect 25770 6502 25816 6554
rect 25520 6500 25576 6502
rect 25600 6500 25656 6502
rect 25680 6500 25736 6502
rect 25760 6500 25816 6502
rect 23938 4664 23994 4720
rect 25520 5466 25576 5468
rect 25600 5466 25656 5468
rect 25680 5466 25736 5468
rect 25760 5466 25816 5468
rect 25520 5414 25566 5466
rect 25566 5414 25576 5466
rect 25600 5414 25630 5466
rect 25630 5414 25642 5466
rect 25642 5414 25656 5466
rect 25680 5414 25694 5466
rect 25694 5414 25706 5466
rect 25706 5414 25736 5466
rect 25760 5414 25770 5466
rect 25770 5414 25816 5466
rect 25520 5412 25576 5414
rect 25600 5412 25656 5414
rect 25680 5412 25736 5414
rect 25760 5412 25816 5414
rect 26054 5208 26110 5264
rect 25520 4378 25576 4380
rect 25600 4378 25656 4380
rect 25680 4378 25736 4380
rect 25760 4378 25816 4380
rect 25520 4326 25566 4378
rect 25566 4326 25576 4378
rect 25600 4326 25630 4378
rect 25630 4326 25642 4378
rect 25642 4326 25656 4378
rect 25680 4326 25694 4378
rect 25694 4326 25706 4378
rect 25706 4326 25736 4378
rect 25760 4326 25770 4378
rect 25770 4326 25816 4378
rect 25520 4324 25576 4326
rect 25600 4324 25656 4326
rect 25680 4324 25736 4326
rect 25760 4324 25816 4326
rect 25520 3290 25576 3292
rect 25600 3290 25656 3292
rect 25680 3290 25736 3292
rect 25760 3290 25816 3292
rect 25520 3238 25566 3290
rect 25566 3238 25576 3290
rect 25600 3238 25630 3290
rect 25630 3238 25642 3290
rect 25642 3238 25656 3290
rect 25680 3238 25694 3290
rect 25694 3238 25706 3290
rect 25706 3238 25736 3290
rect 25760 3238 25770 3290
rect 25770 3238 25816 3290
rect 25520 3236 25576 3238
rect 25600 3236 25656 3238
rect 25680 3236 25736 3238
rect 25760 3236 25816 3238
rect 29614 12538 29670 12540
rect 29694 12538 29750 12540
rect 29774 12538 29830 12540
rect 29854 12538 29910 12540
rect 29614 12486 29660 12538
rect 29660 12486 29670 12538
rect 29694 12486 29724 12538
rect 29724 12486 29736 12538
rect 29736 12486 29750 12538
rect 29774 12486 29788 12538
rect 29788 12486 29800 12538
rect 29800 12486 29830 12538
rect 29854 12486 29864 12538
rect 29864 12486 29910 12538
rect 29614 12484 29670 12486
rect 29694 12484 29750 12486
rect 29774 12484 29830 12486
rect 29854 12484 29910 12486
rect 33322 15408 33378 15464
rect 33708 15258 33764 15260
rect 33788 15258 33844 15260
rect 33868 15258 33924 15260
rect 33948 15258 34004 15260
rect 33708 15206 33754 15258
rect 33754 15206 33764 15258
rect 33788 15206 33818 15258
rect 33818 15206 33830 15258
rect 33830 15206 33844 15258
rect 33868 15206 33882 15258
rect 33882 15206 33894 15258
rect 33894 15206 33924 15258
rect 33948 15206 33958 15258
rect 33958 15206 34004 15258
rect 33708 15204 33764 15206
rect 33788 15204 33844 15206
rect 33868 15204 33924 15206
rect 33948 15204 34004 15206
rect 29614 11450 29670 11452
rect 29694 11450 29750 11452
rect 29774 11450 29830 11452
rect 29854 11450 29910 11452
rect 29614 11398 29660 11450
rect 29660 11398 29670 11450
rect 29694 11398 29724 11450
rect 29724 11398 29736 11450
rect 29736 11398 29750 11450
rect 29774 11398 29788 11450
rect 29788 11398 29800 11450
rect 29800 11398 29830 11450
rect 29854 11398 29864 11450
rect 29864 11398 29910 11450
rect 29614 11396 29670 11398
rect 29694 11396 29750 11398
rect 29774 11396 29830 11398
rect 29854 11396 29910 11398
rect 33708 14170 33764 14172
rect 33788 14170 33844 14172
rect 33868 14170 33924 14172
rect 33948 14170 34004 14172
rect 33708 14118 33754 14170
rect 33754 14118 33764 14170
rect 33788 14118 33818 14170
rect 33818 14118 33830 14170
rect 33830 14118 33844 14170
rect 33868 14118 33882 14170
rect 33882 14118 33894 14170
rect 33894 14118 33924 14170
rect 33948 14118 33958 14170
rect 33958 14118 34004 14170
rect 33708 14116 33764 14118
rect 33788 14116 33844 14118
rect 33868 14116 33924 14118
rect 33948 14116 34004 14118
rect 33708 13082 33764 13084
rect 33788 13082 33844 13084
rect 33868 13082 33924 13084
rect 33948 13082 34004 13084
rect 33708 13030 33754 13082
rect 33754 13030 33764 13082
rect 33788 13030 33818 13082
rect 33818 13030 33830 13082
rect 33830 13030 33844 13082
rect 33868 13030 33882 13082
rect 33882 13030 33894 13082
rect 33894 13030 33924 13082
rect 33948 13030 33958 13082
rect 33958 13030 34004 13082
rect 33708 13028 33764 13030
rect 33788 13028 33844 13030
rect 33868 13028 33924 13030
rect 33948 13028 34004 13030
rect 33322 12552 33378 12608
rect 33708 11994 33764 11996
rect 33788 11994 33844 11996
rect 33868 11994 33924 11996
rect 33948 11994 34004 11996
rect 33708 11942 33754 11994
rect 33754 11942 33764 11994
rect 33788 11942 33818 11994
rect 33818 11942 33830 11994
rect 33830 11942 33844 11994
rect 33868 11942 33882 11994
rect 33882 11942 33894 11994
rect 33894 11942 33924 11994
rect 33948 11942 33958 11994
rect 33958 11942 34004 11994
rect 33708 11940 33764 11942
rect 33788 11940 33844 11942
rect 33868 11940 33924 11942
rect 33948 11940 34004 11942
rect 31482 11192 31538 11248
rect 33708 10906 33764 10908
rect 33788 10906 33844 10908
rect 33868 10906 33924 10908
rect 33948 10906 34004 10908
rect 33708 10854 33754 10906
rect 33754 10854 33764 10906
rect 33788 10854 33818 10906
rect 33818 10854 33830 10906
rect 33830 10854 33844 10906
rect 33868 10854 33882 10906
rect 33882 10854 33894 10906
rect 33894 10854 33924 10906
rect 33948 10854 33958 10906
rect 33958 10854 34004 10906
rect 33708 10852 33764 10854
rect 33788 10852 33844 10854
rect 33868 10852 33924 10854
rect 33948 10852 34004 10854
rect 29614 10362 29670 10364
rect 29694 10362 29750 10364
rect 29774 10362 29830 10364
rect 29854 10362 29910 10364
rect 29614 10310 29660 10362
rect 29660 10310 29670 10362
rect 29694 10310 29724 10362
rect 29724 10310 29736 10362
rect 29736 10310 29750 10362
rect 29774 10310 29788 10362
rect 29788 10310 29800 10362
rect 29800 10310 29830 10362
rect 29854 10310 29864 10362
rect 29864 10310 29910 10362
rect 29614 10308 29670 10310
rect 29694 10308 29750 10310
rect 29774 10308 29830 10310
rect 29854 10308 29910 10310
rect 29614 9274 29670 9276
rect 29694 9274 29750 9276
rect 29774 9274 29830 9276
rect 29854 9274 29910 9276
rect 29614 9222 29660 9274
rect 29660 9222 29670 9274
rect 29694 9222 29724 9274
rect 29724 9222 29736 9274
rect 29736 9222 29750 9274
rect 29774 9222 29788 9274
rect 29788 9222 29800 9274
rect 29800 9222 29830 9274
rect 29854 9222 29864 9274
rect 29864 9222 29910 9274
rect 29614 9220 29670 9222
rect 29694 9220 29750 9222
rect 29774 9220 29830 9222
rect 29854 9220 29910 9222
rect 29614 8186 29670 8188
rect 29694 8186 29750 8188
rect 29774 8186 29830 8188
rect 29854 8186 29910 8188
rect 29614 8134 29660 8186
rect 29660 8134 29670 8186
rect 29694 8134 29724 8186
rect 29724 8134 29736 8186
rect 29736 8134 29750 8186
rect 29774 8134 29788 8186
rect 29788 8134 29800 8186
rect 29800 8134 29830 8186
rect 29854 8134 29864 8186
rect 29864 8134 29910 8186
rect 29614 8132 29670 8134
rect 29694 8132 29750 8134
rect 29774 8132 29830 8134
rect 29854 8132 29910 8134
rect 26422 5752 26478 5808
rect 27526 5752 27582 5808
rect 26698 5652 26700 5672
rect 26700 5652 26752 5672
rect 26752 5652 26754 5672
rect 26698 5616 26754 5652
rect 25520 2202 25576 2204
rect 25600 2202 25656 2204
rect 25680 2202 25736 2204
rect 25760 2202 25816 2204
rect 25520 2150 25566 2202
rect 25566 2150 25576 2202
rect 25600 2150 25630 2202
rect 25630 2150 25642 2202
rect 25642 2150 25656 2202
rect 25680 2150 25694 2202
rect 25694 2150 25706 2202
rect 25706 2150 25736 2202
rect 25760 2150 25770 2202
rect 25770 2150 25816 2202
rect 25520 2148 25576 2150
rect 25600 2148 25656 2150
rect 25680 2148 25736 2150
rect 25760 2148 25816 2150
rect 29182 5244 29184 5264
rect 29184 5244 29236 5264
rect 29236 5244 29238 5264
rect 29182 5208 29238 5244
rect 29614 7098 29670 7100
rect 29694 7098 29750 7100
rect 29774 7098 29830 7100
rect 29854 7098 29910 7100
rect 29614 7046 29660 7098
rect 29660 7046 29670 7098
rect 29694 7046 29724 7098
rect 29724 7046 29736 7098
rect 29736 7046 29750 7098
rect 29774 7046 29788 7098
rect 29788 7046 29800 7098
rect 29800 7046 29830 7098
rect 29854 7046 29864 7098
rect 29864 7046 29910 7098
rect 29614 7044 29670 7046
rect 29694 7044 29750 7046
rect 29774 7044 29830 7046
rect 29854 7044 29910 7046
rect 29614 6010 29670 6012
rect 29694 6010 29750 6012
rect 29774 6010 29830 6012
rect 29854 6010 29910 6012
rect 29614 5958 29660 6010
rect 29660 5958 29670 6010
rect 29694 5958 29724 6010
rect 29724 5958 29736 6010
rect 29736 5958 29750 6010
rect 29774 5958 29788 6010
rect 29788 5958 29800 6010
rect 29800 5958 29830 6010
rect 29854 5958 29864 6010
rect 29864 5958 29910 6010
rect 29614 5956 29670 5958
rect 29694 5956 29750 5958
rect 29774 5956 29830 5958
rect 29854 5956 29910 5958
rect 33708 9818 33764 9820
rect 33788 9818 33844 9820
rect 33868 9818 33924 9820
rect 33948 9818 34004 9820
rect 33708 9766 33754 9818
rect 33754 9766 33764 9818
rect 33788 9766 33818 9818
rect 33818 9766 33830 9818
rect 33830 9766 33844 9818
rect 33868 9766 33882 9818
rect 33882 9766 33894 9818
rect 33894 9766 33924 9818
rect 33948 9766 33958 9818
rect 33958 9766 34004 9818
rect 33708 9764 33764 9766
rect 33788 9764 33844 9766
rect 33868 9764 33924 9766
rect 33948 9764 34004 9766
rect 33322 9560 33378 9616
rect 31298 8472 31354 8528
rect 33708 8730 33764 8732
rect 33788 8730 33844 8732
rect 33868 8730 33924 8732
rect 33948 8730 34004 8732
rect 33708 8678 33754 8730
rect 33754 8678 33764 8730
rect 33788 8678 33818 8730
rect 33818 8678 33830 8730
rect 33830 8678 33844 8730
rect 33868 8678 33882 8730
rect 33882 8678 33894 8730
rect 33894 8678 33924 8730
rect 33948 8678 33958 8730
rect 33958 8678 34004 8730
rect 33708 8676 33764 8678
rect 33788 8676 33844 8678
rect 33868 8676 33924 8678
rect 33948 8676 34004 8678
rect 30746 5752 30802 5808
rect 29614 4922 29670 4924
rect 29694 4922 29750 4924
rect 29774 4922 29830 4924
rect 29854 4922 29910 4924
rect 29614 4870 29660 4922
rect 29660 4870 29670 4922
rect 29694 4870 29724 4922
rect 29724 4870 29736 4922
rect 29736 4870 29750 4922
rect 29774 4870 29788 4922
rect 29788 4870 29800 4922
rect 29800 4870 29830 4922
rect 29854 4870 29864 4922
rect 29864 4870 29910 4922
rect 29614 4868 29670 4870
rect 29694 4868 29750 4870
rect 29774 4868 29830 4870
rect 29854 4868 29910 4870
rect 29614 3834 29670 3836
rect 29694 3834 29750 3836
rect 29774 3834 29830 3836
rect 29854 3834 29910 3836
rect 29614 3782 29660 3834
rect 29660 3782 29670 3834
rect 29694 3782 29724 3834
rect 29724 3782 29736 3834
rect 29736 3782 29750 3834
rect 29774 3782 29788 3834
rect 29788 3782 29800 3834
rect 29800 3782 29830 3834
rect 29854 3782 29864 3834
rect 29864 3782 29910 3834
rect 29614 3780 29670 3782
rect 29694 3780 29750 3782
rect 29774 3780 29830 3782
rect 29854 3780 29910 3782
rect 29614 2746 29670 2748
rect 29694 2746 29750 2748
rect 29774 2746 29830 2748
rect 29854 2746 29910 2748
rect 29614 2694 29660 2746
rect 29660 2694 29670 2746
rect 29694 2694 29724 2746
rect 29724 2694 29736 2746
rect 29736 2694 29750 2746
rect 29774 2694 29788 2746
rect 29788 2694 29800 2746
rect 29800 2694 29830 2746
rect 29854 2694 29864 2746
rect 29864 2694 29910 2746
rect 29614 2692 29670 2694
rect 29694 2692 29750 2694
rect 29774 2692 29830 2694
rect 29854 2692 29910 2694
rect 29550 1672 29606 1728
rect 33708 7642 33764 7644
rect 33788 7642 33844 7644
rect 33868 7642 33924 7644
rect 33948 7642 34004 7644
rect 33708 7590 33754 7642
rect 33754 7590 33764 7642
rect 33788 7590 33818 7642
rect 33818 7590 33830 7642
rect 33830 7590 33844 7642
rect 33868 7590 33882 7642
rect 33882 7590 33894 7642
rect 33894 7590 33924 7642
rect 33948 7590 33958 7642
rect 33958 7590 34004 7642
rect 33708 7588 33764 7590
rect 33788 7588 33844 7590
rect 33868 7588 33924 7590
rect 33948 7588 34004 7590
rect 33322 7112 33378 7168
rect 31482 5752 31538 5808
rect 31574 4528 31630 4584
rect 32218 4664 32274 4720
rect 33708 6554 33764 6556
rect 33788 6554 33844 6556
rect 33868 6554 33924 6556
rect 33948 6554 34004 6556
rect 33708 6502 33754 6554
rect 33754 6502 33764 6554
rect 33788 6502 33818 6554
rect 33818 6502 33830 6554
rect 33830 6502 33844 6554
rect 33868 6502 33882 6554
rect 33882 6502 33894 6554
rect 33894 6502 33924 6554
rect 33948 6502 33958 6554
rect 33958 6502 34004 6554
rect 33708 6500 33764 6502
rect 33788 6500 33844 6502
rect 33868 6500 33924 6502
rect 33948 6500 34004 6502
rect 33506 5616 33562 5672
rect 33708 5466 33764 5468
rect 33788 5466 33844 5468
rect 33868 5466 33924 5468
rect 33948 5466 34004 5468
rect 33708 5414 33754 5466
rect 33754 5414 33764 5466
rect 33788 5414 33818 5466
rect 33818 5414 33830 5466
rect 33830 5414 33844 5466
rect 33868 5414 33882 5466
rect 33882 5414 33894 5466
rect 33894 5414 33924 5466
rect 33948 5414 33958 5466
rect 33958 5414 34004 5466
rect 33708 5412 33764 5414
rect 33788 5412 33844 5414
rect 33868 5412 33924 5414
rect 33948 5412 34004 5414
rect 33708 4378 33764 4380
rect 33788 4378 33844 4380
rect 33868 4378 33924 4380
rect 33948 4378 34004 4380
rect 33708 4326 33754 4378
rect 33754 4326 33764 4378
rect 33788 4326 33818 4378
rect 33818 4326 33830 4378
rect 33830 4326 33844 4378
rect 33868 4326 33882 4378
rect 33882 4326 33894 4378
rect 33894 4326 33924 4378
rect 33948 4326 33958 4378
rect 33958 4326 34004 4378
rect 33708 4324 33764 4326
rect 33788 4324 33844 4326
rect 33868 4324 33924 4326
rect 33948 4324 34004 4326
rect 33708 3290 33764 3292
rect 33788 3290 33844 3292
rect 33868 3290 33924 3292
rect 33948 3290 34004 3292
rect 33708 3238 33754 3290
rect 33754 3238 33764 3290
rect 33788 3238 33818 3290
rect 33818 3238 33830 3290
rect 33830 3238 33844 3290
rect 33868 3238 33882 3290
rect 33882 3238 33894 3290
rect 33894 3238 33924 3290
rect 33948 3238 33958 3290
rect 33958 3238 34004 3290
rect 33708 3236 33764 3238
rect 33788 3236 33844 3238
rect 33868 3236 33924 3238
rect 33948 3236 34004 3238
rect 33506 3032 33562 3088
rect 33708 2202 33764 2204
rect 33788 2202 33844 2204
rect 33868 2202 33924 2204
rect 33948 2202 34004 2204
rect 33708 2150 33754 2202
rect 33754 2150 33764 2202
rect 33788 2150 33818 2202
rect 33818 2150 33830 2202
rect 33830 2150 33844 2202
rect 33868 2150 33882 2202
rect 33882 2150 33894 2202
rect 33894 2150 33924 2202
rect 33948 2150 33958 2202
rect 33958 2150 34004 2202
rect 33708 2148 33764 2150
rect 33788 2148 33844 2150
rect 33868 2148 33924 2150
rect 33948 2148 34004 2150
<< metal3 >>
rect 31293 33010 31359 33013
rect 34200 33010 35000 33040
rect 31293 33008 35000 33010
rect 31293 32952 31298 33008
rect 31354 32952 35000 33008
rect 31293 32950 35000 32952
rect 31293 32947 31359 32950
rect 34200 32920 35000 32950
rect 9134 32672 9450 32673
rect 9134 32608 9140 32672
rect 9204 32608 9220 32672
rect 9284 32608 9300 32672
rect 9364 32608 9380 32672
rect 9444 32608 9450 32672
rect 9134 32607 9450 32608
rect 17322 32672 17638 32673
rect 17322 32608 17328 32672
rect 17392 32608 17408 32672
rect 17472 32608 17488 32672
rect 17552 32608 17568 32672
rect 17632 32608 17638 32672
rect 17322 32607 17638 32608
rect 25510 32672 25826 32673
rect 25510 32608 25516 32672
rect 25580 32608 25596 32672
rect 25660 32608 25676 32672
rect 25740 32608 25756 32672
rect 25820 32608 25826 32672
rect 25510 32607 25826 32608
rect 33698 32672 34014 32673
rect 33698 32608 33704 32672
rect 33768 32608 33784 32672
rect 33848 32608 33864 32672
rect 33928 32608 33944 32672
rect 34008 32608 34014 32672
rect 33698 32607 34014 32608
rect 5040 32128 5356 32129
rect 5040 32064 5046 32128
rect 5110 32064 5126 32128
rect 5190 32064 5206 32128
rect 5270 32064 5286 32128
rect 5350 32064 5356 32128
rect 5040 32063 5356 32064
rect 13228 32128 13544 32129
rect 13228 32064 13234 32128
rect 13298 32064 13314 32128
rect 13378 32064 13394 32128
rect 13458 32064 13474 32128
rect 13538 32064 13544 32128
rect 13228 32063 13544 32064
rect 21416 32128 21732 32129
rect 21416 32064 21422 32128
rect 21486 32064 21502 32128
rect 21566 32064 21582 32128
rect 21646 32064 21662 32128
rect 21726 32064 21732 32128
rect 21416 32063 21732 32064
rect 29604 32128 29920 32129
rect 29604 32064 29610 32128
rect 29674 32064 29690 32128
rect 29754 32064 29770 32128
rect 29834 32064 29850 32128
rect 29914 32064 29920 32128
rect 29604 32063 29920 32064
rect 28950 31726 34162 31786
rect 0 31650 800 31680
rect 4061 31650 4127 31653
rect 0 31648 4127 31650
rect 0 31592 4066 31648
rect 4122 31592 4127 31648
rect 0 31590 4127 31592
rect 0 31560 800 31590
rect 4061 31587 4127 31590
rect 9134 31584 9450 31585
rect 9134 31520 9140 31584
rect 9204 31520 9220 31584
rect 9284 31520 9300 31584
rect 9364 31520 9380 31584
rect 9444 31520 9450 31584
rect 9134 31519 9450 31520
rect 17322 31584 17638 31585
rect 17322 31520 17328 31584
rect 17392 31520 17408 31584
rect 17472 31520 17488 31584
rect 17552 31520 17568 31584
rect 17632 31520 17638 31584
rect 17322 31519 17638 31520
rect 25510 31584 25826 31585
rect 25510 31520 25516 31584
rect 25580 31520 25596 31584
rect 25660 31520 25676 31584
rect 25740 31520 25756 31584
rect 25820 31520 25826 31584
rect 25510 31519 25826 31520
rect 27429 31378 27495 31381
rect 28950 31378 29010 31726
rect 34102 31684 34162 31726
rect 34102 31680 34346 31684
rect 34102 31624 35000 31680
rect 33698 31584 34014 31585
rect 33698 31520 33704 31584
rect 33768 31520 33784 31584
rect 33848 31520 33864 31584
rect 33928 31520 33944 31584
rect 34008 31520 34014 31584
rect 34200 31560 35000 31624
rect 33698 31519 34014 31520
rect 27429 31376 29010 31378
rect 27429 31320 27434 31376
rect 27490 31320 29010 31376
rect 27429 31318 29010 31320
rect 27429 31315 27495 31318
rect 5040 31040 5356 31041
rect 5040 30976 5046 31040
rect 5110 30976 5126 31040
rect 5190 30976 5206 31040
rect 5270 30976 5286 31040
rect 5350 30976 5356 31040
rect 5040 30975 5356 30976
rect 13228 31040 13544 31041
rect 13228 30976 13234 31040
rect 13298 30976 13314 31040
rect 13378 30976 13394 31040
rect 13458 30976 13474 31040
rect 13538 30976 13544 31040
rect 13228 30975 13544 30976
rect 21416 31040 21732 31041
rect 21416 30976 21422 31040
rect 21486 30976 21502 31040
rect 21566 30976 21582 31040
rect 21646 30976 21662 31040
rect 21726 30976 21732 31040
rect 21416 30975 21732 30976
rect 29604 31040 29920 31041
rect 29604 30976 29610 31040
rect 29674 30976 29690 31040
rect 29754 30976 29770 31040
rect 29834 30976 29850 31040
rect 29914 30976 29920 31040
rect 29604 30975 29920 30976
rect 9134 30496 9450 30497
rect 9134 30432 9140 30496
rect 9204 30432 9220 30496
rect 9284 30432 9300 30496
rect 9364 30432 9380 30496
rect 9444 30432 9450 30496
rect 9134 30431 9450 30432
rect 17322 30496 17638 30497
rect 17322 30432 17328 30496
rect 17392 30432 17408 30496
rect 17472 30432 17488 30496
rect 17552 30432 17568 30496
rect 17632 30432 17638 30496
rect 17322 30431 17638 30432
rect 25510 30496 25826 30497
rect 25510 30432 25516 30496
rect 25580 30432 25596 30496
rect 25660 30432 25676 30496
rect 25740 30432 25756 30496
rect 25820 30432 25826 30496
rect 25510 30431 25826 30432
rect 33698 30496 34014 30497
rect 33698 30432 33704 30496
rect 33768 30432 33784 30496
rect 33848 30432 33864 30496
rect 33928 30432 33944 30496
rect 34008 30432 34014 30496
rect 33698 30431 34014 30432
rect 0 30290 800 30320
rect 1393 30290 1459 30293
rect 0 30288 1459 30290
rect 0 30232 1398 30288
rect 1454 30232 1459 30288
rect 0 30230 1459 30232
rect 0 30200 800 30230
rect 1393 30227 1459 30230
rect 32949 30290 33015 30293
rect 34200 30290 35000 30320
rect 32949 30288 35000 30290
rect 32949 30232 32954 30288
rect 33010 30232 35000 30288
rect 32949 30230 35000 30232
rect 32949 30227 33015 30230
rect 34200 30200 35000 30230
rect 5040 29952 5356 29953
rect 5040 29888 5046 29952
rect 5110 29888 5126 29952
rect 5190 29888 5206 29952
rect 5270 29888 5286 29952
rect 5350 29888 5356 29952
rect 5040 29887 5356 29888
rect 13228 29952 13544 29953
rect 13228 29888 13234 29952
rect 13298 29888 13314 29952
rect 13378 29888 13394 29952
rect 13458 29888 13474 29952
rect 13538 29888 13544 29952
rect 13228 29887 13544 29888
rect 21416 29952 21732 29953
rect 21416 29888 21422 29952
rect 21486 29888 21502 29952
rect 21566 29888 21582 29952
rect 21646 29888 21662 29952
rect 21726 29888 21732 29952
rect 21416 29887 21732 29888
rect 29604 29952 29920 29953
rect 29604 29888 29610 29952
rect 29674 29888 29690 29952
rect 29754 29888 29770 29952
rect 29834 29888 29850 29952
rect 29914 29888 29920 29952
rect 29604 29887 29920 29888
rect 9134 29408 9450 29409
rect 9134 29344 9140 29408
rect 9204 29344 9220 29408
rect 9284 29344 9300 29408
rect 9364 29344 9380 29408
rect 9444 29344 9450 29408
rect 9134 29343 9450 29344
rect 17322 29408 17638 29409
rect 17322 29344 17328 29408
rect 17392 29344 17408 29408
rect 17472 29344 17488 29408
rect 17552 29344 17568 29408
rect 17632 29344 17638 29408
rect 17322 29343 17638 29344
rect 25510 29408 25826 29409
rect 25510 29344 25516 29408
rect 25580 29344 25596 29408
rect 25660 29344 25676 29408
rect 25740 29344 25756 29408
rect 25820 29344 25826 29408
rect 25510 29343 25826 29344
rect 33698 29408 34014 29409
rect 33698 29344 33704 29408
rect 33768 29344 33784 29408
rect 33848 29344 33864 29408
rect 33928 29344 33944 29408
rect 34008 29344 34014 29408
rect 33698 29343 34014 29344
rect 0 28930 800 28960
rect 3325 28930 3391 28933
rect 0 28928 3391 28930
rect 0 28872 3330 28928
rect 3386 28872 3391 28928
rect 0 28870 3391 28872
rect 0 28840 800 28870
rect 3325 28867 3391 28870
rect 31477 28930 31543 28933
rect 34200 28930 35000 28960
rect 31477 28928 35000 28930
rect 31477 28872 31482 28928
rect 31538 28872 35000 28928
rect 31477 28870 35000 28872
rect 31477 28867 31543 28870
rect 5040 28864 5356 28865
rect 5040 28800 5046 28864
rect 5110 28800 5126 28864
rect 5190 28800 5206 28864
rect 5270 28800 5286 28864
rect 5350 28800 5356 28864
rect 5040 28799 5356 28800
rect 13228 28864 13544 28865
rect 13228 28800 13234 28864
rect 13298 28800 13314 28864
rect 13378 28800 13394 28864
rect 13458 28800 13474 28864
rect 13538 28800 13544 28864
rect 13228 28799 13544 28800
rect 21416 28864 21732 28865
rect 21416 28800 21422 28864
rect 21486 28800 21502 28864
rect 21566 28800 21582 28864
rect 21646 28800 21662 28864
rect 21726 28800 21732 28864
rect 21416 28799 21732 28800
rect 29604 28864 29920 28865
rect 29604 28800 29610 28864
rect 29674 28800 29690 28864
rect 29754 28800 29770 28864
rect 29834 28800 29850 28864
rect 29914 28800 29920 28864
rect 34200 28840 35000 28870
rect 29604 28799 29920 28800
rect 9134 28320 9450 28321
rect 9134 28256 9140 28320
rect 9204 28256 9220 28320
rect 9284 28256 9300 28320
rect 9364 28256 9380 28320
rect 9444 28256 9450 28320
rect 9134 28255 9450 28256
rect 17322 28320 17638 28321
rect 17322 28256 17328 28320
rect 17392 28256 17408 28320
rect 17472 28256 17488 28320
rect 17552 28256 17568 28320
rect 17632 28256 17638 28320
rect 17322 28255 17638 28256
rect 25510 28320 25826 28321
rect 25510 28256 25516 28320
rect 25580 28256 25596 28320
rect 25660 28256 25676 28320
rect 25740 28256 25756 28320
rect 25820 28256 25826 28320
rect 25510 28255 25826 28256
rect 33698 28320 34014 28321
rect 33698 28256 33704 28320
rect 33768 28256 33784 28320
rect 33848 28256 33864 28320
rect 33928 28256 33944 28320
rect 34008 28256 34014 28320
rect 33698 28255 34014 28256
rect 5040 27776 5356 27777
rect 5040 27712 5046 27776
rect 5110 27712 5126 27776
rect 5190 27712 5206 27776
rect 5270 27712 5286 27776
rect 5350 27712 5356 27776
rect 5040 27711 5356 27712
rect 13228 27776 13544 27777
rect 13228 27712 13234 27776
rect 13298 27712 13314 27776
rect 13378 27712 13394 27776
rect 13458 27712 13474 27776
rect 13538 27712 13544 27776
rect 13228 27711 13544 27712
rect 21416 27776 21732 27777
rect 21416 27712 21422 27776
rect 21486 27712 21502 27776
rect 21566 27712 21582 27776
rect 21646 27712 21662 27776
rect 21726 27712 21732 27776
rect 21416 27711 21732 27712
rect 29604 27776 29920 27777
rect 29604 27712 29610 27776
rect 29674 27712 29690 27776
rect 29754 27712 29770 27776
rect 29834 27712 29850 27776
rect 29914 27712 29920 27776
rect 29604 27711 29920 27712
rect 0 27570 800 27600
rect 2773 27570 2839 27573
rect 0 27568 2839 27570
rect 0 27512 2778 27568
rect 2834 27512 2839 27568
rect 0 27510 2839 27512
rect 0 27480 800 27510
rect 2773 27507 2839 27510
rect 31477 27570 31543 27573
rect 34200 27570 35000 27600
rect 31477 27568 35000 27570
rect 31477 27512 31482 27568
rect 31538 27512 35000 27568
rect 31477 27510 35000 27512
rect 31477 27507 31543 27510
rect 34200 27480 35000 27510
rect 9134 27232 9450 27233
rect 9134 27168 9140 27232
rect 9204 27168 9220 27232
rect 9284 27168 9300 27232
rect 9364 27168 9380 27232
rect 9444 27168 9450 27232
rect 9134 27167 9450 27168
rect 17322 27232 17638 27233
rect 17322 27168 17328 27232
rect 17392 27168 17408 27232
rect 17472 27168 17488 27232
rect 17552 27168 17568 27232
rect 17632 27168 17638 27232
rect 17322 27167 17638 27168
rect 25510 27232 25826 27233
rect 25510 27168 25516 27232
rect 25580 27168 25596 27232
rect 25660 27168 25676 27232
rect 25740 27168 25756 27232
rect 25820 27168 25826 27232
rect 25510 27167 25826 27168
rect 33698 27232 34014 27233
rect 33698 27168 33704 27232
rect 33768 27168 33784 27232
rect 33848 27168 33864 27232
rect 33928 27168 33944 27232
rect 34008 27168 34014 27232
rect 33698 27167 34014 27168
rect 5040 26688 5356 26689
rect 5040 26624 5046 26688
rect 5110 26624 5126 26688
rect 5190 26624 5206 26688
rect 5270 26624 5286 26688
rect 5350 26624 5356 26688
rect 5040 26623 5356 26624
rect 13228 26688 13544 26689
rect 13228 26624 13234 26688
rect 13298 26624 13314 26688
rect 13378 26624 13394 26688
rect 13458 26624 13474 26688
rect 13538 26624 13544 26688
rect 13228 26623 13544 26624
rect 21416 26688 21732 26689
rect 21416 26624 21422 26688
rect 21486 26624 21502 26688
rect 21566 26624 21582 26688
rect 21646 26624 21662 26688
rect 21726 26624 21732 26688
rect 21416 26623 21732 26624
rect 29604 26688 29920 26689
rect 29604 26624 29610 26688
rect 29674 26624 29690 26688
rect 29754 26624 29770 26688
rect 29834 26624 29850 26688
rect 29914 26624 29920 26688
rect 29604 26623 29920 26624
rect 33317 26346 33383 26349
rect 33317 26344 34162 26346
rect 33317 26288 33322 26344
rect 33378 26288 34162 26344
rect 33317 26286 34162 26288
rect 33317 26283 33383 26286
rect 34102 26244 34162 26286
rect 34102 26240 34346 26244
rect 0 26210 800 26240
rect 1577 26210 1643 26213
rect 0 26208 1643 26210
rect 0 26152 1582 26208
rect 1638 26152 1643 26208
rect 34102 26184 35000 26240
rect 0 26150 1643 26152
rect 0 26120 800 26150
rect 1577 26147 1643 26150
rect 9134 26144 9450 26145
rect 9134 26080 9140 26144
rect 9204 26080 9220 26144
rect 9284 26080 9300 26144
rect 9364 26080 9380 26144
rect 9444 26080 9450 26144
rect 9134 26079 9450 26080
rect 17322 26144 17638 26145
rect 17322 26080 17328 26144
rect 17392 26080 17408 26144
rect 17472 26080 17488 26144
rect 17552 26080 17568 26144
rect 17632 26080 17638 26144
rect 17322 26079 17638 26080
rect 25510 26144 25826 26145
rect 25510 26080 25516 26144
rect 25580 26080 25596 26144
rect 25660 26080 25676 26144
rect 25740 26080 25756 26144
rect 25820 26080 25826 26144
rect 25510 26079 25826 26080
rect 33698 26144 34014 26145
rect 33698 26080 33704 26144
rect 33768 26080 33784 26144
rect 33848 26080 33864 26144
rect 33928 26080 33944 26144
rect 34008 26080 34014 26144
rect 34200 26120 35000 26184
rect 33698 26079 34014 26080
rect 5040 25600 5356 25601
rect 5040 25536 5046 25600
rect 5110 25536 5126 25600
rect 5190 25536 5206 25600
rect 5270 25536 5286 25600
rect 5350 25536 5356 25600
rect 5040 25535 5356 25536
rect 13228 25600 13544 25601
rect 13228 25536 13234 25600
rect 13298 25536 13314 25600
rect 13378 25536 13394 25600
rect 13458 25536 13474 25600
rect 13538 25536 13544 25600
rect 13228 25535 13544 25536
rect 21416 25600 21732 25601
rect 21416 25536 21422 25600
rect 21486 25536 21502 25600
rect 21566 25536 21582 25600
rect 21646 25536 21662 25600
rect 21726 25536 21732 25600
rect 21416 25535 21732 25536
rect 29604 25600 29920 25601
rect 29604 25536 29610 25600
rect 29674 25536 29690 25600
rect 29754 25536 29770 25600
rect 29834 25536 29850 25600
rect 29914 25536 29920 25600
rect 29604 25535 29920 25536
rect 9134 25056 9450 25057
rect 9134 24992 9140 25056
rect 9204 24992 9220 25056
rect 9284 24992 9300 25056
rect 9364 24992 9380 25056
rect 9444 24992 9450 25056
rect 9134 24991 9450 24992
rect 17322 25056 17638 25057
rect 17322 24992 17328 25056
rect 17392 24992 17408 25056
rect 17472 24992 17488 25056
rect 17552 24992 17568 25056
rect 17632 24992 17638 25056
rect 17322 24991 17638 24992
rect 25510 25056 25826 25057
rect 25510 24992 25516 25056
rect 25580 24992 25596 25056
rect 25660 24992 25676 25056
rect 25740 24992 25756 25056
rect 25820 24992 25826 25056
rect 25510 24991 25826 24992
rect 33698 25056 34014 25057
rect 33698 24992 33704 25056
rect 33768 24992 33784 25056
rect 33848 24992 33864 25056
rect 33928 24992 33944 25056
rect 34008 24992 34014 25056
rect 33698 24991 34014 24992
rect 0 24850 800 24880
rect 2773 24850 2839 24853
rect 0 24848 2839 24850
rect 0 24792 2778 24848
rect 2834 24792 2839 24848
rect 0 24790 2839 24792
rect 0 24760 800 24790
rect 2773 24787 2839 24790
rect 31109 24850 31175 24853
rect 34200 24850 35000 24880
rect 31109 24848 35000 24850
rect 31109 24792 31114 24848
rect 31170 24792 35000 24848
rect 31109 24790 35000 24792
rect 31109 24787 31175 24790
rect 34200 24760 35000 24790
rect 5040 24512 5356 24513
rect 5040 24448 5046 24512
rect 5110 24448 5126 24512
rect 5190 24448 5206 24512
rect 5270 24448 5286 24512
rect 5350 24448 5356 24512
rect 5040 24447 5356 24448
rect 13228 24512 13544 24513
rect 13228 24448 13234 24512
rect 13298 24448 13314 24512
rect 13378 24448 13394 24512
rect 13458 24448 13474 24512
rect 13538 24448 13544 24512
rect 13228 24447 13544 24448
rect 21416 24512 21732 24513
rect 21416 24448 21422 24512
rect 21486 24448 21502 24512
rect 21566 24448 21582 24512
rect 21646 24448 21662 24512
rect 21726 24448 21732 24512
rect 21416 24447 21732 24448
rect 29604 24512 29920 24513
rect 29604 24448 29610 24512
rect 29674 24448 29690 24512
rect 29754 24448 29770 24512
rect 29834 24448 29850 24512
rect 29914 24448 29920 24512
rect 29604 24447 29920 24448
rect 9134 23968 9450 23969
rect 9134 23904 9140 23968
rect 9204 23904 9220 23968
rect 9284 23904 9300 23968
rect 9364 23904 9380 23968
rect 9444 23904 9450 23968
rect 9134 23903 9450 23904
rect 17322 23968 17638 23969
rect 17322 23904 17328 23968
rect 17392 23904 17408 23968
rect 17472 23904 17488 23968
rect 17552 23904 17568 23968
rect 17632 23904 17638 23968
rect 17322 23903 17638 23904
rect 25510 23968 25826 23969
rect 25510 23904 25516 23968
rect 25580 23904 25596 23968
rect 25660 23904 25676 23968
rect 25740 23904 25756 23968
rect 25820 23904 25826 23968
rect 25510 23903 25826 23904
rect 33698 23968 34014 23969
rect 33698 23904 33704 23968
rect 33768 23904 33784 23968
rect 33848 23904 33864 23968
rect 33928 23904 33944 23968
rect 34008 23904 34014 23968
rect 33698 23903 34014 23904
rect 0 23490 800 23520
rect 933 23490 999 23493
rect 0 23488 999 23490
rect 0 23432 938 23488
rect 994 23432 999 23488
rect 0 23430 999 23432
rect 0 23400 800 23430
rect 933 23427 999 23430
rect 33777 23490 33843 23493
rect 34200 23490 35000 23520
rect 33777 23488 35000 23490
rect 33777 23432 33782 23488
rect 33838 23432 35000 23488
rect 33777 23430 35000 23432
rect 33777 23427 33843 23430
rect 5040 23424 5356 23425
rect 5040 23360 5046 23424
rect 5110 23360 5126 23424
rect 5190 23360 5206 23424
rect 5270 23360 5286 23424
rect 5350 23360 5356 23424
rect 5040 23359 5356 23360
rect 13228 23424 13544 23425
rect 13228 23360 13234 23424
rect 13298 23360 13314 23424
rect 13378 23360 13394 23424
rect 13458 23360 13474 23424
rect 13538 23360 13544 23424
rect 13228 23359 13544 23360
rect 21416 23424 21732 23425
rect 21416 23360 21422 23424
rect 21486 23360 21502 23424
rect 21566 23360 21582 23424
rect 21646 23360 21662 23424
rect 21726 23360 21732 23424
rect 21416 23359 21732 23360
rect 29604 23424 29920 23425
rect 29604 23360 29610 23424
rect 29674 23360 29690 23424
rect 29754 23360 29770 23424
rect 29834 23360 29850 23424
rect 29914 23360 29920 23424
rect 34200 23400 35000 23430
rect 29604 23359 29920 23360
rect 9134 22880 9450 22881
rect 9134 22816 9140 22880
rect 9204 22816 9220 22880
rect 9284 22816 9300 22880
rect 9364 22816 9380 22880
rect 9444 22816 9450 22880
rect 9134 22815 9450 22816
rect 17322 22880 17638 22881
rect 17322 22816 17328 22880
rect 17392 22816 17408 22880
rect 17472 22816 17488 22880
rect 17552 22816 17568 22880
rect 17632 22816 17638 22880
rect 17322 22815 17638 22816
rect 25510 22880 25826 22881
rect 25510 22816 25516 22880
rect 25580 22816 25596 22880
rect 25660 22816 25676 22880
rect 25740 22816 25756 22880
rect 25820 22816 25826 22880
rect 25510 22815 25826 22816
rect 33698 22880 34014 22881
rect 33698 22816 33704 22880
rect 33768 22816 33784 22880
rect 33848 22816 33864 22880
rect 33928 22816 33944 22880
rect 34008 22816 34014 22880
rect 33698 22815 34014 22816
rect 1577 22402 1643 22405
rect 982 22400 1643 22402
rect 982 22344 1582 22400
rect 1638 22344 1643 22400
rect 982 22342 1643 22344
rect 0 22130 800 22160
rect 982 22130 1042 22342
rect 1577 22339 1643 22342
rect 5040 22336 5356 22337
rect 5040 22272 5046 22336
rect 5110 22272 5126 22336
rect 5190 22272 5206 22336
rect 5270 22272 5286 22336
rect 5350 22272 5356 22336
rect 5040 22271 5356 22272
rect 13228 22336 13544 22337
rect 13228 22272 13234 22336
rect 13298 22272 13314 22336
rect 13378 22272 13394 22336
rect 13458 22272 13474 22336
rect 13538 22272 13544 22336
rect 13228 22271 13544 22272
rect 21416 22336 21732 22337
rect 21416 22272 21422 22336
rect 21486 22272 21502 22336
rect 21566 22272 21582 22336
rect 21646 22272 21662 22336
rect 21726 22272 21732 22336
rect 21416 22271 21732 22272
rect 29604 22336 29920 22337
rect 29604 22272 29610 22336
rect 29674 22272 29690 22336
rect 29754 22272 29770 22336
rect 29834 22272 29850 22336
rect 29914 22272 29920 22336
rect 29604 22271 29920 22272
rect 0 22070 1042 22130
rect 31477 22130 31543 22133
rect 34200 22130 35000 22160
rect 31477 22128 35000 22130
rect 31477 22072 31482 22128
rect 31538 22072 35000 22128
rect 31477 22070 35000 22072
rect 0 22040 800 22070
rect 31477 22067 31543 22070
rect 34200 22040 35000 22070
rect 9134 21792 9450 21793
rect 9134 21728 9140 21792
rect 9204 21728 9220 21792
rect 9284 21728 9300 21792
rect 9364 21728 9380 21792
rect 9444 21728 9450 21792
rect 9134 21727 9450 21728
rect 17322 21792 17638 21793
rect 17322 21728 17328 21792
rect 17392 21728 17408 21792
rect 17472 21728 17488 21792
rect 17552 21728 17568 21792
rect 17632 21728 17638 21792
rect 17322 21727 17638 21728
rect 25510 21792 25826 21793
rect 25510 21728 25516 21792
rect 25580 21728 25596 21792
rect 25660 21728 25676 21792
rect 25740 21728 25756 21792
rect 25820 21728 25826 21792
rect 25510 21727 25826 21728
rect 33698 21792 34014 21793
rect 33698 21728 33704 21792
rect 33768 21728 33784 21792
rect 33848 21728 33864 21792
rect 33928 21728 33944 21792
rect 34008 21728 34014 21792
rect 33698 21727 34014 21728
rect 5040 21248 5356 21249
rect 5040 21184 5046 21248
rect 5110 21184 5126 21248
rect 5190 21184 5206 21248
rect 5270 21184 5286 21248
rect 5350 21184 5356 21248
rect 5040 21183 5356 21184
rect 13228 21248 13544 21249
rect 13228 21184 13234 21248
rect 13298 21184 13314 21248
rect 13378 21184 13394 21248
rect 13458 21184 13474 21248
rect 13538 21184 13544 21248
rect 13228 21183 13544 21184
rect 21416 21248 21732 21249
rect 21416 21184 21422 21248
rect 21486 21184 21502 21248
rect 21566 21184 21582 21248
rect 21646 21184 21662 21248
rect 21726 21184 21732 21248
rect 21416 21183 21732 21184
rect 29604 21248 29920 21249
rect 29604 21184 29610 21248
rect 29674 21184 29690 21248
rect 29754 21184 29770 21248
rect 29834 21184 29850 21248
rect 29914 21184 29920 21248
rect 29604 21183 29920 21184
rect 33317 20906 33383 20909
rect 33317 20904 34162 20906
rect 33317 20848 33322 20904
rect 33378 20848 34162 20904
rect 33317 20846 34162 20848
rect 33317 20843 33383 20846
rect 34102 20804 34162 20846
rect 34102 20800 34346 20804
rect 0 20770 800 20800
rect 933 20770 999 20773
rect 0 20768 999 20770
rect 0 20712 938 20768
rect 994 20712 999 20768
rect 34102 20744 35000 20800
rect 0 20710 999 20712
rect 0 20680 800 20710
rect 933 20707 999 20710
rect 9134 20704 9450 20705
rect 9134 20640 9140 20704
rect 9204 20640 9220 20704
rect 9284 20640 9300 20704
rect 9364 20640 9380 20704
rect 9444 20640 9450 20704
rect 9134 20639 9450 20640
rect 17322 20704 17638 20705
rect 17322 20640 17328 20704
rect 17392 20640 17408 20704
rect 17472 20640 17488 20704
rect 17552 20640 17568 20704
rect 17632 20640 17638 20704
rect 17322 20639 17638 20640
rect 25510 20704 25826 20705
rect 25510 20640 25516 20704
rect 25580 20640 25596 20704
rect 25660 20640 25676 20704
rect 25740 20640 25756 20704
rect 25820 20640 25826 20704
rect 25510 20639 25826 20640
rect 33698 20704 34014 20705
rect 33698 20640 33704 20704
rect 33768 20640 33784 20704
rect 33848 20640 33864 20704
rect 33928 20640 33944 20704
rect 34008 20640 34014 20704
rect 34200 20680 35000 20744
rect 33698 20639 34014 20640
rect 5040 20160 5356 20161
rect 5040 20096 5046 20160
rect 5110 20096 5126 20160
rect 5190 20096 5206 20160
rect 5270 20096 5286 20160
rect 5350 20096 5356 20160
rect 5040 20095 5356 20096
rect 13228 20160 13544 20161
rect 13228 20096 13234 20160
rect 13298 20096 13314 20160
rect 13378 20096 13394 20160
rect 13458 20096 13474 20160
rect 13538 20096 13544 20160
rect 13228 20095 13544 20096
rect 21416 20160 21732 20161
rect 21416 20096 21422 20160
rect 21486 20096 21502 20160
rect 21566 20096 21582 20160
rect 21646 20096 21662 20160
rect 21726 20096 21732 20160
rect 21416 20095 21732 20096
rect 29604 20160 29920 20161
rect 29604 20096 29610 20160
rect 29674 20096 29690 20160
rect 29754 20096 29770 20160
rect 29834 20096 29850 20160
rect 29914 20096 29920 20160
rect 29604 20095 29920 20096
rect 9134 19616 9450 19617
rect 9134 19552 9140 19616
rect 9204 19552 9220 19616
rect 9284 19552 9300 19616
rect 9364 19552 9380 19616
rect 9444 19552 9450 19616
rect 9134 19551 9450 19552
rect 17322 19616 17638 19617
rect 17322 19552 17328 19616
rect 17392 19552 17408 19616
rect 17472 19552 17488 19616
rect 17552 19552 17568 19616
rect 17632 19552 17638 19616
rect 17322 19551 17638 19552
rect 25510 19616 25826 19617
rect 25510 19552 25516 19616
rect 25580 19552 25596 19616
rect 25660 19552 25676 19616
rect 25740 19552 25756 19616
rect 25820 19552 25826 19616
rect 25510 19551 25826 19552
rect 33698 19616 34014 19617
rect 33698 19552 33704 19616
rect 33768 19552 33784 19616
rect 33848 19552 33864 19616
rect 33928 19552 33944 19616
rect 34008 19552 34014 19616
rect 33698 19551 34014 19552
rect 0 19410 800 19440
rect 933 19410 999 19413
rect 0 19408 999 19410
rect 0 19352 938 19408
rect 994 19352 999 19408
rect 0 19350 999 19352
rect 0 19320 800 19350
rect 933 19347 999 19350
rect 33317 19410 33383 19413
rect 34200 19410 35000 19440
rect 33317 19408 35000 19410
rect 33317 19352 33322 19408
rect 33378 19352 35000 19408
rect 33317 19350 35000 19352
rect 33317 19347 33383 19350
rect 34200 19320 35000 19350
rect 5040 19072 5356 19073
rect 5040 19008 5046 19072
rect 5110 19008 5126 19072
rect 5190 19008 5206 19072
rect 5270 19008 5286 19072
rect 5350 19008 5356 19072
rect 5040 19007 5356 19008
rect 13228 19072 13544 19073
rect 13228 19008 13234 19072
rect 13298 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13544 19072
rect 13228 19007 13544 19008
rect 21416 19072 21732 19073
rect 21416 19008 21422 19072
rect 21486 19008 21502 19072
rect 21566 19008 21582 19072
rect 21646 19008 21662 19072
rect 21726 19008 21732 19072
rect 21416 19007 21732 19008
rect 29604 19072 29920 19073
rect 29604 19008 29610 19072
rect 29674 19008 29690 19072
rect 29754 19008 29770 19072
rect 29834 19008 29850 19072
rect 29914 19008 29920 19072
rect 29604 19007 29920 19008
rect 9134 18528 9450 18529
rect 9134 18464 9140 18528
rect 9204 18464 9220 18528
rect 9284 18464 9300 18528
rect 9364 18464 9380 18528
rect 9444 18464 9450 18528
rect 9134 18463 9450 18464
rect 17322 18528 17638 18529
rect 17322 18464 17328 18528
rect 17392 18464 17408 18528
rect 17472 18464 17488 18528
rect 17552 18464 17568 18528
rect 17632 18464 17638 18528
rect 17322 18463 17638 18464
rect 25510 18528 25826 18529
rect 25510 18464 25516 18528
rect 25580 18464 25596 18528
rect 25660 18464 25676 18528
rect 25740 18464 25756 18528
rect 25820 18464 25826 18528
rect 25510 18463 25826 18464
rect 33698 18528 34014 18529
rect 33698 18464 33704 18528
rect 33768 18464 33784 18528
rect 33848 18464 33864 18528
rect 33928 18464 33944 18528
rect 34008 18464 34014 18528
rect 33698 18463 34014 18464
rect 0 18050 800 18080
rect 1301 18050 1367 18053
rect 0 18048 1367 18050
rect 0 17992 1306 18048
rect 1362 17992 1367 18048
rect 0 17990 1367 17992
rect 0 17960 800 17990
rect 1301 17987 1367 17990
rect 33317 18050 33383 18053
rect 34200 18050 35000 18080
rect 33317 18048 35000 18050
rect 33317 17992 33322 18048
rect 33378 17992 35000 18048
rect 33317 17990 35000 17992
rect 33317 17987 33383 17990
rect 5040 17984 5356 17985
rect 5040 17920 5046 17984
rect 5110 17920 5126 17984
rect 5190 17920 5206 17984
rect 5270 17920 5286 17984
rect 5350 17920 5356 17984
rect 5040 17919 5356 17920
rect 13228 17984 13544 17985
rect 13228 17920 13234 17984
rect 13298 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13544 17984
rect 13228 17919 13544 17920
rect 21416 17984 21732 17985
rect 21416 17920 21422 17984
rect 21486 17920 21502 17984
rect 21566 17920 21582 17984
rect 21646 17920 21662 17984
rect 21726 17920 21732 17984
rect 21416 17919 21732 17920
rect 29604 17984 29920 17985
rect 29604 17920 29610 17984
rect 29674 17920 29690 17984
rect 29754 17920 29770 17984
rect 29834 17920 29850 17984
rect 29914 17920 29920 17984
rect 34200 17960 35000 17990
rect 29604 17919 29920 17920
rect 9134 17440 9450 17441
rect 9134 17376 9140 17440
rect 9204 17376 9220 17440
rect 9284 17376 9300 17440
rect 9364 17376 9380 17440
rect 9444 17376 9450 17440
rect 9134 17375 9450 17376
rect 17322 17440 17638 17441
rect 17322 17376 17328 17440
rect 17392 17376 17408 17440
rect 17472 17376 17488 17440
rect 17552 17376 17568 17440
rect 17632 17376 17638 17440
rect 17322 17375 17638 17376
rect 25510 17440 25826 17441
rect 25510 17376 25516 17440
rect 25580 17376 25596 17440
rect 25660 17376 25676 17440
rect 25740 17376 25756 17440
rect 25820 17376 25826 17440
rect 25510 17375 25826 17376
rect 33698 17440 34014 17441
rect 33698 17376 33704 17440
rect 33768 17376 33784 17440
rect 33848 17376 33864 17440
rect 33928 17376 33944 17440
rect 34008 17376 34014 17440
rect 33698 17375 34014 17376
rect 5040 16896 5356 16897
rect 5040 16832 5046 16896
rect 5110 16832 5126 16896
rect 5190 16832 5206 16896
rect 5270 16832 5286 16896
rect 5350 16832 5356 16896
rect 5040 16831 5356 16832
rect 13228 16896 13544 16897
rect 13228 16832 13234 16896
rect 13298 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13544 16896
rect 13228 16831 13544 16832
rect 21416 16896 21732 16897
rect 21416 16832 21422 16896
rect 21486 16832 21502 16896
rect 21566 16832 21582 16896
rect 21646 16832 21662 16896
rect 21726 16832 21732 16896
rect 21416 16831 21732 16832
rect 29604 16896 29920 16897
rect 29604 16832 29610 16896
rect 29674 16832 29690 16896
rect 29754 16832 29770 16896
rect 29834 16832 29850 16896
rect 29914 16832 29920 16896
rect 29604 16831 29920 16832
rect 0 16690 800 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 800 16630
rect 1577 16627 1643 16630
rect 31477 16690 31543 16693
rect 34200 16690 35000 16720
rect 31477 16688 35000 16690
rect 31477 16632 31482 16688
rect 31538 16632 35000 16688
rect 31477 16630 35000 16632
rect 31477 16627 31543 16630
rect 34200 16600 35000 16630
rect 9134 16352 9450 16353
rect 9134 16288 9140 16352
rect 9204 16288 9220 16352
rect 9284 16288 9300 16352
rect 9364 16288 9380 16352
rect 9444 16288 9450 16352
rect 9134 16287 9450 16288
rect 17322 16352 17638 16353
rect 17322 16288 17328 16352
rect 17392 16288 17408 16352
rect 17472 16288 17488 16352
rect 17552 16288 17568 16352
rect 17632 16288 17638 16352
rect 17322 16287 17638 16288
rect 25510 16352 25826 16353
rect 25510 16288 25516 16352
rect 25580 16288 25596 16352
rect 25660 16288 25676 16352
rect 25740 16288 25756 16352
rect 25820 16288 25826 16352
rect 25510 16287 25826 16288
rect 33698 16352 34014 16353
rect 33698 16288 33704 16352
rect 33768 16288 33784 16352
rect 33848 16288 33864 16352
rect 33928 16288 33944 16352
rect 34008 16288 34014 16352
rect 33698 16287 34014 16288
rect 5040 15808 5356 15809
rect 5040 15744 5046 15808
rect 5110 15744 5126 15808
rect 5190 15744 5206 15808
rect 5270 15744 5286 15808
rect 5350 15744 5356 15808
rect 5040 15743 5356 15744
rect 13228 15808 13544 15809
rect 13228 15744 13234 15808
rect 13298 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13544 15808
rect 13228 15743 13544 15744
rect 21416 15808 21732 15809
rect 21416 15744 21422 15808
rect 21486 15744 21502 15808
rect 21566 15744 21582 15808
rect 21646 15744 21662 15808
rect 21726 15744 21732 15808
rect 21416 15743 21732 15744
rect 29604 15808 29920 15809
rect 29604 15744 29610 15808
rect 29674 15744 29690 15808
rect 29754 15744 29770 15808
rect 29834 15744 29850 15808
rect 29914 15744 29920 15808
rect 29604 15743 29920 15744
rect 33317 15466 33383 15469
rect 33317 15464 34162 15466
rect 33317 15408 33322 15464
rect 33378 15408 34162 15464
rect 33317 15406 34162 15408
rect 33317 15403 33383 15406
rect 34102 15364 34162 15406
rect 34102 15360 34346 15364
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 34102 15304 35000 15360
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 9134 15264 9450 15265
rect 9134 15200 9140 15264
rect 9204 15200 9220 15264
rect 9284 15200 9300 15264
rect 9364 15200 9380 15264
rect 9444 15200 9450 15264
rect 9134 15199 9450 15200
rect 17322 15264 17638 15265
rect 17322 15200 17328 15264
rect 17392 15200 17408 15264
rect 17472 15200 17488 15264
rect 17552 15200 17568 15264
rect 17632 15200 17638 15264
rect 17322 15199 17638 15200
rect 25510 15264 25826 15265
rect 25510 15200 25516 15264
rect 25580 15200 25596 15264
rect 25660 15200 25676 15264
rect 25740 15200 25756 15264
rect 25820 15200 25826 15264
rect 25510 15199 25826 15200
rect 33698 15264 34014 15265
rect 33698 15200 33704 15264
rect 33768 15200 33784 15264
rect 33848 15200 33864 15264
rect 33928 15200 33944 15264
rect 34008 15200 34014 15264
rect 34200 15240 35000 15304
rect 33698 15199 34014 15200
rect 5040 14720 5356 14721
rect 5040 14656 5046 14720
rect 5110 14656 5126 14720
rect 5190 14656 5206 14720
rect 5270 14656 5286 14720
rect 5350 14656 5356 14720
rect 5040 14655 5356 14656
rect 13228 14720 13544 14721
rect 13228 14656 13234 14720
rect 13298 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13544 14720
rect 13228 14655 13544 14656
rect 21416 14720 21732 14721
rect 21416 14656 21422 14720
rect 21486 14656 21502 14720
rect 21566 14656 21582 14720
rect 21646 14656 21662 14720
rect 21726 14656 21732 14720
rect 21416 14655 21732 14656
rect 29604 14720 29920 14721
rect 29604 14656 29610 14720
rect 29674 14656 29690 14720
rect 29754 14656 29770 14720
rect 29834 14656 29850 14720
rect 29914 14656 29920 14720
rect 29604 14655 29920 14656
rect 9134 14176 9450 14177
rect 9134 14112 9140 14176
rect 9204 14112 9220 14176
rect 9284 14112 9300 14176
rect 9364 14112 9380 14176
rect 9444 14112 9450 14176
rect 9134 14111 9450 14112
rect 17322 14176 17638 14177
rect 17322 14112 17328 14176
rect 17392 14112 17408 14176
rect 17472 14112 17488 14176
rect 17552 14112 17568 14176
rect 17632 14112 17638 14176
rect 17322 14111 17638 14112
rect 25510 14176 25826 14177
rect 25510 14112 25516 14176
rect 25580 14112 25596 14176
rect 25660 14112 25676 14176
rect 25740 14112 25756 14176
rect 25820 14112 25826 14176
rect 25510 14111 25826 14112
rect 33698 14176 34014 14177
rect 33698 14112 33704 14176
rect 33768 14112 33784 14176
rect 33848 14112 33864 14176
rect 33928 14112 33944 14176
rect 34008 14112 34014 14176
rect 33698 14111 34014 14112
rect 0 13970 800 14000
rect 1301 13970 1367 13973
rect 0 13968 1367 13970
rect 0 13912 1306 13968
rect 1362 13912 1367 13968
rect 0 13910 1367 13912
rect 0 13880 800 13910
rect 1301 13907 1367 13910
rect 31109 13970 31175 13973
rect 34200 13970 35000 14000
rect 31109 13968 35000 13970
rect 31109 13912 31114 13968
rect 31170 13912 35000 13968
rect 31109 13910 35000 13912
rect 31109 13907 31175 13910
rect 34200 13880 35000 13910
rect 5040 13632 5356 13633
rect 5040 13568 5046 13632
rect 5110 13568 5126 13632
rect 5190 13568 5206 13632
rect 5270 13568 5286 13632
rect 5350 13568 5356 13632
rect 5040 13567 5356 13568
rect 13228 13632 13544 13633
rect 13228 13568 13234 13632
rect 13298 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13544 13632
rect 13228 13567 13544 13568
rect 21416 13632 21732 13633
rect 21416 13568 21422 13632
rect 21486 13568 21502 13632
rect 21566 13568 21582 13632
rect 21646 13568 21662 13632
rect 21726 13568 21732 13632
rect 21416 13567 21732 13568
rect 29604 13632 29920 13633
rect 29604 13568 29610 13632
rect 29674 13568 29690 13632
rect 29754 13568 29770 13632
rect 29834 13568 29850 13632
rect 29914 13568 29920 13632
rect 29604 13567 29920 13568
rect 9134 13088 9450 13089
rect 9134 13024 9140 13088
rect 9204 13024 9220 13088
rect 9284 13024 9300 13088
rect 9364 13024 9380 13088
rect 9444 13024 9450 13088
rect 9134 13023 9450 13024
rect 17322 13088 17638 13089
rect 17322 13024 17328 13088
rect 17392 13024 17408 13088
rect 17472 13024 17488 13088
rect 17552 13024 17568 13088
rect 17632 13024 17638 13088
rect 17322 13023 17638 13024
rect 25510 13088 25826 13089
rect 25510 13024 25516 13088
rect 25580 13024 25596 13088
rect 25660 13024 25676 13088
rect 25740 13024 25756 13088
rect 25820 13024 25826 13088
rect 25510 13023 25826 13024
rect 33698 13088 34014 13089
rect 33698 13024 33704 13088
rect 33768 13024 33784 13088
rect 33848 13024 33864 13088
rect 33928 13024 33944 13088
rect 34008 13024 34014 13088
rect 33698 13023 34014 13024
rect 0 12610 800 12640
rect 33317 12610 33383 12613
rect 34200 12610 35000 12640
rect 0 12550 1640 12610
rect 0 12520 800 12550
rect 1580 12477 1640 12550
rect 33317 12608 35000 12610
rect 33317 12552 33322 12608
rect 33378 12552 35000 12608
rect 33317 12550 35000 12552
rect 33317 12547 33383 12550
rect 5040 12544 5356 12545
rect 5040 12480 5046 12544
rect 5110 12480 5126 12544
rect 5190 12480 5206 12544
rect 5270 12480 5286 12544
rect 5350 12480 5356 12544
rect 5040 12479 5356 12480
rect 13228 12544 13544 12545
rect 13228 12480 13234 12544
rect 13298 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13544 12544
rect 13228 12479 13544 12480
rect 21416 12544 21732 12545
rect 21416 12480 21422 12544
rect 21486 12480 21502 12544
rect 21566 12480 21582 12544
rect 21646 12480 21662 12544
rect 21726 12480 21732 12544
rect 21416 12479 21732 12480
rect 29604 12544 29920 12545
rect 29604 12480 29610 12544
rect 29674 12480 29690 12544
rect 29754 12480 29770 12544
rect 29834 12480 29850 12544
rect 29914 12480 29920 12544
rect 34200 12520 35000 12550
rect 29604 12479 29920 12480
rect 1577 12472 1643 12477
rect 1577 12416 1582 12472
rect 1638 12416 1643 12472
rect 1577 12411 1643 12416
rect 9134 12000 9450 12001
rect 9134 11936 9140 12000
rect 9204 11936 9220 12000
rect 9284 11936 9300 12000
rect 9364 11936 9380 12000
rect 9444 11936 9450 12000
rect 9134 11935 9450 11936
rect 17322 12000 17638 12001
rect 17322 11936 17328 12000
rect 17392 11936 17408 12000
rect 17472 11936 17488 12000
rect 17552 11936 17568 12000
rect 17632 11936 17638 12000
rect 17322 11935 17638 11936
rect 25510 12000 25826 12001
rect 25510 11936 25516 12000
rect 25580 11936 25596 12000
rect 25660 11936 25676 12000
rect 25740 11936 25756 12000
rect 25820 11936 25826 12000
rect 25510 11935 25826 11936
rect 33698 12000 34014 12001
rect 33698 11936 33704 12000
rect 33768 11936 33784 12000
rect 33848 11936 33864 12000
rect 33928 11936 33944 12000
rect 34008 11936 34014 12000
rect 33698 11935 34014 11936
rect 5040 11456 5356 11457
rect 5040 11392 5046 11456
rect 5110 11392 5126 11456
rect 5190 11392 5206 11456
rect 5270 11392 5286 11456
rect 5350 11392 5356 11456
rect 5040 11391 5356 11392
rect 13228 11456 13544 11457
rect 13228 11392 13234 11456
rect 13298 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13544 11456
rect 13228 11391 13544 11392
rect 21416 11456 21732 11457
rect 21416 11392 21422 11456
rect 21486 11392 21502 11456
rect 21566 11392 21582 11456
rect 21646 11392 21662 11456
rect 21726 11392 21732 11456
rect 21416 11391 21732 11392
rect 29604 11456 29920 11457
rect 29604 11392 29610 11456
rect 29674 11392 29690 11456
rect 29754 11392 29770 11456
rect 29834 11392 29850 11456
rect 29914 11392 29920 11456
rect 29604 11391 29920 11392
rect 0 11250 800 11280
rect 1301 11250 1367 11253
rect 0 11248 1367 11250
rect 0 11192 1306 11248
rect 1362 11192 1367 11248
rect 0 11190 1367 11192
rect 0 11160 800 11190
rect 1301 11187 1367 11190
rect 31477 11250 31543 11253
rect 34200 11250 35000 11280
rect 31477 11248 35000 11250
rect 31477 11192 31482 11248
rect 31538 11192 35000 11248
rect 31477 11190 35000 11192
rect 31477 11187 31543 11190
rect 34200 11160 35000 11190
rect 9134 10912 9450 10913
rect 9134 10848 9140 10912
rect 9204 10848 9220 10912
rect 9284 10848 9300 10912
rect 9364 10848 9380 10912
rect 9444 10848 9450 10912
rect 9134 10847 9450 10848
rect 17322 10912 17638 10913
rect 17322 10848 17328 10912
rect 17392 10848 17408 10912
rect 17472 10848 17488 10912
rect 17552 10848 17568 10912
rect 17632 10848 17638 10912
rect 17322 10847 17638 10848
rect 25510 10912 25826 10913
rect 25510 10848 25516 10912
rect 25580 10848 25596 10912
rect 25660 10848 25676 10912
rect 25740 10848 25756 10912
rect 25820 10848 25826 10912
rect 25510 10847 25826 10848
rect 33698 10912 34014 10913
rect 33698 10848 33704 10912
rect 33768 10848 33784 10912
rect 33848 10848 33864 10912
rect 33928 10848 33944 10912
rect 34008 10848 34014 10912
rect 33698 10847 34014 10848
rect 5040 10368 5356 10369
rect 5040 10304 5046 10368
rect 5110 10304 5126 10368
rect 5190 10304 5206 10368
rect 5270 10304 5286 10368
rect 5350 10304 5356 10368
rect 5040 10303 5356 10304
rect 13228 10368 13544 10369
rect 13228 10304 13234 10368
rect 13298 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13544 10368
rect 13228 10303 13544 10304
rect 21416 10368 21732 10369
rect 21416 10304 21422 10368
rect 21486 10304 21502 10368
rect 21566 10304 21582 10368
rect 21646 10304 21662 10368
rect 21726 10304 21732 10368
rect 21416 10303 21732 10304
rect 29604 10368 29920 10369
rect 29604 10304 29610 10368
rect 29674 10304 29690 10368
rect 29754 10304 29770 10368
rect 29834 10304 29850 10368
rect 29914 10304 29920 10368
rect 29604 10303 29920 10304
rect 0 9890 800 9920
rect 0 9830 1640 9890
rect 0 9800 800 9830
rect 1580 9757 1640 9830
rect 9134 9824 9450 9825
rect 9134 9760 9140 9824
rect 9204 9760 9220 9824
rect 9284 9760 9300 9824
rect 9364 9760 9380 9824
rect 9444 9760 9450 9824
rect 9134 9759 9450 9760
rect 17322 9824 17638 9825
rect 17322 9760 17328 9824
rect 17392 9760 17408 9824
rect 17472 9760 17488 9824
rect 17552 9760 17568 9824
rect 17632 9760 17638 9824
rect 17322 9759 17638 9760
rect 25510 9824 25826 9825
rect 25510 9760 25516 9824
rect 25580 9760 25596 9824
rect 25660 9760 25676 9824
rect 25740 9760 25756 9824
rect 25820 9760 25826 9824
rect 25510 9759 25826 9760
rect 33698 9824 34014 9825
rect 33698 9760 33704 9824
rect 33768 9760 33784 9824
rect 33848 9760 33864 9824
rect 33928 9760 33944 9824
rect 34008 9760 34014 9824
rect 34200 9800 35000 9920
rect 33698 9759 34014 9760
rect 1577 9752 1643 9757
rect 1577 9696 1582 9752
rect 1638 9696 1643 9752
rect 1577 9691 1643 9696
rect 34470 9690 34530 9800
rect 34102 9630 34530 9690
rect 33317 9618 33383 9621
rect 34102 9618 34162 9630
rect 33317 9616 34162 9618
rect 33317 9560 33322 9616
rect 33378 9560 34162 9616
rect 33317 9558 34162 9560
rect 33317 9555 33383 9558
rect 5040 9280 5356 9281
rect 5040 9216 5046 9280
rect 5110 9216 5126 9280
rect 5190 9216 5206 9280
rect 5270 9216 5286 9280
rect 5350 9216 5356 9280
rect 5040 9215 5356 9216
rect 13228 9280 13544 9281
rect 13228 9216 13234 9280
rect 13298 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13544 9280
rect 13228 9215 13544 9216
rect 21416 9280 21732 9281
rect 21416 9216 21422 9280
rect 21486 9216 21502 9280
rect 21566 9216 21582 9280
rect 21646 9216 21662 9280
rect 21726 9216 21732 9280
rect 21416 9215 21732 9216
rect 29604 9280 29920 9281
rect 29604 9216 29610 9280
rect 29674 9216 29690 9280
rect 29754 9216 29770 9280
rect 29834 9216 29850 9280
rect 29914 9216 29920 9280
rect 29604 9215 29920 9216
rect 9134 8736 9450 8737
rect 9134 8672 9140 8736
rect 9204 8672 9220 8736
rect 9284 8672 9300 8736
rect 9364 8672 9380 8736
rect 9444 8672 9450 8736
rect 9134 8671 9450 8672
rect 17322 8736 17638 8737
rect 17322 8672 17328 8736
rect 17392 8672 17408 8736
rect 17472 8672 17488 8736
rect 17552 8672 17568 8736
rect 17632 8672 17638 8736
rect 17322 8671 17638 8672
rect 25510 8736 25826 8737
rect 25510 8672 25516 8736
rect 25580 8672 25596 8736
rect 25660 8672 25676 8736
rect 25740 8672 25756 8736
rect 25820 8672 25826 8736
rect 25510 8671 25826 8672
rect 33698 8736 34014 8737
rect 33698 8672 33704 8736
rect 33768 8672 33784 8736
rect 33848 8672 33864 8736
rect 33928 8672 33944 8736
rect 34008 8672 34014 8736
rect 33698 8671 34014 8672
rect 0 8530 800 8560
rect 31293 8530 31359 8533
rect 34200 8530 35000 8560
rect 0 8470 1640 8530
rect 0 8440 800 8470
rect 1580 8397 1640 8470
rect 31293 8528 35000 8530
rect 31293 8472 31298 8528
rect 31354 8472 35000 8528
rect 31293 8470 35000 8472
rect 31293 8467 31359 8470
rect 34200 8440 35000 8470
rect 1577 8392 1643 8397
rect 1577 8336 1582 8392
rect 1638 8336 1643 8392
rect 1577 8331 1643 8336
rect 5040 8192 5356 8193
rect 5040 8128 5046 8192
rect 5110 8128 5126 8192
rect 5190 8128 5206 8192
rect 5270 8128 5286 8192
rect 5350 8128 5356 8192
rect 5040 8127 5356 8128
rect 13228 8192 13544 8193
rect 13228 8128 13234 8192
rect 13298 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13544 8192
rect 13228 8127 13544 8128
rect 21416 8192 21732 8193
rect 21416 8128 21422 8192
rect 21486 8128 21502 8192
rect 21566 8128 21582 8192
rect 21646 8128 21662 8192
rect 21726 8128 21732 8192
rect 21416 8127 21732 8128
rect 29604 8192 29920 8193
rect 29604 8128 29610 8192
rect 29674 8128 29690 8192
rect 29754 8128 29770 8192
rect 29834 8128 29850 8192
rect 29914 8128 29920 8192
rect 29604 8127 29920 8128
rect 9134 7648 9450 7649
rect 9134 7584 9140 7648
rect 9204 7584 9220 7648
rect 9284 7584 9300 7648
rect 9364 7584 9380 7648
rect 9444 7584 9450 7648
rect 9134 7583 9450 7584
rect 17322 7648 17638 7649
rect 17322 7584 17328 7648
rect 17392 7584 17408 7648
rect 17472 7584 17488 7648
rect 17552 7584 17568 7648
rect 17632 7584 17638 7648
rect 17322 7583 17638 7584
rect 25510 7648 25826 7649
rect 25510 7584 25516 7648
rect 25580 7584 25596 7648
rect 25660 7584 25676 7648
rect 25740 7584 25756 7648
rect 25820 7584 25826 7648
rect 25510 7583 25826 7584
rect 33698 7648 34014 7649
rect 33698 7584 33704 7648
rect 33768 7584 33784 7648
rect 33848 7584 33864 7648
rect 33928 7584 33944 7648
rect 34008 7584 34014 7648
rect 33698 7583 34014 7584
rect 0 7170 800 7200
rect 33317 7170 33383 7173
rect 34200 7170 35000 7200
rect 0 7110 1640 7170
rect 0 7080 800 7110
rect 1580 7037 1640 7110
rect 33317 7168 35000 7170
rect 33317 7112 33322 7168
rect 33378 7112 35000 7168
rect 33317 7110 35000 7112
rect 33317 7107 33383 7110
rect 5040 7104 5356 7105
rect 5040 7040 5046 7104
rect 5110 7040 5126 7104
rect 5190 7040 5206 7104
rect 5270 7040 5286 7104
rect 5350 7040 5356 7104
rect 5040 7039 5356 7040
rect 13228 7104 13544 7105
rect 13228 7040 13234 7104
rect 13298 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13544 7104
rect 13228 7039 13544 7040
rect 21416 7104 21732 7105
rect 21416 7040 21422 7104
rect 21486 7040 21502 7104
rect 21566 7040 21582 7104
rect 21646 7040 21662 7104
rect 21726 7040 21732 7104
rect 21416 7039 21732 7040
rect 29604 7104 29920 7105
rect 29604 7040 29610 7104
rect 29674 7040 29690 7104
rect 29754 7040 29770 7104
rect 29834 7040 29850 7104
rect 29914 7040 29920 7104
rect 34200 7080 35000 7110
rect 29604 7039 29920 7040
rect 1577 7032 1643 7037
rect 1577 6976 1582 7032
rect 1638 6976 1643 7032
rect 1577 6971 1643 6976
rect 9134 6560 9450 6561
rect 9134 6496 9140 6560
rect 9204 6496 9220 6560
rect 9284 6496 9300 6560
rect 9364 6496 9380 6560
rect 9444 6496 9450 6560
rect 9134 6495 9450 6496
rect 17322 6560 17638 6561
rect 17322 6496 17328 6560
rect 17392 6496 17408 6560
rect 17472 6496 17488 6560
rect 17552 6496 17568 6560
rect 17632 6496 17638 6560
rect 17322 6495 17638 6496
rect 25510 6560 25826 6561
rect 25510 6496 25516 6560
rect 25580 6496 25596 6560
rect 25660 6496 25676 6560
rect 25740 6496 25756 6560
rect 25820 6496 25826 6560
rect 25510 6495 25826 6496
rect 33698 6560 34014 6561
rect 33698 6496 33704 6560
rect 33768 6496 33784 6560
rect 33848 6496 33864 6560
rect 33928 6496 33944 6560
rect 34008 6496 34014 6560
rect 33698 6495 34014 6496
rect 5040 6016 5356 6017
rect 5040 5952 5046 6016
rect 5110 5952 5126 6016
rect 5190 5952 5206 6016
rect 5270 5952 5286 6016
rect 5350 5952 5356 6016
rect 5040 5951 5356 5952
rect 13228 6016 13544 6017
rect 13228 5952 13234 6016
rect 13298 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13544 6016
rect 13228 5951 13544 5952
rect 21416 6016 21732 6017
rect 21416 5952 21422 6016
rect 21486 5952 21502 6016
rect 21566 5952 21582 6016
rect 21646 5952 21662 6016
rect 21726 5952 21732 6016
rect 21416 5951 21732 5952
rect 29604 6016 29920 6017
rect 29604 5952 29610 6016
rect 29674 5952 29690 6016
rect 29754 5952 29770 6016
rect 29834 5952 29850 6016
rect 29914 5952 29920 6016
rect 29604 5951 29920 5952
rect 0 5810 800 5840
rect 1301 5810 1367 5813
rect 0 5808 1367 5810
rect 0 5752 1306 5808
rect 1362 5752 1367 5808
rect 0 5750 1367 5752
rect 0 5720 800 5750
rect 1301 5747 1367 5750
rect 26417 5810 26483 5813
rect 27521 5810 27587 5813
rect 30741 5810 30807 5813
rect 26417 5808 30807 5810
rect 26417 5752 26422 5808
rect 26478 5752 27526 5808
rect 27582 5752 30746 5808
rect 30802 5752 30807 5808
rect 26417 5750 30807 5752
rect 26417 5747 26483 5750
rect 27521 5747 27587 5750
rect 30741 5747 30807 5750
rect 31477 5810 31543 5813
rect 34200 5810 35000 5840
rect 31477 5808 35000 5810
rect 31477 5752 31482 5808
rect 31538 5752 35000 5808
rect 31477 5750 35000 5752
rect 31477 5747 31543 5750
rect 34200 5720 35000 5750
rect 26693 5674 26759 5677
rect 33501 5674 33567 5677
rect 26693 5672 33567 5674
rect 26693 5616 26698 5672
rect 26754 5616 33506 5672
rect 33562 5616 33567 5672
rect 26693 5614 33567 5616
rect 26693 5611 26759 5614
rect 33501 5611 33567 5614
rect 9134 5472 9450 5473
rect 9134 5408 9140 5472
rect 9204 5408 9220 5472
rect 9284 5408 9300 5472
rect 9364 5408 9380 5472
rect 9444 5408 9450 5472
rect 9134 5407 9450 5408
rect 17322 5472 17638 5473
rect 17322 5408 17328 5472
rect 17392 5408 17408 5472
rect 17472 5408 17488 5472
rect 17552 5408 17568 5472
rect 17632 5408 17638 5472
rect 17322 5407 17638 5408
rect 25510 5472 25826 5473
rect 25510 5408 25516 5472
rect 25580 5408 25596 5472
rect 25660 5408 25676 5472
rect 25740 5408 25756 5472
rect 25820 5408 25826 5472
rect 25510 5407 25826 5408
rect 33698 5472 34014 5473
rect 33698 5408 33704 5472
rect 33768 5408 33784 5472
rect 33848 5408 33864 5472
rect 33928 5408 33944 5472
rect 34008 5408 34014 5472
rect 33698 5407 34014 5408
rect 26049 5266 26115 5269
rect 29177 5266 29243 5269
rect 26049 5264 29243 5266
rect 26049 5208 26054 5264
rect 26110 5208 29182 5264
rect 29238 5208 29243 5264
rect 26049 5206 29243 5208
rect 26049 5203 26115 5206
rect 29177 5203 29243 5206
rect 5040 4928 5356 4929
rect 5040 4864 5046 4928
rect 5110 4864 5126 4928
rect 5190 4864 5206 4928
rect 5270 4864 5286 4928
rect 5350 4864 5356 4928
rect 5040 4863 5356 4864
rect 13228 4928 13544 4929
rect 13228 4864 13234 4928
rect 13298 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13544 4928
rect 13228 4863 13544 4864
rect 21416 4928 21732 4929
rect 21416 4864 21422 4928
rect 21486 4864 21502 4928
rect 21566 4864 21582 4928
rect 21646 4864 21662 4928
rect 21726 4864 21732 4928
rect 21416 4863 21732 4864
rect 29604 4928 29920 4929
rect 29604 4864 29610 4928
rect 29674 4864 29690 4928
rect 29754 4864 29770 4928
rect 29834 4864 29850 4928
rect 29914 4864 29920 4928
rect 29604 4863 29920 4864
rect 23933 4722 23999 4725
rect 32213 4722 32279 4725
rect 23933 4720 32279 4722
rect 23933 4664 23938 4720
rect 23994 4664 32218 4720
rect 32274 4664 32279 4720
rect 23933 4662 32279 4664
rect 23933 4659 23999 4662
rect 32213 4659 32279 4662
rect 31569 4586 31635 4589
rect 31569 4584 34162 4586
rect 31569 4528 31574 4584
rect 31630 4528 34162 4584
rect 31569 4526 34162 4528
rect 31569 4523 31635 4526
rect 34102 4484 34162 4526
rect 34102 4480 34346 4484
rect 0 4450 800 4480
rect 0 4390 1640 4450
rect 34102 4424 35000 4480
rect 0 4360 800 4390
rect 1580 4181 1640 4390
rect 9134 4384 9450 4385
rect 9134 4320 9140 4384
rect 9204 4320 9220 4384
rect 9284 4320 9300 4384
rect 9364 4320 9380 4384
rect 9444 4320 9450 4384
rect 9134 4319 9450 4320
rect 17322 4384 17638 4385
rect 17322 4320 17328 4384
rect 17392 4320 17408 4384
rect 17472 4320 17488 4384
rect 17552 4320 17568 4384
rect 17632 4320 17638 4384
rect 17322 4319 17638 4320
rect 25510 4384 25826 4385
rect 25510 4320 25516 4384
rect 25580 4320 25596 4384
rect 25660 4320 25676 4384
rect 25740 4320 25756 4384
rect 25820 4320 25826 4384
rect 25510 4319 25826 4320
rect 33698 4384 34014 4385
rect 33698 4320 33704 4384
rect 33768 4320 33784 4384
rect 33848 4320 33864 4384
rect 33928 4320 33944 4384
rect 34008 4320 34014 4384
rect 34200 4360 35000 4424
rect 33698 4319 34014 4320
rect 1577 4176 1643 4181
rect 1577 4120 1582 4176
rect 1638 4120 1643 4176
rect 1577 4115 1643 4120
rect 5040 3840 5356 3841
rect 5040 3776 5046 3840
rect 5110 3776 5126 3840
rect 5190 3776 5206 3840
rect 5270 3776 5286 3840
rect 5350 3776 5356 3840
rect 5040 3775 5356 3776
rect 13228 3840 13544 3841
rect 13228 3776 13234 3840
rect 13298 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13544 3840
rect 13228 3775 13544 3776
rect 21416 3840 21732 3841
rect 21416 3776 21422 3840
rect 21486 3776 21502 3840
rect 21566 3776 21582 3840
rect 21646 3776 21662 3840
rect 21726 3776 21732 3840
rect 21416 3775 21732 3776
rect 29604 3840 29920 3841
rect 29604 3776 29610 3840
rect 29674 3776 29690 3840
rect 29754 3776 29770 3840
rect 29834 3776 29850 3840
rect 29914 3776 29920 3840
rect 29604 3775 29920 3776
rect 9134 3296 9450 3297
rect 9134 3232 9140 3296
rect 9204 3232 9220 3296
rect 9284 3232 9300 3296
rect 9364 3232 9380 3296
rect 9444 3232 9450 3296
rect 9134 3231 9450 3232
rect 17322 3296 17638 3297
rect 17322 3232 17328 3296
rect 17392 3232 17408 3296
rect 17472 3232 17488 3296
rect 17552 3232 17568 3296
rect 17632 3232 17638 3296
rect 17322 3231 17638 3232
rect 25510 3296 25826 3297
rect 25510 3232 25516 3296
rect 25580 3232 25596 3296
rect 25660 3232 25676 3296
rect 25740 3232 25756 3296
rect 25820 3232 25826 3296
rect 25510 3231 25826 3232
rect 33698 3296 34014 3297
rect 33698 3232 33704 3296
rect 33768 3232 33784 3296
rect 33848 3232 33864 3296
rect 33928 3232 33944 3296
rect 34008 3232 34014 3296
rect 33698 3231 34014 3232
rect 0 3090 800 3120
rect 33501 3090 33567 3093
rect 34200 3090 35000 3120
rect 0 3030 1640 3090
rect 0 3000 800 3030
rect 1580 2821 1640 3030
rect 33501 3088 35000 3090
rect 33501 3032 33506 3088
rect 33562 3032 35000 3088
rect 33501 3030 35000 3032
rect 33501 3027 33567 3030
rect 34200 3000 35000 3030
rect 1577 2816 1643 2821
rect 1577 2760 1582 2816
rect 1638 2760 1643 2816
rect 1577 2755 1643 2760
rect 5040 2752 5356 2753
rect 5040 2688 5046 2752
rect 5110 2688 5126 2752
rect 5190 2688 5206 2752
rect 5270 2688 5286 2752
rect 5350 2688 5356 2752
rect 5040 2687 5356 2688
rect 13228 2752 13544 2753
rect 13228 2688 13234 2752
rect 13298 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13544 2752
rect 13228 2687 13544 2688
rect 21416 2752 21732 2753
rect 21416 2688 21422 2752
rect 21486 2688 21502 2752
rect 21566 2688 21582 2752
rect 21646 2688 21662 2752
rect 21726 2688 21732 2752
rect 21416 2687 21732 2688
rect 29604 2752 29920 2753
rect 29604 2688 29610 2752
rect 29674 2688 29690 2752
rect 29754 2688 29770 2752
rect 29834 2688 29850 2752
rect 29914 2688 29920 2752
rect 29604 2687 29920 2688
rect 9134 2208 9450 2209
rect 9134 2144 9140 2208
rect 9204 2144 9220 2208
rect 9284 2144 9300 2208
rect 9364 2144 9380 2208
rect 9444 2144 9450 2208
rect 9134 2143 9450 2144
rect 17322 2208 17638 2209
rect 17322 2144 17328 2208
rect 17392 2144 17408 2208
rect 17472 2144 17488 2208
rect 17552 2144 17568 2208
rect 17632 2144 17638 2208
rect 17322 2143 17638 2144
rect 25510 2208 25826 2209
rect 25510 2144 25516 2208
rect 25580 2144 25596 2208
rect 25660 2144 25676 2208
rect 25740 2144 25756 2208
rect 25820 2144 25826 2208
rect 25510 2143 25826 2144
rect 33698 2208 34014 2209
rect 33698 2144 33704 2208
rect 33768 2144 33784 2208
rect 33848 2144 33864 2208
rect 33928 2144 33944 2208
rect 34008 2144 34014 2208
rect 33698 2143 34014 2144
rect 29545 1730 29611 1733
rect 34200 1730 35000 1760
rect 29545 1728 35000 1730
rect 29545 1672 29550 1728
rect 29606 1672 35000 1728
rect 29545 1670 35000 1672
rect 29545 1667 29611 1670
rect 34200 1640 35000 1670
<< via3 >>
rect 9140 32668 9204 32672
rect 9140 32612 9144 32668
rect 9144 32612 9200 32668
rect 9200 32612 9204 32668
rect 9140 32608 9204 32612
rect 9220 32668 9284 32672
rect 9220 32612 9224 32668
rect 9224 32612 9280 32668
rect 9280 32612 9284 32668
rect 9220 32608 9284 32612
rect 9300 32668 9364 32672
rect 9300 32612 9304 32668
rect 9304 32612 9360 32668
rect 9360 32612 9364 32668
rect 9300 32608 9364 32612
rect 9380 32668 9444 32672
rect 9380 32612 9384 32668
rect 9384 32612 9440 32668
rect 9440 32612 9444 32668
rect 9380 32608 9444 32612
rect 17328 32668 17392 32672
rect 17328 32612 17332 32668
rect 17332 32612 17388 32668
rect 17388 32612 17392 32668
rect 17328 32608 17392 32612
rect 17408 32668 17472 32672
rect 17408 32612 17412 32668
rect 17412 32612 17468 32668
rect 17468 32612 17472 32668
rect 17408 32608 17472 32612
rect 17488 32668 17552 32672
rect 17488 32612 17492 32668
rect 17492 32612 17548 32668
rect 17548 32612 17552 32668
rect 17488 32608 17552 32612
rect 17568 32668 17632 32672
rect 17568 32612 17572 32668
rect 17572 32612 17628 32668
rect 17628 32612 17632 32668
rect 17568 32608 17632 32612
rect 25516 32668 25580 32672
rect 25516 32612 25520 32668
rect 25520 32612 25576 32668
rect 25576 32612 25580 32668
rect 25516 32608 25580 32612
rect 25596 32668 25660 32672
rect 25596 32612 25600 32668
rect 25600 32612 25656 32668
rect 25656 32612 25660 32668
rect 25596 32608 25660 32612
rect 25676 32668 25740 32672
rect 25676 32612 25680 32668
rect 25680 32612 25736 32668
rect 25736 32612 25740 32668
rect 25676 32608 25740 32612
rect 25756 32668 25820 32672
rect 25756 32612 25760 32668
rect 25760 32612 25816 32668
rect 25816 32612 25820 32668
rect 25756 32608 25820 32612
rect 33704 32668 33768 32672
rect 33704 32612 33708 32668
rect 33708 32612 33764 32668
rect 33764 32612 33768 32668
rect 33704 32608 33768 32612
rect 33784 32668 33848 32672
rect 33784 32612 33788 32668
rect 33788 32612 33844 32668
rect 33844 32612 33848 32668
rect 33784 32608 33848 32612
rect 33864 32668 33928 32672
rect 33864 32612 33868 32668
rect 33868 32612 33924 32668
rect 33924 32612 33928 32668
rect 33864 32608 33928 32612
rect 33944 32668 34008 32672
rect 33944 32612 33948 32668
rect 33948 32612 34004 32668
rect 34004 32612 34008 32668
rect 33944 32608 34008 32612
rect 5046 32124 5110 32128
rect 5046 32068 5050 32124
rect 5050 32068 5106 32124
rect 5106 32068 5110 32124
rect 5046 32064 5110 32068
rect 5126 32124 5190 32128
rect 5126 32068 5130 32124
rect 5130 32068 5186 32124
rect 5186 32068 5190 32124
rect 5126 32064 5190 32068
rect 5206 32124 5270 32128
rect 5206 32068 5210 32124
rect 5210 32068 5266 32124
rect 5266 32068 5270 32124
rect 5206 32064 5270 32068
rect 5286 32124 5350 32128
rect 5286 32068 5290 32124
rect 5290 32068 5346 32124
rect 5346 32068 5350 32124
rect 5286 32064 5350 32068
rect 13234 32124 13298 32128
rect 13234 32068 13238 32124
rect 13238 32068 13294 32124
rect 13294 32068 13298 32124
rect 13234 32064 13298 32068
rect 13314 32124 13378 32128
rect 13314 32068 13318 32124
rect 13318 32068 13374 32124
rect 13374 32068 13378 32124
rect 13314 32064 13378 32068
rect 13394 32124 13458 32128
rect 13394 32068 13398 32124
rect 13398 32068 13454 32124
rect 13454 32068 13458 32124
rect 13394 32064 13458 32068
rect 13474 32124 13538 32128
rect 13474 32068 13478 32124
rect 13478 32068 13534 32124
rect 13534 32068 13538 32124
rect 13474 32064 13538 32068
rect 21422 32124 21486 32128
rect 21422 32068 21426 32124
rect 21426 32068 21482 32124
rect 21482 32068 21486 32124
rect 21422 32064 21486 32068
rect 21502 32124 21566 32128
rect 21502 32068 21506 32124
rect 21506 32068 21562 32124
rect 21562 32068 21566 32124
rect 21502 32064 21566 32068
rect 21582 32124 21646 32128
rect 21582 32068 21586 32124
rect 21586 32068 21642 32124
rect 21642 32068 21646 32124
rect 21582 32064 21646 32068
rect 21662 32124 21726 32128
rect 21662 32068 21666 32124
rect 21666 32068 21722 32124
rect 21722 32068 21726 32124
rect 21662 32064 21726 32068
rect 29610 32124 29674 32128
rect 29610 32068 29614 32124
rect 29614 32068 29670 32124
rect 29670 32068 29674 32124
rect 29610 32064 29674 32068
rect 29690 32124 29754 32128
rect 29690 32068 29694 32124
rect 29694 32068 29750 32124
rect 29750 32068 29754 32124
rect 29690 32064 29754 32068
rect 29770 32124 29834 32128
rect 29770 32068 29774 32124
rect 29774 32068 29830 32124
rect 29830 32068 29834 32124
rect 29770 32064 29834 32068
rect 29850 32124 29914 32128
rect 29850 32068 29854 32124
rect 29854 32068 29910 32124
rect 29910 32068 29914 32124
rect 29850 32064 29914 32068
rect 9140 31580 9204 31584
rect 9140 31524 9144 31580
rect 9144 31524 9200 31580
rect 9200 31524 9204 31580
rect 9140 31520 9204 31524
rect 9220 31580 9284 31584
rect 9220 31524 9224 31580
rect 9224 31524 9280 31580
rect 9280 31524 9284 31580
rect 9220 31520 9284 31524
rect 9300 31580 9364 31584
rect 9300 31524 9304 31580
rect 9304 31524 9360 31580
rect 9360 31524 9364 31580
rect 9300 31520 9364 31524
rect 9380 31580 9444 31584
rect 9380 31524 9384 31580
rect 9384 31524 9440 31580
rect 9440 31524 9444 31580
rect 9380 31520 9444 31524
rect 17328 31580 17392 31584
rect 17328 31524 17332 31580
rect 17332 31524 17388 31580
rect 17388 31524 17392 31580
rect 17328 31520 17392 31524
rect 17408 31580 17472 31584
rect 17408 31524 17412 31580
rect 17412 31524 17468 31580
rect 17468 31524 17472 31580
rect 17408 31520 17472 31524
rect 17488 31580 17552 31584
rect 17488 31524 17492 31580
rect 17492 31524 17548 31580
rect 17548 31524 17552 31580
rect 17488 31520 17552 31524
rect 17568 31580 17632 31584
rect 17568 31524 17572 31580
rect 17572 31524 17628 31580
rect 17628 31524 17632 31580
rect 17568 31520 17632 31524
rect 25516 31580 25580 31584
rect 25516 31524 25520 31580
rect 25520 31524 25576 31580
rect 25576 31524 25580 31580
rect 25516 31520 25580 31524
rect 25596 31580 25660 31584
rect 25596 31524 25600 31580
rect 25600 31524 25656 31580
rect 25656 31524 25660 31580
rect 25596 31520 25660 31524
rect 25676 31580 25740 31584
rect 25676 31524 25680 31580
rect 25680 31524 25736 31580
rect 25736 31524 25740 31580
rect 25676 31520 25740 31524
rect 25756 31580 25820 31584
rect 25756 31524 25760 31580
rect 25760 31524 25816 31580
rect 25816 31524 25820 31580
rect 25756 31520 25820 31524
rect 33704 31580 33768 31584
rect 33704 31524 33708 31580
rect 33708 31524 33764 31580
rect 33764 31524 33768 31580
rect 33704 31520 33768 31524
rect 33784 31580 33848 31584
rect 33784 31524 33788 31580
rect 33788 31524 33844 31580
rect 33844 31524 33848 31580
rect 33784 31520 33848 31524
rect 33864 31580 33928 31584
rect 33864 31524 33868 31580
rect 33868 31524 33924 31580
rect 33924 31524 33928 31580
rect 33864 31520 33928 31524
rect 33944 31580 34008 31584
rect 33944 31524 33948 31580
rect 33948 31524 34004 31580
rect 34004 31524 34008 31580
rect 33944 31520 34008 31524
rect 5046 31036 5110 31040
rect 5046 30980 5050 31036
rect 5050 30980 5106 31036
rect 5106 30980 5110 31036
rect 5046 30976 5110 30980
rect 5126 31036 5190 31040
rect 5126 30980 5130 31036
rect 5130 30980 5186 31036
rect 5186 30980 5190 31036
rect 5126 30976 5190 30980
rect 5206 31036 5270 31040
rect 5206 30980 5210 31036
rect 5210 30980 5266 31036
rect 5266 30980 5270 31036
rect 5206 30976 5270 30980
rect 5286 31036 5350 31040
rect 5286 30980 5290 31036
rect 5290 30980 5346 31036
rect 5346 30980 5350 31036
rect 5286 30976 5350 30980
rect 13234 31036 13298 31040
rect 13234 30980 13238 31036
rect 13238 30980 13294 31036
rect 13294 30980 13298 31036
rect 13234 30976 13298 30980
rect 13314 31036 13378 31040
rect 13314 30980 13318 31036
rect 13318 30980 13374 31036
rect 13374 30980 13378 31036
rect 13314 30976 13378 30980
rect 13394 31036 13458 31040
rect 13394 30980 13398 31036
rect 13398 30980 13454 31036
rect 13454 30980 13458 31036
rect 13394 30976 13458 30980
rect 13474 31036 13538 31040
rect 13474 30980 13478 31036
rect 13478 30980 13534 31036
rect 13534 30980 13538 31036
rect 13474 30976 13538 30980
rect 21422 31036 21486 31040
rect 21422 30980 21426 31036
rect 21426 30980 21482 31036
rect 21482 30980 21486 31036
rect 21422 30976 21486 30980
rect 21502 31036 21566 31040
rect 21502 30980 21506 31036
rect 21506 30980 21562 31036
rect 21562 30980 21566 31036
rect 21502 30976 21566 30980
rect 21582 31036 21646 31040
rect 21582 30980 21586 31036
rect 21586 30980 21642 31036
rect 21642 30980 21646 31036
rect 21582 30976 21646 30980
rect 21662 31036 21726 31040
rect 21662 30980 21666 31036
rect 21666 30980 21722 31036
rect 21722 30980 21726 31036
rect 21662 30976 21726 30980
rect 29610 31036 29674 31040
rect 29610 30980 29614 31036
rect 29614 30980 29670 31036
rect 29670 30980 29674 31036
rect 29610 30976 29674 30980
rect 29690 31036 29754 31040
rect 29690 30980 29694 31036
rect 29694 30980 29750 31036
rect 29750 30980 29754 31036
rect 29690 30976 29754 30980
rect 29770 31036 29834 31040
rect 29770 30980 29774 31036
rect 29774 30980 29830 31036
rect 29830 30980 29834 31036
rect 29770 30976 29834 30980
rect 29850 31036 29914 31040
rect 29850 30980 29854 31036
rect 29854 30980 29910 31036
rect 29910 30980 29914 31036
rect 29850 30976 29914 30980
rect 9140 30492 9204 30496
rect 9140 30436 9144 30492
rect 9144 30436 9200 30492
rect 9200 30436 9204 30492
rect 9140 30432 9204 30436
rect 9220 30492 9284 30496
rect 9220 30436 9224 30492
rect 9224 30436 9280 30492
rect 9280 30436 9284 30492
rect 9220 30432 9284 30436
rect 9300 30492 9364 30496
rect 9300 30436 9304 30492
rect 9304 30436 9360 30492
rect 9360 30436 9364 30492
rect 9300 30432 9364 30436
rect 9380 30492 9444 30496
rect 9380 30436 9384 30492
rect 9384 30436 9440 30492
rect 9440 30436 9444 30492
rect 9380 30432 9444 30436
rect 17328 30492 17392 30496
rect 17328 30436 17332 30492
rect 17332 30436 17388 30492
rect 17388 30436 17392 30492
rect 17328 30432 17392 30436
rect 17408 30492 17472 30496
rect 17408 30436 17412 30492
rect 17412 30436 17468 30492
rect 17468 30436 17472 30492
rect 17408 30432 17472 30436
rect 17488 30492 17552 30496
rect 17488 30436 17492 30492
rect 17492 30436 17548 30492
rect 17548 30436 17552 30492
rect 17488 30432 17552 30436
rect 17568 30492 17632 30496
rect 17568 30436 17572 30492
rect 17572 30436 17628 30492
rect 17628 30436 17632 30492
rect 17568 30432 17632 30436
rect 25516 30492 25580 30496
rect 25516 30436 25520 30492
rect 25520 30436 25576 30492
rect 25576 30436 25580 30492
rect 25516 30432 25580 30436
rect 25596 30492 25660 30496
rect 25596 30436 25600 30492
rect 25600 30436 25656 30492
rect 25656 30436 25660 30492
rect 25596 30432 25660 30436
rect 25676 30492 25740 30496
rect 25676 30436 25680 30492
rect 25680 30436 25736 30492
rect 25736 30436 25740 30492
rect 25676 30432 25740 30436
rect 25756 30492 25820 30496
rect 25756 30436 25760 30492
rect 25760 30436 25816 30492
rect 25816 30436 25820 30492
rect 25756 30432 25820 30436
rect 33704 30492 33768 30496
rect 33704 30436 33708 30492
rect 33708 30436 33764 30492
rect 33764 30436 33768 30492
rect 33704 30432 33768 30436
rect 33784 30492 33848 30496
rect 33784 30436 33788 30492
rect 33788 30436 33844 30492
rect 33844 30436 33848 30492
rect 33784 30432 33848 30436
rect 33864 30492 33928 30496
rect 33864 30436 33868 30492
rect 33868 30436 33924 30492
rect 33924 30436 33928 30492
rect 33864 30432 33928 30436
rect 33944 30492 34008 30496
rect 33944 30436 33948 30492
rect 33948 30436 34004 30492
rect 34004 30436 34008 30492
rect 33944 30432 34008 30436
rect 5046 29948 5110 29952
rect 5046 29892 5050 29948
rect 5050 29892 5106 29948
rect 5106 29892 5110 29948
rect 5046 29888 5110 29892
rect 5126 29948 5190 29952
rect 5126 29892 5130 29948
rect 5130 29892 5186 29948
rect 5186 29892 5190 29948
rect 5126 29888 5190 29892
rect 5206 29948 5270 29952
rect 5206 29892 5210 29948
rect 5210 29892 5266 29948
rect 5266 29892 5270 29948
rect 5206 29888 5270 29892
rect 5286 29948 5350 29952
rect 5286 29892 5290 29948
rect 5290 29892 5346 29948
rect 5346 29892 5350 29948
rect 5286 29888 5350 29892
rect 13234 29948 13298 29952
rect 13234 29892 13238 29948
rect 13238 29892 13294 29948
rect 13294 29892 13298 29948
rect 13234 29888 13298 29892
rect 13314 29948 13378 29952
rect 13314 29892 13318 29948
rect 13318 29892 13374 29948
rect 13374 29892 13378 29948
rect 13314 29888 13378 29892
rect 13394 29948 13458 29952
rect 13394 29892 13398 29948
rect 13398 29892 13454 29948
rect 13454 29892 13458 29948
rect 13394 29888 13458 29892
rect 13474 29948 13538 29952
rect 13474 29892 13478 29948
rect 13478 29892 13534 29948
rect 13534 29892 13538 29948
rect 13474 29888 13538 29892
rect 21422 29948 21486 29952
rect 21422 29892 21426 29948
rect 21426 29892 21482 29948
rect 21482 29892 21486 29948
rect 21422 29888 21486 29892
rect 21502 29948 21566 29952
rect 21502 29892 21506 29948
rect 21506 29892 21562 29948
rect 21562 29892 21566 29948
rect 21502 29888 21566 29892
rect 21582 29948 21646 29952
rect 21582 29892 21586 29948
rect 21586 29892 21642 29948
rect 21642 29892 21646 29948
rect 21582 29888 21646 29892
rect 21662 29948 21726 29952
rect 21662 29892 21666 29948
rect 21666 29892 21722 29948
rect 21722 29892 21726 29948
rect 21662 29888 21726 29892
rect 29610 29948 29674 29952
rect 29610 29892 29614 29948
rect 29614 29892 29670 29948
rect 29670 29892 29674 29948
rect 29610 29888 29674 29892
rect 29690 29948 29754 29952
rect 29690 29892 29694 29948
rect 29694 29892 29750 29948
rect 29750 29892 29754 29948
rect 29690 29888 29754 29892
rect 29770 29948 29834 29952
rect 29770 29892 29774 29948
rect 29774 29892 29830 29948
rect 29830 29892 29834 29948
rect 29770 29888 29834 29892
rect 29850 29948 29914 29952
rect 29850 29892 29854 29948
rect 29854 29892 29910 29948
rect 29910 29892 29914 29948
rect 29850 29888 29914 29892
rect 9140 29404 9204 29408
rect 9140 29348 9144 29404
rect 9144 29348 9200 29404
rect 9200 29348 9204 29404
rect 9140 29344 9204 29348
rect 9220 29404 9284 29408
rect 9220 29348 9224 29404
rect 9224 29348 9280 29404
rect 9280 29348 9284 29404
rect 9220 29344 9284 29348
rect 9300 29404 9364 29408
rect 9300 29348 9304 29404
rect 9304 29348 9360 29404
rect 9360 29348 9364 29404
rect 9300 29344 9364 29348
rect 9380 29404 9444 29408
rect 9380 29348 9384 29404
rect 9384 29348 9440 29404
rect 9440 29348 9444 29404
rect 9380 29344 9444 29348
rect 17328 29404 17392 29408
rect 17328 29348 17332 29404
rect 17332 29348 17388 29404
rect 17388 29348 17392 29404
rect 17328 29344 17392 29348
rect 17408 29404 17472 29408
rect 17408 29348 17412 29404
rect 17412 29348 17468 29404
rect 17468 29348 17472 29404
rect 17408 29344 17472 29348
rect 17488 29404 17552 29408
rect 17488 29348 17492 29404
rect 17492 29348 17548 29404
rect 17548 29348 17552 29404
rect 17488 29344 17552 29348
rect 17568 29404 17632 29408
rect 17568 29348 17572 29404
rect 17572 29348 17628 29404
rect 17628 29348 17632 29404
rect 17568 29344 17632 29348
rect 25516 29404 25580 29408
rect 25516 29348 25520 29404
rect 25520 29348 25576 29404
rect 25576 29348 25580 29404
rect 25516 29344 25580 29348
rect 25596 29404 25660 29408
rect 25596 29348 25600 29404
rect 25600 29348 25656 29404
rect 25656 29348 25660 29404
rect 25596 29344 25660 29348
rect 25676 29404 25740 29408
rect 25676 29348 25680 29404
rect 25680 29348 25736 29404
rect 25736 29348 25740 29404
rect 25676 29344 25740 29348
rect 25756 29404 25820 29408
rect 25756 29348 25760 29404
rect 25760 29348 25816 29404
rect 25816 29348 25820 29404
rect 25756 29344 25820 29348
rect 33704 29404 33768 29408
rect 33704 29348 33708 29404
rect 33708 29348 33764 29404
rect 33764 29348 33768 29404
rect 33704 29344 33768 29348
rect 33784 29404 33848 29408
rect 33784 29348 33788 29404
rect 33788 29348 33844 29404
rect 33844 29348 33848 29404
rect 33784 29344 33848 29348
rect 33864 29404 33928 29408
rect 33864 29348 33868 29404
rect 33868 29348 33924 29404
rect 33924 29348 33928 29404
rect 33864 29344 33928 29348
rect 33944 29404 34008 29408
rect 33944 29348 33948 29404
rect 33948 29348 34004 29404
rect 34004 29348 34008 29404
rect 33944 29344 34008 29348
rect 5046 28860 5110 28864
rect 5046 28804 5050 28860
rect 5050 28804 5106 28860
rect 5106 28804 5110 28860
rect 5046 28800 5110 28804
rect 5126 28860 5190 28864
rect 5126 28804 5130 28860
rect 5130 28804 5186 28860
rect 5186 28804 5190 28860
rect 5126 28800 5190 28804
rect 5206 28860 5270 28864
rect 5206 28804 5210 28860
rect 5210 28804 5266 28860
rect 5266 28804 5270 28860
rect 5206 28800 5270 28804
rect 5286 28860 5350 28864
rect 5286 28804 5290 28860
rect 5290 28804 5346 28860
rect 5346 28804 5350 28860
rect 5286 28800 5350 28804
rect 13234 28860 13298 28864
rect 13234 28804 13238 28860
rect 13238 28804 13294 28860
rect 13294 28804 13298 28860
rect 13234 28800 13298 28804
rect 13314 28860 13378 28864
rect 13314 28804 13318 28860
rect 13318 28804 13374 28860
rect 13374 28804 13378 28860
rect 13314 28800 13378 28804
rect 13394 28860 13458 28864
rect 13394 28804 13398 28860
rect 13398 28804 13454 28860
rect 13454 28804 13458 28860
rect 13394 28800 13458 28804
rect 13474 28860 13538 28864
rect 13474 28804 13478 28860
rect 13478 28804 13534 28860
rect 13534 28804 13538 28860
rect 13474 28800 13538 28804
rect 21422 28860 21486 28864
rect 21422 28804 21426 28860
rect 21426 28804 21482 28860
rect 21482 28804 21486 28860
rect 21422 28800 21486 28804
rect 21502 28860 21566 28864
rect 21502 28804 21506 28860
rect 21506 28804 21562 28860
rect 21562 28804 21566 28860
rect 21502 28800 21566 28804
rect 21582 28860 21646 28864
rect 21582 28804 21586 28860
rect 21586 28804 21642 28860
rect 21642 28804 21646 28860
rect 21582 28800 21646 28804
rect 21662 28860 21726 28864
rect 21662 28804 21666 28860
rect 21666 28804 21722 28860
rect 21722 28804 21726 28860
rect 21662 28800 21726 28804
rect 29610 28860 29674 28864
rect 29610 28804 29614 28860
rect 29614 28804 29670 28860
rect 29670 28804 29674 28860
rect 29610 28800 29674 28804
rect 29690 28860 29754 28864
rect 29690 28804 29694 28860
rect 29694 28804 29750 28860
rect 29750 28804 29754 28860
rect 29690 28800 29754 28804
rect 29770 28860 29834 28864
rect 29770 28804 29774 28860
rect 29774 28804 29830 28860
rect 29830 28804 29834 28860
rect 29770 28800 29834 28804
rect 29850 28860 29914 28864
rect 29850 28804 29854 28860
rect 29854 28804 29910 28860
rect 29910 28804 29914 28860
rect 29850 28800 29914 28804
rect 9140 28316 9204 28320
rect 9140 28260 9144 28316
rect 9144 28260 9200 28316
rect 9200 28260 9204 28316
rect 9140 28256 9204 28260
rect 9220 28316 9284 28320
rect 9220 28260 9224 28316
rect 9224 28260 9280 28316
rect 9280 28260 9284 28316
rect 9220 28256 9284 28260
rect 9300 28316 9364 28320
rect 9300 28260 9304 28316
rect 9304 28260 9360 28316
rect 9360 28260 9364 28316
rect 9300 28256 9364 28260
rect 9380 28316 9444 28320
rect 9380 28260 9384 28316
rect 9384 28260 9440 28316
rect 9440 28260 9444 28316
rect 9380 28256 9444 28260
rect 17328 28316 17392 28320
rect 17328 28260 17332 28316
rect 17332 28260 17388 28316
rect 17388 28260 17392 28316
rect 17328 28256 17392 28260
rect 17408 28316 17472 28320
rect 17408 28260 17412 28316
rect 17412 28260 17468 28316
rect 17468 28260 17472 28316
rect 17408 28256 17472 28260
rect 17488 28316 17552 28320
rect 17488 28260 17492 28316
rect 17492 28260 17548 28316
rect 17548 28260 17552 28316
rect 17488 28256 17552 28260
rect 17568 28316 17632 28320
rect 17568 28260 17572 28316
rect 17572 28260 17628 28316
rect 17628 28260 17632 28316
rect 17568 28256 17632 28260
rect 25516 28316 25580 28320
rect 25516 28260 25520 28316
rect 25520 28260 25576 28316
rect 25576 28260 25580 28316
rect 25516 28256 25580 28260
rect 25596 28316 25660 28320
rect 25596 28260 25600 28316
rect 25600 28260 25656 28316
rect 25656 28260 25660 28316
rect 25596 28256 25660 28260
rect 25676 28316 25740 28320
rect 25676 28260 25680 28316
rect 25680 28260 25736 28316
rect 25736 28260 25740 28316
rect 25676 28256 25740 28260
rect 25756 28316 25820 28320
rect 25756 28260 25760 28316
rect 25760 28260 25816 28316
rect 25816 28260 25820 28316
rect 25756 28256 25820 28260
rect 33704 28316 33768 28320
rect 33704 28260 33708 28316
rect 33708 28260 33764 28316
rect 33764 28260 33768 28316
rect 33704 28256 33768 28260
rect 33784 28316 33848 28320
rect 33784 28260 33788 28316
rect 33788 28260 33844 28316
rect 33844 28260 33848 28316
rect 33784 28256 33848 28260
rect 33864 28316 33928 28320
rect 33864 28260 33868 28316
rect 33868 28260 33924 28316
rect 33924 28260 33928 28316
rect 33864 28256 33928 28260
rect 33944 28316 34008 28320
rect 33944 28260 33948 28316
rect 33948 28260 34004 28316
rect 34004 28260 34008 28316
rect 33944 28256 34008 28260
rect 5046 27772 5110 27776
rect 5046 27716 5050 27772
rect 5050 27716 5106 27772
rect 5106 27716 5110 27772
rect 5046 27712 5110 27716
rect 5126 27772 5190 27776
rect 5126 27716 5130 27772
rect 5130 27716 5186 27772
rect 5186 27716 5190 27772
rect 5126 27712 5190 27716
rect 5206 27772 5270 27776
rect 5206 27716 5210 27772
rect 5210 27716 5266 27772
rect 5266 27716 5270 27772
rect 5206 27712 5270 27716
rect 5286 27772 5350 27776
rect 5286 27716 5290 27772
rect 5290 27716 5346 27772
rect 5346 27716 5350 27772
rect 5286 27712 5350 27716
rect 13234 27772 13298 27776
rect 13234 27716 13238 27772
rect 13238 27716 13294 27772
rect 13294 27716 13298 27772
rect 13234 27712 13298 27716
rect 13314 27772 13378 27776
rect 13314 27716 13318 27772
rect 13318 27716 13374 27772
rect 13374 27716 13378 27772
rect 13314 27712 13378 27716
rect 13394 27772 13458 27776
rect 13394 27716 13398 27772
rect 13398 27716 13454 27772
rect 13454 27716 13458 27772
rect 13394 27712 13458 27716
rect 13474 27772 13538 27776
rect 13474 27716 13478 27772
rect 13478 27716 13534 27772
rect 13534 27716 13538 27772
rect 13474 27712 13538 27716
rect 21422 27772 21486 27776
rect 21422 27716 21426 27772
rect 21426 27716 21482 27772
rect 21482 27716 21486 27772
rect 21422 27712 21486 27716
rect 21502 27772 21566 27776
rect 21502 27716 21506 27772
rect 21506 27716 21562 27772
rect 21562 27716 21566 27772
rect 21502 27712 21566 27716
rect 21582 27772 21646 27776
rect 21582 27716 21586 27772
rect 21586 27716 21642 27772
rect 21642 27716 21646 27772
rect 21582 27712 21646 27716
rect 21662 27772 21726 27776
rect 21662 27716 21666 27772
rect 21666 27716 21722 27772
rect 21722 27716 21726 27772
rect 21662 27712 21726 27716
rect 29610 27772 29674 27776
rect 29610 27716 29614 27772
rect 29614 27716 29670 27772
rect 29670 27716 29674 27772
rect 29610 27712 29674 27716
rect 29690 27772 29754 27776
rect 29690 27716 29694 27772
rect 29694 27716 29750 27772
rect 29750 27716 29754 27772
rect 29690 27712 29754 27716
rect 29770 27772 29834 27776
rect 29770 27716 29774 27772
rect 29774 27716 29830 27772
rect 29830 27716 29834 27772
rect 29770 27712 29834 27716
rect 29850 27772 29914 27776
rect 29850 27716 29854 27772
rect 29854 27716 29910 27772
rect 29910 27716 29914 27772
rect 29850 27712 29914 27716
rect 9140 27228 9204 27232
rect 9140 27172 9144 27228
rect 9144 27172 9200 27228
rect 9200 27172 9204 27228
rect 9140 27168 9204 27172
rect 9220 27228 9284 27232
rect 9220 27172 9224 27228
rect 9224 27172 9280 27228
rect 9280 27172 9284 27228
rect 9220 27168 9284 27172
rect 9300 27228 9364 27232
rect 9300 27172 9304 27228
rect 9304 27172 9360 27228
rect 9360 27172 9364 27228
rect 9300 27168 9364 27172
rect 9380 27228 9444 27232
rect 9380 27172 9384 27228
rect 9384 27172 9440 27228
rect 9440 27172 9444 27228
rect 9380 27168 9444 27172
rect 17328 27228 17392 27232
rect 17328 27172 17332 27228
rect 17332 27172 17388 27228
rect 17388 27172 17392 27228
rect 17328 27168 17392 27172
rect 17408 27228 17472 27232
rect 17408 27172 17412 27228
rect 17412 27172 17468 27228
rect 17468 27172 17472 27228
rect 17408 27168 17472 27172
rect 17488 27228 17552 27232
rect 17488 27172 17492 27228
rect 17492 27172 17548 27228
rect 17548 27172 17552 27228
rect 17488 27168 17552 27172
rect 17568 27228 17632 27232
rect 17568 27172 17572 27228
rect 17572 27172 17628 27228
rect 17628 27172 17632 27228
rect 17568 27168 17632 27172
rect 25516 27228 25580 27232
rect 25516 27172 25520 27228
rect 25520 27172 25576 27228
rect 25576 27172 25580 27228
rect 25516 27168 25580 27172
rect 25596 27228 25660 27232
rect 25596 27172 25600 27228
rect 25600 27172 25656 27228
rect 25656 27172 25660 27228
rect 25596 27168 25660 27172
rect 25676 27228 25740 27232
rect 25676 27172 25680 27228
rect 25680 27172 25736 27228
rect 25736 27172 25740 27228
rect 25676 27168 25740 27172
rect 25756 27228 25820 27232
rect 25756 27172 25760 27228
rect 25760 27172 25816 27228
rect 25816 27172 25820 27228
rect 25756 27168 25820 27172
rect 33704 27228 33768 27232
rect 33704 27172 33708 27228
rect 33708 27172 33764 27228
rect 33764 27172 33768 27228
rect 33704 27168 33768 27172
rect 33784 27228 33848 27232
rect 33784 27172 33788 27228
rect 33788 27172 33844 27228
rect 33844 27172 33848 27228
rect 33784 27168 33848 27172
rect 33864 27228 33928 27232
rect 33864 27172 33868 27228
rect 33868 27172 33924 27228
rect 33924 27172 33928 27228
rect 33864 27168 33928 27172
rect 33944 27228 34008 27232
rect 33944 27172 33948 27228
rect 33948 27172 34004 27228
rect 34004 27172 34008 27228
rect 33944 27168 34008 27172
rect 5046 26684 5110 26688
rect 5046 26628 5050 26684
rect 5050 26628 5106 26684
rect 5106 26628 5110 26684
rect 5046 26624 5110 26628
rect 5126 26684 5190 26688
rect 5126 26628 5130 26684
rect 5130 26628 5186 26684
rect 5186 26628 5190 26684
rect 5126 26624 5190 26628
rect 5206 26684 5270 26688
rect 5206 26628 5210 26684
rect 5210 26628 5266 26684
rect 5266 26628 5270 26684
rect 5206 26624 5270 26628
rect 5286 26684 5350 26688
rect 5286 26628 5290 26684
rect 5290 26628 5346 26684
rect 5346 26628 5350 26684
rect 5286 26624 5350 26628
rect 13234 26684 13298 26688
rect 13234 26628 13238 26684
rect 13238 26628 13294 26684
rect 13294 26628 13298 26684
rect 13234 26624 13298 26628
rect 13314 26684 13378 26688
rect 13314 26628 13318 26684
rect 13318 26628 13374 26684
rect 13374 26628 13378 26684
rect 13314 26624 13378 26628
rect 13394 26684 13458 26688
rect 13394 26628 13398 26684
rect 13398 26628 13454 26684
rect 13454 26628 13458 26684
rect 13394 26624 13458 26628
rect 13474 26684 13538 26688
rect 13474 26628 13478 26684
rect 13478 26628 13534 26684
rect 13534 26628 13538 26684
rect 13474 26624 13538 26628
rect 21422 26684 21486 26688
rect 21422 26628 21426 26684
rect 21426 26628 21482 26684
rect 21482 26628 21486 26684
rect 21422 26624 21486 26628
rect 21502 26684 21566 26688
rect 21502 26628 21506 26684
rect 21506 26628 21562 26684
rect 21562 26628 21566 26684
rect 21502 26624 21566 26628
rect 21582 26684 21646 26688
rect 21582 26628 21586 26684
rect 21586 26628 21642 26684
rect 21642 26628 21646 26684
rect 21582 26624 21646 26628
rect 21662 26684 21726 26688
rect 21662 26628 21666 26684
rect 21666 26628 21722 26684
rect 21722 26628 21726 26684
rect 21662 26624 21726 26628
rect 29610 26684 29674 26688
rect 29610 26628 29614 26684
rect 29614 26628 29670 26684
rect 29670 26628 29674 26684
rect 29610 26624 29674 26628
rect 29690 26684 29754 26688
rect 29690 26628 29694 26684
rect 29694 26628 29750 26684
rect 29750 26628 29754 26684
rect 29690 26624 29754 26628
rect 29770 26684 29834 26688
rect 29770 26628 29774 26684
rect 29774 26628 29830 26684
rect 29830 26628 29834 26684
rect 29770 26624 29834 26628
rect 29850 26684 29914 26688
rect 29850 26628 29854 26684
rect 29854 26628 29910 26684
rect 29910 26628 29914 26684
rect 29850 26624 29914 26628
rect 9140 26140 9204 26144
rect 9140 26084 9144 26140
rect 9144 26084 9200 26140
rect 9200 26084 9204 26140
rect 9140 26080 9204 26084
rect 9220 26140 9284 26144
rect 9220 26084 9224 26140
rect 9224 26084 9280 26140
rect 9280 26084 9284 26140
rect 9220 26080 9284 26084
rect 9300 26140 9364 26144
rect 9300 26084 9304 26140
rect 9304 26084 9360 26140
rect 9360 26084 9364 26140
rect 9300 26080 9364 26084
rect 9380 26140 9444 26144
rect 9380 26084 9384 26140
rect 9384 26084 9440 26140
rect 9440 26084 9444 26140
rect 9380 26080 9444 26084
rect 17328 26140 17392 26144
rect 17328 26084 17332 26140
rect 17332 26084 17388 26140
rect 17388 26084 17392 26140
rect 17328 26080 17392 26084
rect 17408 26140 17472 26144
rect 17408 26084 17412 26140
rect 17412 26084 17468 26140
rect 17468 26084 17472 26140
rect 17408 26080 17472 26084
rect 17488 26140 17552 26144
rect 17488 26084 17492 26140
rect 17492 26084 17548 26140
rect 17548 26084 17552 26140
rect 17488 26080 17552 26084
rect 17568 26140 17632 26144
rect 17568 26084 17572 26140
rect 17572 26084 17628 26140
rect 17628 26084 17632 26140
rect 17568 26080 17632 26084
rect 25516 26140 25580 26144
rect 25516 26084 25520 26140
rect 25520 26084 25576 26140
rect 25576 26084 25580 26140
rect 25516 26080 25580 26084
rect 25596 26140 25660 26144
rect 25596 26084 25600 26140
rect 25600 26084 25656 26140
rect 25656 26084 25660 26140
rect 25596 26080 25660 26084
rect 25676 26140 25740 26144
rect 25676 26084 25680 26140
rect 25680 26084 25736 26140
rect 25736 26084 25740 26140
rect 25676 26080 25740 26084
rect 25756 26140 25820 26144
rect 25756 26084 25760 26140
rect 25760 26084 25816 26140
rect 25816 26084 25820 26140
rect 25756 26080 25820 26084
rect 33704 26140 33768 26144
rect 33704 26084 33708 26140
rect 33708 26084 33764 26140
rect 33764 26084 33768 26140
rect 33704 26080 33768 26084
rect 33784 26140 33848 26144
rect 33784 26084 33788 26140
rect 33788 26084 33844 26140
rect 33844 26084 33848 26140
rect 33784 26080 33848 26084
rect 33864 26140 33928 26144
rect 33864 26084 33868 26140
rect 33868 26084 33924 26140
rect 33924 26084 33928 26140
rect 33864 26080 33928 26084
rect 33944 26140 34008 26144
rect 33944 26084 33948 26140
rect 33948 26084 34004 26140
rect 34004 26084 34008 26140
rect 33944 26080 34008 26084
rect 5046 25596 5110 25600
rect 5046 25540 5050 25596
rect 5050 25540 5106 25596
rect 5106 25540 5110 25596
rect 5046 25536 5110 25540
rect 5126 25596 5190 25600
rect 5126 25540 5130 25596
rect 5130 25540 5186 25596
rect 5186 25540 5190 25596
rect 5126 25536 5190 25540
rect 5206 25596 5270 25600
rect 5206 25540 5210 25596
rect 5210 25540 5266 25596
rect 5266 25540 5270 25596
rect 5206 25536 5270 25540
rect 5286 25596 5350 25600
rect 5286 25540 5290 25596
rect 5290 25540 5346 25596
rect 5346 25540 5350 25596
rect 5286 25536 5350 25540
rect 13234 25596 13298 25600
rect 13234 25540 13238 25596
rect 13238 25540 13294 25596
rect 13294 25540 13298 25596
rect 13234 25536 13298 25540
rect 13314 25596 13378 25600
rect 13314 25540 13318 25596
rect 13318 25540 13374 25596
rect 13374 25540 13378 25596
rect 13314 25536 13378 25540
rect 13394 25596 13458 25600
rect 13394 25540 13398 25596
rect 13398 25540 13454 25596
rect 13454 25540 13458 25596
rect 13394 25536 13458 25540
rect 13474 25596 13538 25600
rect 13474 25540 13478 25596
rect 13478 25540 13534 25596
rect 13534 25540 13538 25596
rect 13474 25536 13538 25540
rect 21422 25596 21486 25600
rect 21422 25540 21426 25596
rect 21426 25540 21482 25596
rect 21482 25540 21486 25596
rect 21422 25536 21486 25540
rect 21502 25596 21566 25600
rect 21502 25540 21506 25596
rect 21506 25540 21562 25596
rect 21562 25540 21566 25596
rect 21502 25536 21566 25540
rect 21582 25596 21646 25600
rect 21582 25540 21586 25596
rect 21586 25540 21642 25596
rect 21642 25540 21646 25596
rect 21582 25536 21646 25540
rect 21662 25596 21726 25600
rect 21662 25540 21666 25596
rect 21666 25540 21722 25596
rect 21722 25540 21726 25596
rect 21662 25536 21726 25540
rect 29610 25596 29674 25600
rect 29610 25540 29614 25596
rect 29614 25540 29670 25596
rect 29670 25540 29674 25596
rect 29610 25536 29674 25540
rect 29690 25596 29754 25600
rect 29690 25540 29694 25596
rect 29694 25540 29750 25596
rect 29750 25540 29754 25596
rect 29690 25536 29754 25540
rect 29770 25596 29834 25600
rect 29770 25540 29774 25596
rect 29774 25540 29830 25596
rect 29830 25540 29834 25596
rect 29770 25536 29834 25540
rect 29850 25596 29914 25600
rect 29850 25540 29854 25596
rect 29854 25540 29910 25596
rect 29910 25540 29914 25596
rect 29850 25536 29914 25540
rect 9140 25052 9204 25056
rect 9140 24996 9144 25052
rect 9144 24996 9200 25052
rect 9200 24996 9204 25052
rect 9140 24992 9204 24996
rect 9220 25052 9284 25056
rect 9220 24996 9224 25052
rect 9224 24996 9280 25052
rect 9280 24996 9284 25052
rect 9220 24992 9284 24996
rect 9300 25052 9364 25056
rect 9300 24996 9304 25052
rect 9304 24996 9360 25052
rect 9360 24996 9364 25052
rect 9300 24992 9364 24996
rect 9380 25052 9444 25056
rect 9380 24996 9384 25052
rect 9384 24996 9440 25052
rect 9440 24996 9444 25052
rect 9380 24992 9444 24996
rect 17328 25052 17392 25056
rect 17328 24996 17332 25052
rect 17332 24996 17388 25052
rect 17388 24996 17392 25052
rect 17328 24992 17392 24996
rect 17408 25052 17472 25056
rect 17408 24996 17412 25052
rect 17412 24996 17468 25052
rect 17468 24996 17472 25052
rect 17408 24992 17472 24996
rect 17488 25052 17552 25056
rect 17488 24996 17492 25052
rect 17492 24996 17548 25052
rect 17548 24996 17552 25052
rect 17488 24992 17552 24996
rect 17568 25052 17632 25056
rect 17568 24996 17572 25052
rect 17572 24996 17628 25052
rect 17628 24996 17632 25052
rect 17568 24992 17632 24996
rect 25516 25052 25580 25056
rect 25516 24996 25520 25052
rect 25520 24996 25576 25052
rect 25576 24996 25580 25052
rect 25516 24992 25580 24996
rect 25596 25052 25660 25056
rect 25596 24996 25600 25052
rect 25600 24996 25656 25052
rect 25656 24996 25660 25052
rect 25596 24992 25660 24996
rect 25676 25052 25740 25056
rect 25676 24996 25680 25052
rect 25680 24996 25736 25052
rect 25736 24996 25740 25052
rect 25676 24992 25740 24996
rect 25756 25052 25820 25056
rect 25756 24996 25760 25052
rect 25760 24996 25816 25052
rect 25816 24996 25820 25052
rect 25756 24992 25820 24996
rect 33704 25052 33768 25056
rect 33704 24996 33708 25052
rect 33708 24996 33764 25052
rect 33764 24996 33768 25052
rect 33704 24992 33768 24996
rect 33784 25052 33848 25056
rect 33784 24996 33788 25052
rect 33788 24996 33844 25052
rect 33844 24996 33848 25052
rect 33784 24992 33848 24996
rect 33864 25052 33928 25056
rect 33864 24996 33868 25052
rect 33868 24996 33924 25052
rect 33924 24996 33928 25052
rect 33864 24992 33928 24996
rect 33944 25052 34008 25056
rect 33944 24996 33948 25052
rect 33948 24996 34004 25052
rect 34004 24996 34008 25052
rect 33944 24992 34008 24996
rect 5046 24508 5110 24512
rect 5046 24452 5050 24508
rect 5050 24452 5106 24508
rect 5106 24452 5110 24508
rect 5046 24448 5110 24452
rect 5126 24508 5190 24512
rect 5126 24452 5130 24508
rect 5130 24452 5186 24508
rect 5186 24452 5190 24508
rect 5126 24448 5190 24452
rect 5206 24508 5270 24512
rect 5206 24452 5210 24508
rect 5210 24452 5266 24508
rect 5266 24452 5270 24508
rect 5206 24448 5270 24452
rect 5286 24508 5350 24512
rect 5286 24452 5290 24508
rect 5290 24452 5346 24508
rect 5346 24452 5350 24508
rect 5286 24448 5350 24452
rect 13234 24508 13298 24512
rect 13234 24452 13238 24508
rect 13238 24452 13294 24508
rect 13294 24452 13298 24508
rect 13234 24448 13298 24452
rect 13314 24508 13378 24512
rect 13314 24452 13318 24508
rect 13318 24452 13374 24508
rect 13374 24452 13378 24508
rect 13314 24448 13378 24452
rect 13394 24508 13458 24512
rect 13394 24452 13398 24508
rect 13398 24452 13454 24508
rect 13454 24452 13458 24508
rect 13394 24448 13458 24452
rect 13474 24508 13538 24512
rect 13474 24452 13478 24508
rect 13478 24452 13534 24508
rect 13534 24452 13538 24508
rect 13474 24448 13538 24452
rect 21422 24508 21486 24512
rect 21422 24452 21426 24508
rect 21426 24452 21482 24508
rect 21482 24452 21486 24508
rect 21422 24448 21486 24452
rect 21502 24508 21566 24512
rect 21502 24452 21506 24508
rect 21506 24452 21562 24508
rect 21562 24452 21566 24508
rect 21502 24448 21566 24452
rect 21582 24508 21646 24512
rect 21582 24452 21586 24508
rect 21586 24452 21642 24508
rect 21642 24452 21646 24508
rect 21582 24448 21646 24452
rect 21662 24508 21726 24512
rect 21662 24452 21666 24508
rect 21666 24452 21722 24508
rect 21722 24452 21726 24508
rect 21662 24448 21726 24452
rect 29610 24508 29674 24512
rect 29610 24452 29614 24508
rect 29614 24452 29670 24508
rect 29670 24452 29674 24508
rect 29610 24448 29674 24452
rect 29690 24508 29754 24512
rect 29690 24452 29694 24508
rect 29694 24452 29750 24508
rect 29750 24452 29754 24508
rect 29690 24448 29754 24452
rect 29770 24508 29834 24512
rect 29770 24452 29774 24508
rect 29774 24452 29830 24508
rect 29830 24452 29834 24508
rect 29770 24448 29834 24452
rect 29850 24508 29914 24512
rect 29850 24452 29854 24508
rect 29854 24452 29910 24508
rect 29910 24452 29914 24508
rect 29850 24448 29914 24452
rect 9140 23964 9204 23968
rect 9140 23908 9144 23964
rect 9144 23908 9200 23964
rect 9200 23908 9204 23964
rect 9140 23904 9204 23908
rect 9220 23964 9284 23968
rect 9220 23908 9224 23964
rect 9224 23908 9280 23964
rect 9280 23908 9284 23964
rect 9220 23904 9284 23908
rect 9300 23964 9364 23968
rect 9300 23908 9304 23964
rect 9304 23908 9360 23964
rect 9360 23908 9364 23964
rect 9300 23904 9364 23908
rect 9380 23964 9444 23968
rect 9380 23908 9384 23964
rect 9384 23908 9440 23964
rect 9440 23908 9444 23964
rect 9380 23904 9444 23908
rect 17328 23964 17392 23968
rect 17328 23908 17332 23964
rect 17332 23908 17388 23964
rect 17388 23908 17392 23964
rect 17328 23904 17392 23908
rect 17408 23964 17472 23968
rect 17408 23908 17412 23964
rect 17412 23908 17468 23964
rect 17468 23908 17472 23964
rect 17408 23904 17472 23908
rect 17488 23964 17552 23968
rect 17488 23908 17492 23964
rect 17492 23908 17548 23964
rect 17548 23908 17552 23964
rect 17488 23904 17552 23908
rect 17568 23964 17632 23968
rect 17568 23908 17572 23964
rect 17572 23908 17628 23964
rect 17628 23908 17632 23964
rect 17568 23904 17632 23908
rect 25516 23964 25580 23968
rect 25516 23908 25520 23964
rect 25520 23908 25576 23964
rect 25576 23908 25580 23964
rect 25516 23904 25580 23908
rect 25596 23964 25660 23968
rect 25596 23908 25600 23964
rect 25600 23908 25656 23964
rect 25656 23908 25660 23964
rect 25596 23904 25660 23908
rect 25676 23964 25740 23968
rect 25676 23908 25680 23964
rect 25680 23908 25736 23964
rect 25736 23908 25740 23964
rect 25676 23904 25740 23908
rect 25756 23964 25820 23968
rect 25756 23908 25760 23964
rect 25760 23908 25816 23964
rect 25816 23908 25820 23964
rect 25756 23904 25820 23908
rect 33704 23964 33768 23968
rect 33704 23908 33708 23964
rect 33708 23908 33764 23964
rect 33764 23908 33768 23964
rect 33704 23904 33768 23908
rect 33784 23964 33848 23968
rect 33784 23908 33788 23964
rect 33788 23908 33844 23964
rect 33844 23908 33848 23964
rect 33784 23904 33848 23908
rect 33864 23964 33928 23968
rect 33864 23908 33868 23964
rect 33868 23908 33924 23964
rect 33924 23908 33928 23964
rect 33864 23904 33928 23908
rect 33944 23964 34008 23968
rect 33944 23908 33948 23964
rect 33948 23908 34004 23964
rect 34004 23908 34008 23964
rect 33944 23904 34008 23908
rect 5046 23420 5110 23424
rect 5046 23364 5050 23420
rect 5050 23364 5106 23420
rect 5106 23364 5110 23420
rect 5046 23360 5110 23364
rect 5126 23420 5190 23424
rect 5126 23364 5130 23420
rect 5130 23364 5186 23420
rect 5186 23364 5190 23420
rect 5126 23360 5190 23364
rect 5206 23420 5270 23424
rect 5206 23364 5210 23420
rect 5210 23364 5266 23420
rect 5266 23364 5270 23420
rect 5206 23360 5270 23364
rect 5286 23420 5350 23424
rect 5286 23364 5290 23420
rect 5290 23364 5346 23420
rect 5346 23364 5350 23420
rect 5286 23360 5350 23364
rect 13234 23420 13298 23424
rect 13234 23364 13238 23420
rect 13238 23364 13294 23420
rect 13294 23364 13298 23420
rect 13234 23360 13298 23364
rect 13314 23420 13378 23424
rect 13314 23364 13318 23420
rect 13318 23364 13374 23420
rect 13374 23364 13378 23420
rect 13314 23360 13378 23364
rect 13394 23420 13458 23424
rect 13394 23364 13398 23420
rect 13398 23364 13454 23420
rect 13454 23364 13458 23420
rect 13394 23360 13458 23364
rect 13474 23420 13538 23424
rect 13474 23364 13478 23420
rect 13478 23364 13534 23420
rect 13534 23364 13538 23420
rect 13474 23360 13538 23364
rect 21422 23420 21486 23424
rect 21422 23364 21426 23420
rect 21426 23364 21482 23420
rect 21482 23364 21486 23420
rect 21422 23360 21486 23364
rect 21502 23420 21566 23424
rect 21502 23364 21506 23420
rect 21506 23364 21562 23420
rect 21562 23364 21566 23420
rect 21502 23360 21566 23364
rect 21582 23420 21646 23424
rect 21582 23364 21586 23420
rect 21586 23364 21642 23420
rect 21642 23364 21646 23420
rect 21582 23360 21646 23364
rect 21662 23420 21726 23424
rect 21662 23364 21666 23420
rect 21666 23364 21722 23420
rect 21722 23364 21726 23420
rect 21662 23360 21726 23364
rect 29610 23420 29674 23424
rect 29610 23364 29614 23420
rect 29614 23364 29670 23420
rect 29670 23364 29674 23420
rect 29610 23360 29674 23364
rect 29690 23420 29754 23424
rect 29690 23364 29694 23420
rect 29694 23364 29750 23420
rect 29750 23364 29754 23420
rect 29690 23360 29754 23364
rect 29770 23420 29834 23424
rect 29770 23364 29774 23420
rect 29774 23364 29830 23420
rect 29830 23364 29834 23420
rect 29770 23360 29834 23364
rect 29850 23420 29914 23424
rect 29850 23364 29854 23420
rect 29854 23364 29910 23420
rect 29910 23364 29914 23420
rect 29850 23360 29914 23364
rect 9140 22876 9204 22880
rect 9140 22820 9144 22876
rect 9144 22820 9200 22876
rect 9200 22820 9204 22876
rect 9140 22816 9204 22820
rect 9220 22876 9284 22880
rect 9220 22820 9224 22876
rect 9224 22820 9280 22876
rect 9280 22820 9284 22876
rect 9220 22816 9284 22820
rect 9300 22876 9364 22880
rect 9300 22820 9304 22876
rect 9304 22820 9360 22876
rect 9360 22820 9364 22876
rect 9300 22816 9364 22820
rect 9380 22876 9444 22880
rect 9380 22820 9384 22876
rect 9384 22820 9440 22876
rect 9440 22820 9444 22876
rect 9380 22816 9444 22820
rect 17328 22876 17392 22880
rect 17328 22820 17332 22876
rect 17332 22820 17388 22876
rect 17388 22820 17392 22876
rect 17328 22816 17392 22820
rect 17408 22876 17472 22880
rect 17408 22820 17412 22876
rect 17412 22820 17468 22876
rect 17468 22820 17472 22876
rect 17408 22816 17472 22820
rect 17488 22876 17552 22880
rect 17488 22820 17492 22876
rect 17492 22820 17548 22876
rect 17548 22820 17552 22876
rect 17488 22816 17552 22820
rect 17568 22876 17632 22880
rect 17568 22820 17572 22876
rect 17572 22820 17628 22876
rect 17628 22820 17632 22876
rect 17568 22816 17632 22820
rect 25516 22876 25580 22880
rect 25516 22820 25520 22876
rect 25520 22820 25576 22876
rect 25576 22820 25580 22876
rect 25516 22816 25580 22820
rect 25596 22876 25660 22880
rect 25596 22820 25600 22876
rect 25600 22820 25656 22876
rect 25656 22820 25660 22876
rect 25596 22816 25660 22820
rect 25676 22876 25740 22880
rect 25676 22820 25680 22876
rect 25680 22820 25736 22876
rect 25736 22820 25740 22876
rect 25676 22816 25740 22820
rect 25756 22876 25820 22880
rect 25756 22820 25760 22876
rect 25760 22820 25816 22876
rect 25816 22820 25820 22876
rect 25756 22816 25820 22820
rect 33704 22876 33768 22880
rect 33704 22820 33708 22876
rect 33708 22820 33764 22876
rect 33764 22820 33768 22876
rect 33704 22816 33768 22820
rect 33784 22876 33848 22880
rect 33784 22820 33788 22876
rect 33788 22820 33844 22876
rect 33844 22820 33848 22876
rect 33784 22816 33848 22820
rect 33864 22876 33928 22880
rect 33864 22820 33868 22876
rect 33868 22820 33924 22876
rect 33924 22820 33928 22876
rect 33864 22816 33928 22820
rect 33944 22876 34008 22880
rect 33944 22820 33948 22876
rect 33948 22820 34004 22876
rect 34004 22820 34008 22876
rect 33944 22816 34008 22820
rect 5046 22332 5110 22336
rect 5046 22276 5050 22332
rect 5050 22276 5106 22332
rect 5106 22276 5110 22332
rect 5046 22272 5110 22276
rect 5126 22332 5190 22336
rect 5126 22276 5130 22332
rect 5130 22276 5186 22332
rect 5186 22276 5190 22332
rect 5126 22272 5190 22276
rect 5206 22332 5270 22336
rect 5206 22276 5210 22332
rect 5210 22276 5266 22332
rect 5266 22276 5270 22332
rect 5206 22272 5270 22276
rect 5286 22332 5350 22336
rect 5286 22276 5290 22332
rect 5290 22276 5346 22332
rect 5346 22276 5350 22332
rect 5286 22272 5350 22276
rect 13234 22332 13298 22336
rect 13234 22276 13238 22332
rect 13238 22276 13294 22332
rect 13294 22276 13298 22332
rect 13234 22272 13298 22276
rect 13314 22332 13378 22336
rect 13314 22276 13318 22332
rect 13318 22276 13374 22332
rect 13374 22276 13378 22332
rect 13314 22272 13378 22276
rect 13394 22332 13458 22336
rect 13394 22276 13398 22332
rect 13398 22276 13454 22332
rect 13454 22276 13458 22332
rect 13394 22272 13458 22276
rect 13474 22332 13538 22336
rect 13474 22276 13478 22332
rect 13478 22276 13534 22332
rect 13534 22276 13538 22332
rect 13474 22272 13538 22276
rect 21422 22332 21486 22336
rect 21422 22276 21426 22332
rect 21426 22276 21482 22332
rect 21482 22276 21486 22332
rect 21422 22272 21486 22276
rect 21502 22332 21566 22336
rect 21502 22276 21506 22332
rect 21506 22276 21562 22332
rect 21562 22276 21566 22332
rect 21502 22272 21566 22276
rect 21582 22332 21646 22336
rect 21582 22276 21586 22332
rect 21586 22276 21642 22332
rect 21642 22276 21646 22332
rect 21582 22272 21646 22276
rect 21662 22332 21726 22336
rect 21662 22276 21666 22332
rect 21666 22276 21722 22332
rect 21722 22276 21726 22332
rect 21662 22272 21726 22276
rect 29610 22332 29674 22336
rect 29610 22276 29614 22332
rect 29614 22276 29670 22332
rect 29670 22276 29674 22332
rect 29610 22272 29674 22276
rect 29690 22332 29754 22336
rect 29690 22276 29694 22332
rect 29694 22276 29750 22332
rect 29750 22276 29754 22332
rect 29690 22272 29754 22276
rect 29770 22332 29834 22336
rect 29770 22276 29774 22332
rect 29774 22276 29830 22332
rect 29830 22276 29834 22332
rect 29770 22272 29834 22276
rect 29850 22332 29914 22336
rect 29850 22276 29854 22332
rect 29854 22276 29910 22332
rect 29910 22276 29914 22332
rect 29850 22272 29914 22276
rect 9140 21788 9204 21792
rect 9140 21732 9144 21788
rect 9144 21732 9200 21788
rect 9200 21732 9204 21788
rect 9140 21728 9204 21732
rect 9220 21788 9284 21792
rect 9220 21732 9224 21788
rect 9224 21732 9280 21788
rect 9280 21732 9284 21788
rect 9220 21728 9284 21732
rect 9300 21788 9364 21792
rect 9300 21732 9304 21788
rect 9304 21732 9360 21788
rect 9360 21732 9364 21788
rect 9300 21728 9364 21732
rect 9380 21788 9444 21792
rect 9380 21732 9384 21788
rect 9384 21732 9440 21788
rect 9440 21732 9444 21788
rect 9380 21728 9444 21732
rect 17328 21788 17392 21792
rect 17328 21732 17332 21788
rect 17332 21732 17388 21788
rect 17388 21732 17392 21788
rect 17328 21728 17392 21732
rect 17408 21788 17472 21792
rect 17408 21732 17412 21788
rect 17412 21732 17468 21788
rect 17468 21732 17472 21788
rect 17408 21728 17472 21732
rect 17488 21788 17552 21792
rect 17488 21732 17492 21788
rect 17492 21732 17548 21788
rect 17548 21732 17552 21788
rect 17488 21728 17552 21732
rect 17568 21788 17632 21792
rect 17568 21732 17572 21788
rect 17572 21732 17628 21788
rect 17628 21732 17632 21788
rect 17568 21728 17632 21732
rect 25516 21788 25580 21792
rect 25516 21732 25520 21788
rect 25520 21732 25576 21788
rect 25576 21732 25580 21788
rect 25516 21728 25580 21732
rect 25596 21788 25660 21792
rect 25596 21732 25600 21788
rect 25600 21732 25656 21788
rect 25656 21732 25660 21788
rect 25596 21728 25660 21732
rect 25676 21788 25740 21792
rect 25676 21732 25680 21788
rect 25680 21732 25736 21788
rect 25736 21732 25740 21788
rect 25676 21728 25740 21732
rect 25756 21788 25820 21792
rect 25756 21732 25760 21788
rect 25760 21732 25816 21788
rect 25816 21732 25820 21788
rect 25756 21728 25820 21732
rect 33704 21788 33768 21792
rect 33704 21732 33708 21788
rect 33708 21732 33764 21788
rect 33764 21732 33768 21788
rect 33704 21728 33768 21732
rect 33784 21788 33848 21792
rect 33784 21732 33788 21788
rect 33788 21732 33844 21788
rect 33844 21732 33848 21788
rect 33784 21728 33848 21732
rect 33864 21788 33928 21792
rect 33864 21732 33868 21788
rect 33868 21732 33924 21788
rect 33924 21732 33928 21788
rect 33864 21728 33928 21732
rect 33944 21788 34008 21792
rect 33944 21732 33948 21788
rect 33948 21732 34004 21788
rect 34004 21732 34008 21788
rect 33944 21728 34008 21732
rect 5046 21244 5110 21248
rect 5046 21188 5050 21244
rect 5050 21188 5106 21244
rect 5106 21188 5110 21244
rect 5046 21184 5110 21188
rect 5126 21244 5190 21248
rect 5126 21188 5130 21244
rect 5130 21188 5186 21244
rect 5186 21188 5190 21244
rect 5126 21184 5190 21188
rect 5206 21244 5270 21248
rect 5206 21188 5210 21244
rect 5210 21188 5266 21244
rect 5266 21188 5270 21244
rect 5206 21184 5270 21188
rect 5286 21244 5350 21248
rect 5286 21188 5290 21244
rect 5290 21188 5346 21244
rect 5346 21188 5350 21244
rect 5286 21184 5350 21188
rect 13234 21244 13298 21248
rect 13234 21188 13238 21244
rect 13238 21188 13294 21244
rect 13294 21188 13298 21244
rect 13234 21184 13298 21188
rect 13314 21244 13378 21248
rect 13314 21188 13318 21244
rect 13318 21188 13374 21244
rect 13374 21188 13378 21244
rect 13314 21184 13378 21188
rect 13394 21244 13458 21248
rect 13394 21188 13398 21244
rect 13398 21188 13454 21244
rect 13454 21188 13458 21244
rect 13394 21184 13458 21188
rect 13474 21244 13538 21248
rect 13474 21188 13478 21244
rect 13478 21188 13534 21244
rect 13534 21188 13538 21244
rect 13474 21184 13538 21188
rect 21422 21244 21486 21248
rect 21422 21188 21426 21244
rect 21426 21188 21482 21244
rect 21482 21188 21486 21244
rect 21422 21184 21486 21188
rect 21502 21244 21566 21248
rect 21502 21188 21506 21244
rect 21506 21188 21562 21244
rect 21562 21188 21566 21244
rect 21502 21184 21566 21188
rect 21582 21244 21646 21248
rect 21582 21188 21586 21244
rect 21586 21188 21642 21244
rect 21642 21188 21646 21244
rect 21582 21184 21646 21188
rect 21662 21244 21726 21248
rect 21662 21188 21666 21244
rect 21666 21188 21722 21244
rect 21722 21188 21726 21244
rect 21662 21184 21726 21188
rect 29610 21244 29674 21248
rect 29610 21188 29614 21244
rect 29614 21188 29670 21244
rect 29670 21188 29674 21244
rect 29610 21184 29674 21188
rect 29690 21244 29754 21248
rect 29690 21188 29694 21244
rect 29694 21188 29750 21244
rect 29750 21188 29754 21244
rect 29690 21184 29754 21188
rect 29770 21244 29834 21248
rect 29770 21188 29774 21244
rect 29774 21188 29830 21244
rect 29830 21188 29834 21244
rect 29770 21184 29834 21188
rect 29850 21244 29914 21248
rect 29850 21188 29854 21244
rect 29854 21188 29910 21244
rect 29910 21188 29914 21244
rect 29850 21184 29914 21188
rect 9140 20700 9204 20704
rect 9140 20644 9144 20700
rect 9144 20644 9200 20700
rect 9200 20644 9204 20700
rect 9140 20640 9204 20644
rect 9220 20700 9284 20704
rect 9220 20644 9224 20700
rect 9224 20644 9280 20700
rect 9280 20644 9284 20700
rect 9220 20640 9284 20644
rect 9300 20700 9364 20704
rect 9300 20644 9304 20700
rect 9304 20644 9360 20700
rect 9360 20644 9364 20700
rect 9300 20640 9364 20644
rect 9380 20700 9444 20704
rect 9380 20644 9384 20700
rect 9384 20644 9440 20700
rect 9440 20644 9444 20700
rect 9380 20640 9444 20644
rect 17328 20700 17392 20704
rect 17328 20644 17332 20700
rect 17332 20644 17388 20700
rect 17388 20644 17392 20700
rect 17328 20640 17392 20644
rect 17408 20700 17472 20704
rect 17408 20644 17412 20700
rect 17412 20644 17468 20700
rect 17468 20644 17472 20700
rect 17408 20640 17472 20644
rect 17488 20700 17552 20704
rect 17488 20644 17492 20700
rect 17492 20644 17548 20700
rect 17548 20644 17552 20700
rect 17488 20640 17552 20644
rect 17568 20700 17632 20704
rect 17568 20644 17572 20700
rect 17572 20644 17628 20700
rect 17628 20644 17632 20700
rect 17568 20640 17632 20644
rect 25516 20700 25580 20704
rect 25516 20644 25520 20700
rect 25520 20644 25576 20700
rect 25576 20644 25580 20700
rect 25516 20640 25580 20644
rect 25596 20700 25660 20704
rect 25596 20644 25600 20700
rect 25600 20644 25656 20700
rect 25656 20644 25660 20700
rect 25596 20640 25660 20644
rect 25676 20700 25740 20704
rect 25676 20644 25680 20700
rect 25680 20644 25736 20700
rect 25736 20644 25740 20700
rect 25676 20640 25740 20644
rect 25756 20700 25820 20704
rect 25756 20644 25760 20700
rect 25760 20644 25816 20700
rect 25816 20644 25820 20700
rect 25756 20640 25820 20644
rect 33704 20700 33768 20704
rect 33704 20644 33708 20700
rect 33708 20644 33764 20700
rect 33764 20644 33768 20700
rect 33704 20640 33768 20644
rect 33784 20700 33848 20704
rect 33784 20644 33788 20700
rect 33788 20644 33844 20700
rect 33844 20644 33848 20700
rect 33784 20640 33848 20644
rect 33864 20700 33928 20704
rect 33864 20644 33868 20700
rect 33868 20644 33924 20700
rect 33924 20644 33928 20700
rect 33864 20640 33928 20644
rect 33944 20700 34008 20704
rect 33944 20644 33948 20700
rect 33948 20644 34004 20700
rect 34004 20644 34008 20700
rect 33944 20640 34008 20644
rect 5046 20156 5110 20160
rect 5046 20100 5050 20156
rect 5050 20100 5106 20156
rect 5106 20100 5110 20156
rect 5046 20096 5110 20100
rect 5126 20156 5190 20160
rect 5126 20100 5130 20156
rect 5130 20100 5186 20156
rect 5186 20100 5190 20156
rect 5126 20096 5190 20100
rect 5206 20156 5270 20160
rect 5206 20100 5210 20156
rect 5210 20100 5266 20156
rect 5266 20100 5270 20156
rect 5206 20096 5270 20100
rect 5286 20156 5350 20160
rect 5286 20100 5290 20156
rect 5290 20100 5346 20156
rect 5346 20100 5350 20156
rect 5286 20096 5350 20100
rect 13234 20156 13298 20160
rect 13234 20100 13238 20156
rect 13238 20100 13294 20156
rect 13294 20100 13298 20156
rect 13234 20096 13298 20100
rect 13314 20156 13378 20160
rect 13314 20100 13318 20156
rect 13318 20100 13374 20156
rect 13374 20100 13378 20156
rect 13314 20096 13378 20100
rect 13394 20156 13458 20160
rect 13394 20100 13398 20156
rect 13398 20100 13454 20156
rect 13454 20100 13458 20156
rect 13394 20096 13458 20100
rect 13474 20156 13538 20160
rect 13474 20100 13478 20156
rect 13478 20100 13534 20156
rect 13534 20100 13538 20156
rect 13474 20096 13538 20100
rect 21422 20156 21486 20160
rect 21422 20100 21426 20156
rect 21426 20100 21482 20156
rect 21482 20100 21486 20156
rect 21422 20096 21486 20100
rect 21502 20156 21566 20160
rect 21502 20100 21506 20156
rect 21506 20100 21562 20156
rect 21562 20100 21566 20156
rect 21502 20096 21566 20100
rect 21582 20156 21646 20160
rect 21582 20100 21586 20156
rect 21586 20100 21642 20156
rect 21642 20100 21646 20156
rect 21582 20096 21646 20100
rect 21662 20156 21726 20160
rect 21662 20100 21666 20156
rect 21666 20100 21722 20156
rect 21722 20100 21726 20156
rect 21662 20096 21726 20100
rect 29610 20156 29674 20160
rect 29610 20100 29614 20156
rect 29614 20100 29670 20156
rect 29670 20100 29674 20156
rect 29610 20096 29674 20100
rect 29690 20156 29754 20160
rect 29690 20100 29694 20156
rect 29694 20100 29750 20156
rect 29750 20100 29754 20156
rect 29690 20096 29754 20100
rect 29770 20156 29834 20160
rect 29770 20100 29774 20156
rect 29774 20100 29830 20156
rect 29830 20100 29834 20156
rect 29770 20096 29834 20100
rect 29850 20156 29914 20160
rect 29850 20100 29854 20156
rect 29854 20100 29910 20156
rect 29910 20100 29914 20156
rect 29850 20096 29914 20100
rect 9140 19612 9204 19616
rect 9140 19556 9144 19612
rect 9144 19556 9200 19612
rect 9200 19556 9204 19612
rect 9140 19552 9204 19556
rect 9220 19612 9284 19616
rect 9220 19556 9224 19612
rect 9224 19556 9280 19612
rect 9280 19556 9284 19612
rect 9220 19552 9284 19556
rect 9300 19612 9364 19616
rect 9300 19556 9304 19612
rect 9304 19556 9360 19612
rect 9360 19556 9364 19612
rect 9300 19552 9364 19556
rect 9380 19612 9444 19616
rect 9380 19556 9384 19612
rect 9384 19556 9440 19612
rect 9440 19556 9444 19612
rect 9380 19552 9444 19556
rect 17328 19612 17392 19616
rect 17328 19556 17332 19612
rect 17332 19556 17388 19612
rect 17388 19556 17392 19612
rect 17328 19552 17392 19556
rect 17408 19612 17472 19616
rect 17408 19556 17412 19612
rect 17412 19556 17468 19612
rect 17468 19556 17472 19612
rect 17408 19552 17472 19556
rect 17488 19612 17552 19616
rect 17488 19556 17492 19612
rect 17492 19556 17548 19612
rect 17548 19556 17552 19612
rect 17488 19552 17552 19556
rect 17568 19612 17632 19616
rect 17568 19556 17572 19612
rect 17572 19556 17628 19612
rect 17628 19556 17632 19612
rect 17568 19552 17632 19556
rect 25516 19612 25580 19616
rect 25516 19556 25520 19612
rect 25520 19556 25576 19612
rect 25576 19556 25580 19612
rect 25516 19552 25580 19556
rect 25596 19612 25660 19616
rect 25596 19556 25600 19612
rect 25600 19556 25656 19612
rect 25656 19556 25660 19612
rect 25596 19552 25660 19556
rect 25676 19612 25740 19616
rect 25676 19556 25680 19612
rect 25680 19556 25736 19612
rect 25736 19556 25740 19612
rect 25676 19552 25740 19556
rect 25756 19612 25820 19616
rect 25756 19556 25760 19612
rect 25760 19556 25816 19612
rect 25816 19556 25820 19612
rect 25756 19552 25820 19556
rect 33704 19612 33768 19616
rect 33704 19556 33708 19612
rect 33708 19556 33764 19612
rect 33764 19556 33768 19612
rect 33704 19552 33768 19556
rect 33784 19612 33848 19616
rect 33784 19556 33788 19612
rect 33788 19556 33844 19612
rect 33844 19556 33848 19612
rect 33784 19552 33848 19556
rect 33864 19612 33928 19616
rect 33864 19556 33868 19612
rect 33868 19556 33924 19612
rect 33924 19556 33928 19612
rect 33864 19552 33928 19556
rect 33944 19612 34008 19616
rect 33944 19556 33948 19612
rect 33948 19556 34004 19612
rect 34004 19556 34008 19612
rect 33944 19552 34008 19556
rect 5046 19068 5110 19072
rect 5046 19012 5050 19068
rect 5050 19012 5106 19068
rect 5106 19012 5110 19068
rect 5046 19008 5110 19012
rect 5126 19068 5190 19072
rect 5126 19012 5130 19068
rect 5130 19012 5186 19068
rect 5186 19012 5190 19068
rect 5126 19008 5190 19012
rect 5206 19068 5270 19072
rect 5206 19012 5210 19068
rect 5210 19012 5266 19068
rect 5266 19012 5270 19068
rect 5206 19008 5270 19012
rect 5286 19068 5350 19072
rect 5286 19012 5290 19068
rect 5290 19012 5346 19068
rect 5346 19012 5350 19068
rect 5286 19008 5350 19012
rect 13234 19068 13298 19072
rect 13234 19012 13238 19068
rect 13238 19012 13294 19068
rect 13294 19012 13298 19068
rect 13234 19008 13298 19012
rect 13314 19068 13378 19072
rect 13314 19012 13318 19068
rect 13318 19012 13374 19068
rect 13374 19012 13378 19068
rect 13314 19008 13378 19012
rect 13394 19068 13458 19072
rect 13394 19012 13398 19068
rect 13398 19012 13454 19068
rect 13454 19012 13458 19068
rect 13394 19008 13458 19012
rect 13474 19068 13538 19072
rect 13474 19012 13478 19068
rect 13478 19012 13534 19068
rect 13534 19012 13538 19068
rect 13474 19008 13538 19012
rect 21422 19068 21486 19072
rect 21422 19012 21426 19068
rect 21426 19012 21482 19068
rect 21482 19012 21486 19068
rect 21422 19008 21486 19012
rect 21502 19068 21566 19072
rect 21502 19012 21506 19068
rect 21506 19012 21562 19068
rect 21562 19012 21566 19068
rect 21502 19008 21566 19012
rect 21582 19068 21646 19072
rect 21582 19012 21586 19068
rect 21586 19012 21642 19068
rect 21642 19012 21646 19068
rect 21582 19008 21646 19012
rect 21662 19068 21726 19072
rect 21662 19012 21666 19068
rect 21666 19012 21722 19068
rect 21722 19012 21726 19068
rect 21662 19008 21726 19012
rect 29610 19068 29674 19072
rect 29610 19012 29614 19068
rect 29614 19012 29670 19068
rect 29670 19012 29674 19068
rect 29610 19008 29674 19012
rect 29690 19068 29754 19072
rect 29690 19012 29694 19068
rect 29694 19012 29750 19068
rect 29750 19012 29754 19068
rect 29690 19008 29754 19012
rect 29770 19068 29834 19072
rect 29770 19012 29774 19068
rect 29774 19012 29830 19068
rect 29830 19012 29834 19068
rect 29770 19008 29834 19012
rect 29850 19068 29914 19072
rect 29850 19012 29854 19068
rect 29854 19012 29910 19068
rect 29910 19012 29914 19068
rect 29850 19008 29914 19012
rect 9140 18524 9204 18528
rect 9140 18468 9144 18524
rect 9144 18468 9200 18524
rect 9200 18468 9204 18524
rect 9140 18464 9204 18468
rect 9220 18524 9284 18528
rect 9220 18468 9224 18524
rect 9224 18468 9280 18524
rect 9280 18468 9284 18524
rect 9220 18464 9284 18468
rect 9300 18524 9364 18528
rect 9300 18468 9304 18524
rect 9304 18468 9360 18524
rect 9360 18468 9364 18524
rect 9300 18464 9364 18468
rect 9380 18524 9444 18528
rect 9380 18468 9384 18524
rect 9384 18468 9440 18524
rect 9440 18468 9444 18524
rect 9380 18464 9444 18468
rect 17328 18524 17392 18528
rect 17328 18468 17332 18524
rect 17332 18468 17388 18524
rect 17388 18468 17392 18524
rect 17328 18464 17392 18468
rect 17408 18524 17472 18528
rect 17408 18468 17412 18524
rect 17412 18468 17468 18524
rect 17468 18468 17472 18524
rect 17408 18464 17472 18468
rect 17488 18524 17552 18528
rect 17488 18468 17492 18524
rect 17492 18468 17548 18524
rect 17548 18468 17552 18524
rect 17488 18464 17552 18468
rect 17568 18524 17632 18528
rect 17568 18468 17572 18524
rect 17572 18468 17628 18524
rect 17628 18468 17632 18524
rect 17568 18464 17632 18468
rect 25516 18524 25580 18528
rect 25516 18468 25520 18524
rect 25520 18468 25576 18524
rect 25576 18468 25580 18524
rect 25516 18464 25580 18468
rect 25596 18524 25660 18528
rect 25596 18468 25600 18524
rect 25600 18468 25656 18524
rect 25656 18468 25660 18524
rect 25596 18464 25660 18468
rect 25676 18524 25740 18528
rect 25676 18468 25680 18524
rect 25680 18468 25736 18524
rect 25736 18468 25740 18524
rect 25676 18464 25740 18468
rect 25756 18524 25820 18528
rect 25756 18468 25760 18524
rect 25760 18468 25816 18524
rect 25816 18468 25820 18524
rect 25756 18464 25820 18468
rect 33704 18524 33768 18528
rect 33704 18468 33708 18524
rect 33708 18468 33764 18524
rect 33764 18468 33768 18524
rect 33704 18464 33768 18468
rect 33784 18524 33848 18528
rect 33784 18468 33788 18524
rect 33788 18468 33844 18524
rect 33844 18468 33848 18524
rect 33784 18464 33848 18468
rect 33864 18524 33928 18528
rect 33864 18468 33868 18524
rect 33868 18468 33924 18524
rect 33924 18468 33928 18524
rect 33864 18464 33928 18468
rect 33944 18524 34008 18528
rect 33944 18468 33948 18524
rect 33948 18468 34004 18524
rect 34004 18468 34008 18524
rect 33944 18464 34008 18468
rect 5046 17980 5110 17984
rect 5046 17924 5050 17980
rect 5050 17924 5106 17980
rect 5106 17924 5110 17980
rect 5046 17920 5110 17924
rect 5126 17980 5190 17984
rect 5126 17924 5130 17980
rect 5130 17924 5186 17980
rect 5186 17924 5190 17980
rect 5126 17920 5190 17924
rect 5206 17980 5270 17984
rect 5206 17924 5210 17980
rect 5210 17924 5266 17980
rect 5266 17924 5270 17980
rect 5206 17920 5270 17924
rect 5286 17980 5350 17984
rect 5286 17924 5290 17980
rect 5290 17924 5346 17980
rect 5346 17924 5350 17980
rect 5286 17920 5350 17924
rect 13234 17980 13298 17984
rect 13234 17924 13238 17980
rect 13238 17924 13294 17980
rect 13294 17924 13298 17980
rect 13234 17920 13298 17924
rect 13314 17980 13378 17984
rect 13314 17924 13318 17980
rect 13318 17924 13374 17980
rect 13374 17924 13378 17980
rect 13314 17920 13378 17924
rect 13394 17980 13458 17984
rect 13394 17924 13398 17980
rect 13398 17924 13454 17980
rect 13454 17924 13458 17980
rect 13394 17920 13458 17924
rect 13474 17980 13538 17984
rect 13474 17924 13478 17980
rect 13478 17924 13534 17980
rect 13534 17924 13538 17980
rect 13474 17920 13538 17924
rect 21422 17980 21486 17984
rect 21422 17924 21426 17980
rect 21426 17924 21482 17980
rect 21482 17924 21486 17980
rect 21422 17920 21486 17924
rect 21502 17980 21566 17984
rect 21502 17924 21506 17980
rect 21506 17924 21562 17980
rect 21562 17924 21566 17980
rect 21502 17920 21566 17924
rect 21582 17980 21646 17984
rect 21582 17924 21586 17980
rect 21586 17924 21642 17980
rect 21642 17924 21646 17980
rect 21582 17920 21646 17924
rect 21662 17980 21726 17984
rect 21662 17924 21666 17980
rect 21666 17924 21722 17980
rect 21722 17924 21726 17980
rect 21662 17920 21726 17924
rect 29610 17980 29674 17984
rect 29610 17924 29614 17980
rect 29614 17924 29670 17980
rect 29670 17924 29674 17980
rect 29610 17920 29674 17924
rect 29690 17980 29754 17984
rect 29690 17924 29694 17980
rect 29694 17924 29750 17980
rect 29750 17924 29754 17980
rect 29690 17920 29754 17924
rect 29770 17980 29834 17984
rect 29770 17924 29774 17980
rect 29774 17924 29830 17980
rect 29830 17924 29834 17980
rect 29770 17920 29834 17924
rect 29850 17980 29914 17984
rect 29850 17924 29854 17980
rect 29854 17924 29910 17980
rect 29910 17924 29914 17980
rect 29850 17920 29914 17924
rect 9140 17436 9204 17440
rect 9140 17380 9144 17436
rect 9144 17380 9200 17436
rect 9200 17380 9204 17436
rect 9140 17376 9204 17380
rect 9220 17436 9284 17440
rect 9220 17380 9224 17436
rect 9224 17380 9280 17436
rect 9280 17380 9284 17436
rect 9220 17376 9284 17380
rect 9300 17436 9364 17440
rect 9300 17380 9304 17436
rect 9304 17380 9360 17436
rect 9360 17380 9364 17436
rect 9300 17376 9364 17380
rect 9380 17436 9444 17440
rect 9380 17380 9384 17436
rect 9384 17380 9440 17436
rect 9440 17380 9444 17436
rect 9380 17376 9444 17380
rect 17328 17436 17392 17440
rect 17328 17380 17332 17436
rect 17332 17380 17388 17436
rect 17388 17380 17392 17436
rect 17328 17376 17392 17380
rect 17408 17436 17472 17440
rect 17408 17380 17412 17436
rect 17412 17380 17468 17436
rect 17468 17380 17472 17436
rect 17408 17376 17472 17380
rect 17488 17436 17552 17440
rect 17488 17380 17492 17436
rect 17492 17380 17548 17436
rect 17548 17380 17552 17436
rect 17488 17376 17552 17380
rect 17568 17436 17632 17440
rect 17568 17380 17572 17436
rect 17572 17380 17628 17436
rect 17628 17380 17632 17436
rect 17568 17376 17632 17380
rect 25516 17436 25580 17440
rect 25516 17380 25520 17436
rect 25520 17380 25576 17436
rect 25576 17380 25580 17436
rect 25516 17376 25580 17380
rect 25596 17436 25660 17440
rect 25596 17380 25600 17436
rect 25600 17380 25656 17436
rect 25656 17380 25660 17436
rect 25596 17376 25660 17380
rect 25676 17436 25740 17440
rect 25676 17380 25680 17436
rect 25680 17380 25736 17436
rect 25736 17380 25740 17436
rect 25676 17376 25740 17380
rect 25756 17436 25820 17440
rect 25756 17380 25760 17436
rect 25760 17380 25816 17436
rect 25816 17380 25820 17436
rect 25756 17376 25820 17380
rect 33704 17436 33768 17440
rect 33704 17380 33708 17436
rect 33708 17380 33764 17436
rect 33764 17380 33768 17436
rect 33704 17376 33768 17380
rect 33784 17436 33848 17440
rect 33784 17380 33788 17436
rect 33788 17380 33844 17436
rect 33844 17380 33848 17436
rect 33784 17376 33848 17380
rect 33864 17436 33928 17440
rect 33864 17380 33868 17436
rect 33868 17380 33924 17436
rect 33924 17380 33928 17436
rect 33864 17376 33928 17380
rect 33944 17436 34008 17440
rect 33944 17380 33948 17436
rect 33948 17380 34004 17436
rect 34004 17380 34008 17436
rect 33944 17376 34008 17380
rect 5046 16892 5110 16896
rect 5046 16836 5050 16892
rect 5050 16836 5106 16892
rect 5106 16836 5110 16892
rect 5046 16832 5110 16836
rect 5126 16892 5190 16896
rect 5126 16836 5130 16892
rect 5130 16836 5186 16892
rect 5186 16836 5190 16892
rect 5126 16832 5190 16836
rect 5206 16892 5270 16896
rect 5206 16836 5210 16892
rect 5210 16836 5266 16892
rect 5266 16836 5270 16892
rect 5206 16832 5270 16836
rect 5286 16892 5350 16896
rect 5286 16836 5290 16892
rect 5290 16836 5346 16892
rect 5346 16836 5350 16892
rect 5286 16832 5350 16836
rect 13234 16892 13298 16896
rect 13234 16836 13238 16892
rect 13238 16836 13294 16892
rect 13294 16836 13298 16892
rect 13234 16832 13298 16836
rect 13314 16892 13378 16896
rect 13314 16836 13318 16892
rect 13318 16836 13374 16892
rect 13374 16836 13378 16892
rect 13314 16832 13378 16836
rect 13394 16892 13458 16896
rect 13394 16836 13398 16892
rect 13398 16836 13454 16892
rect 13454 16836 13458 16892
rect 13394 16832 13458 16836
rect 13474 16892 13538 16896
rect 13474 16836 13478 16892
rect 13478 16836 13534 16892
rect 13534 16836 13538 16892
rect 13474 16832 13538 16836
rect 21422 16892 21486 16896
rect 21422 16836 21426 16892
rect 21426 16836 21482 16892
rect 21482 16836 21486 16892
rect 21422 16832 21486 16836
rect 21502 16892 21566 16896
rect 21502 16836 21506 16892
rect 21506 16836 21562 16892
rect 21562 16836 21566 16892
rect 21502 16832 21566 16836
rect 21582 16892 21646 16896
rect 21582 16836 21586 16892
rect 21586 16836 21642 16892
rect 21642 16836 21646 16892
rect 21582 16832 21646 16836
rect 21662 16892 21726 16896
rect 21662 16836 21666 16892
rect 21666 16836 21722 16892
rect 21722 16836 21726 16892
rect 21662 16832 21726 16836
rect 29610 16892 29674 16896
rect 29610 16836 29614 16892
rect 29614 16836 29670 16892
rect 29670 16836 29674 16892
rect 29610 16832 29674 16836
rect 29690 16892 29754 16896
rect 29690 16836 29694 16892
rect 29694 16836 29750 16892
rect 29750 16836 29754 16892
rect 29690 16832 29754 16836
rect 29770 16892 29834 16896
rect 29770 16836 29774 16892
rect 29774 16836 29830 16892
rect 29830 16836 29834 16892
rect 29770 16832 29834 16836
rect 29850 16892 29914 16896
rect 29850 16836 29854 16892
rect 29854 16836 29910 16892
rect 29910 16836 29914 16892
rect 29850 16832 29914 16836
rect 9140 16348 9204 16352
rect 9140 16292 9144 16348
rect 9144 16292 9200 16348
rect 9200 16292 9204 16348
rect 9140 16288 9204 16292
rect 9220 16348 9284 16352
rect 9220 16292 9224 16348
rect 9224 16292 9280 16348
rect 9280 16292 9284 16348
rect 9220 16288 9284 16292
rect 9300 16348 9364 16352
rect 9300 16292 9304 16348
rect 9304 16292 9360 16348
rect 9360 16292 9364 16348
rect 9300 16288 9364 16292
rect 9380 16348 9444 16352
rect 9380 16292 9384 16348
rect 9384 16292 9440 16348
rect 9440 16292 9444 16348
rect 9380 16288 9444 16292
rect 17328 16348 17392 16352
rect 17328 16292 17332 16348
rect 17332 16292 17388 16348
rect 17388 16292 17392 16348
rect 17328 16288 17392 16292
rect 17408 16348 17472 16352
rect 17408 16292 17412 16348
rect 17412 16292 17468 16348
rect 17468 16292 17472 16348
rect 17408 16288 17472 16292
rect 17488 16348 17552 16352
rect 17488 16292 17492 16348
rect 17492 16292 17548 16348
rect 17548 16292 17552 16348
rect 17488 16288 17552 16292
rect 17568 16348 17632 16352
rect 17568 16292 17572 16348
rect 17572 16292 17628 16348
rect 17628 16292 17632 16348
rect 17568 16288 17632 16292
rect 25516 16348 25580 16352
rect 25516 16292 25520 16348
rect 25520 16292 25576 16348
rect 25576 16292 25580 16348
rect 25516 16288 25580 16292
rect 25596 16348 25660 16352
rect 25596 16292 25600 16348
rect 25600 16292 25656 16348
rect 25656 16292 25660 16348
rect 25596 16288 25660 16292
rect 25676 16348 25740 16352
rect 25676 16292 25680 16348
rect 25680 16292 25736 16348
rect 25736 16292 25740 16348
rect 25676 16288 25740 16292
rect 25756 16348 25820 16352
rect 25756 16292 25760 16348
rect 25760 16292 25816 16348
rect 25816 16292 25820 16348
rect 25756 16288 25820 16292
rect 33704 16348 33768 16352
rect 33704 16292 33708 16348
rect 33708 16292 33764 16348
rect 33764 16292 33768 16348
rect 33704 16288 33768 16292
rect 33784 16348 33848 16352
rect 33784 16292 33788 16348
rect 33788 16292 33844 16348
rect 33844 16292 33848 16348
rect 33784 16288 33848 16292
rect 33864 16348 33928 16352
rect 33864 16292 33868 16348
rect 33868 16292 33924 16348
rect 33924 16292 33928 16348
rect 33864 16288 33928 16292
rect 33944 16348 34008 16352
rect 33944 16292 33948 16348
rect 33948 16292 34004 16348
rect 34004 16292 34008 16348
rect 33944 16288 34008 16292
rect 5046 15804 5110 15808
rect 5046 15748 5050 15804
rect 5050 15748 5106 15804
rect 5106 15748 5110 15804
rect 5046 15744 5110 15748
rect 5126 15804 5190 15808
rect 5126 15748 5130 15804
rect 5130 15748 5186 15804
rect 5186 15748 5190 15804
rect 5126 15744 5190 15748
rect 5206 15804 5270 15808
rect 5206 15748 5210 15804
rect 5210 15748 5266 15804
rect 5266 15748 5270 15804
rect 5206 15744 5270 15748
rect 5286 15804 5350 15808
rect 5286 15748 5290 15804
rect 5290 15748 5346 15804
rect 5346 15748 5350 15804
rect 5286 15744 5350 15748
rect 13234 15804 13298 15808
rect 13234 15748 13238 15804
rect 13238 15748 13294 15804
rect 13294 15748 13298 15804
rect 13234 15744 13298 15748
rect 13314 15804 13378 15808
rect 13314 15748 13318 15804
rect 13318 15748 13374 15804
rect 13374 15748 13378 15804
rect 13314 15744 13378 15748
rect 13394 15804 13458 15808
rect 13394 15748 13398 15804
rect 13398 15748 13454 15804
rect 13454 15748 13458 15804
rect 13394 15744 13458 15748
rect 13474 15804 13538 15808
rect 13474 15748 13478 15804
rect 13478 15748 13534 15804
rect 13534 15748 13538 15804
rect 13474 15744 13538 15748
rect 21422 15804 21486 15808
rect 21422 15748 21426 15804
rect 21426 15748 21482 15804
rect 21482 15748 21486 15804
rect 21422 15744 21486 15748
rect 21502 15804 21566 15808
rect 21502 15748 21506 15804
rect 21506 15748 21562 15804
rect 21562 15748 21566 15804
rect 21502 15744 21566 15748
rect 21582 15804 21646 15808
rect 21582 15748 21586 15804
rect 21586 15748 21642 15804
rect 21642 15748 21646 15804
rect 21582 15744 21646 15748
rect 21662 15804 21726 15808
rect 21662 15748 21666 15804
rect 21666 15748 21722 15804
rect 21722 15748 21726 15804
rect 21662 15744 21726 15748
rect 29610 15804 29674 15808
rect 29610 15748 29614 15804
rect 29614 15748 29670 15804
rect 29670 15748 29674 15804
rect 29610 15744 29674 15748
rect 29690 15804 29754 15808
rect 29690 15748 29694 15804
rect 29694 15748 29750 15804
rect 29750 15748 29754 15804
rect 29690 15744 29754 15748
rect 29770 15804 29834 15808
rect 29770 15748 29774 15804
rect 29774 15748 29830 15804
rect 29830 15748 29834 15804
rect 29770 15744 29834 15748
rect 29850 15804 29914 15808
rect 29850 15748 29854 15804
rect 29854 15748 29910 15804
rect 29910 15748 29914 15804
rect 29850 15744 29914 15748
rect 9140 15260 9204 15264
rect 9140 15204 9144 15260
rect 9144 15204 9200 15260
rect 9200 15204 9204 15260
rect 9140 15200 9204 15204
rect 9220 15260 9284 15264
rect 9220 15204 9224 15260
rect 9224 15204 9280 15260
rect 9280 15204 9284 15260
rect 9220 15200 9284 15204
rect 9300 15260 9364 15264
rect 9300 15204 9304 15260
rect 9304 15204 9360 15260
rect 9360 15204 9364 15260
rect 9300 15200 9364 15204
rect 9380 15260 9444 15264
rect 9380 15204 9384 15260
rect 9384 15204 9440 15260
rect 9440 15204 9444 15260
rect 9380 15200 9444 15204
rect 17328 15260 17392 15264
rect 17328 15204 17332 15260
rect 17332 15204 17388 15260
rect 17388 15204 17392 15260
rect 17328 15200 17392 15204
rect 17408 15260 17472 15264
rect 17408 15204 17412 15260
rect 17412 15204 17468 15260
rect 17468 15204 17472 15260
rect 17408 15200 17472 15204
rect 17488 15260 17552 15264
rect 17488 15204 17492 15260
rect 17492 15204 17548 15260
rect 17548 15204 17552 15260
rect 17488 15200 17552 15204
rect 17568 15260 17632 15264
rect 17568 15204 17572 15260
rect 17572 15204 17628 15260
rect 17628 15204 17632 15260
rect 17568 15200 17632 15204
rect 25516 15260 25580 15264
rect 25516 15204 25520 15260
rect 25520 15204 25576 15260
rect 25576 15204 25580 15260
rect 25516 15200 25580 15204
rect 25596 15260 25660 15264
rect 25596 15204 25600 15260
rect 25600 15204 25656 15260
rect 25656 15204 25660 15260
rect 25596 15200 25660 15204
rect 25676 15260 25740 15264
rect 25676 15204 25680 15260
rect 25680 15204 25736 15260
rect 25736 15204 25740 15260
rect 25676 15200 25740 15204
rect 25756 15260 25820 15264
rect 25756 15204 25760 15260
rect 25760 15204 25816 15260
rect 25816 15204 25820 15260
rect 25756 15200 25820 15204
rect 33704 15260 33768 15264
rect 33704 15204 33708 15260
rect 33708 15204 33764 15260
rect 33764 15204 33768 15260
rect 33704 15200 33768 15204
rect 33784 15260 33848 15264
rect 33784 15204 33788 15260
rect 33788 15204 33844 15260
rect 33844 15204 33848 15260
rect 33784 15200 33848 15204
rect 33864 15260 33928 15264
rect 33864 15204 33868 15260
rect 33868 15204 33924 15260
rect 33924 15204 33928 15260
rect 33864 15200 33928 15204
rect 33944 15260 34008 15264
rect 33944 15204 33948 15260
rect 33948 15204 34004 15260
rect 34004 15204 34008 15260
rect 33944 15200 34008 15204
rect 5046 14716 5110 14720
rect 5046 14660 5050 14716
rect 5050 14660 5106 14716
rect 5106 14660 5110 14716
rect 5046 14656 5110 14660
rect 5126 14716 5190 14720
rect 5126 14660 5130 14716
rect 5130 14660 5186 14716
rect 5186 14660 5190 14716
rect 5126 14656 5190 14660
rect 5206 14716 5270 14720
rect 5206 14660 5210 14716
rect 5210 14660 5266 14716
rect 5266 14660 5270 14716
rect 5206 14656 5270 14660
rect 5286 14716 5350 14720
rect 5286 14660 5290 14716
rect 5290 14660 5346 14716
rect 5346 14660 5350 14716
rect 5286 14656 5350 14660
rect 13234 14716 13298 14720
rect 13234 14660 13238 14716
rect 13238 14660 13294 14716
rect 13294 14660 13298 14716
rect 13234 14656 13298 14660
rect 13314 14716 13378 14720
rect 13314 14660 13318 14716
rect 13318 14660 13374 14716
rect 13374 14660 13378 14716
rect 13314 14656 13378 14660
rect 13394 14716 13458 14720
rect 13394 14660 13398 14716
rect 13398 14660 13454 14716
rect 13454 14660 13458 14716
rect 13394 14656 13458 14660
rect 13474 14716 13538 14720
rect 13474 14660 13478 14716
rect 13478 14660 13534 14716
rect 13534 14660 13538 14716
rect 13474 14656 13538 14660
rect 21422 14716 21486 14720
rect 21422 14660 21426 14716
rect 21426 14660 21482 14716
rect 21482 14660 21486 14716
rect 21422 14656 21486 14660
rect 21502 14716 21566 14720
rect 21502 14660 21506 14716
rect 21506 14660 21562 14716
rect 21562 14660 21566 14716
rect 21502 14656 21566 14660
rect 21582 14716 21646 14720
rect 21582 14660 21586 14716
rect 21586 14660 21642 14716
rect 21642 14660 21646 14716
rect 21582 14656 21646 14660
rect 21662 14716 21726 14720
rect 21662 14660 21666 14716
rect 21666 14660 21722 14716
rect 21722 14660 21726 14716
rect 21662 14656 21726 14660
rect 29610 14716 29674 14720
rect 29610 14660 29614 14716
rect 29614 14660 29670 14716
rect 29670 14660 29674 14716
rect 29610 14656 29674 14660
rect 29690 14716 29754 14720
rect 29690 14660 29694 14716
rect 29694 14660 29750 14716
rect 29750 14660 29754 14716
rect 29690 14656 29754 14660
rect 29770 14716 29834 14720
rect 29770 14660 29774 14716
rect 29774 14660 29830 14716
rect 29830 14660 29834 14716
rect 29770 14656 29834 14660
rect 29850 14716 29914 14720
rect 29850 14660 29854 14716
rect 29854 14660 29910 14716
rect 29910 14660 29914 14716
rect 29850 14656 29914 14660
rect 9140 14172 9204 14176
rect 9140 14116 9144 14172
rect 9144 14116 9200 14172
rect 9200 14116 9204 14172
rect 9140 14112 9204 14116
rect 9220 14172 9284 14176
rect 9220 14116 9224 14172
rect 9224 14116 9280 14172
rect 9280 14116 9284 14172
rect 9220 14112 9284 14116
rect 9300 14172 9364 14176
rect 9300 14116 9304 14172
rect 9304 14116 9360 14172
rect 9360 14116 9364 14172
rect 9300 14112 9364 14116
rect 9380 14172 9444 14176
rect 9380 14116 9384 14172
rect 9384 14116 9440 14172
rect 9440 14116 9444 14172
rect 9380 14112 9444 14116
rect 17328 14172 17392 14176
rect 17328 14116 17332 14172
rect 17332 14116 17388 14172
rect 17388 14116 17392 14172
rect 17328 14112 17392 14116
rect 17408 14172 17472 14176
rect 17408 14116 17412 14172
rect 17412 14116 17468 14172
rect 17468 14116 17472 14172
rect 17408 14112 17472 14116
rect 17488 14172 17552 14176
rect 17488 14116 17492 14172
rect 17492 14116 17548 14172
rect 17548 14116 17552 14172
rect 17488 14112 17552 14116
rect 17568 14172 17632 14176
rect 17568 14116 17572 14172
rect 17572 14116 17628 14172
rect 17628 14116 17632 14172
rect 17568 14112 17632 14116
rect 25516 14172 25580 14176
rect 25516 14116 25520 14172
rect 25520 14116 25576 14172
rect 25576 14116 25580 14172
rect 25516 14112 25580 14116
rect 25596 14172 25660 14176
rect 25596 14116 25600 14172
rect 25600 14116 25656 14172
rect 25656 14116 25660 14172
rect 25596 14112 25660 14116
rect 25676 14172 25740 14176
rect 25676 14116 25680 14172
rect 25680 14116 25736 14172
rect 25736 14116 25740 14172
rect 25676 14112 25740 14116
rect 25756 14172 25820 14176
rect 25756 14116 25760 14172
rect 25760 14116 25816 14172
rect 25816 14116 25820 14172
rect 25756 14112 25820 14116
rect 33704 14172 33768 14176
rect 33704 14116 33708 14172
rect 33708 14116 33764 14172
rect 33764 14116 33768 14172
rect 33704 14112 33768 14116
rect 33784 14172 33848 14176
rect 33784 14116 33788 14172
rect 33788 14116 33844 14172
rect 33844 14116 33848 14172
rect 33784 14112 33848 14116
rect 33864 14172 33928 14176
rect 33864 14116 33868 14172
rect 33868 14116 33924 14172
rect 33924 14116 33928 14172
rect 33864 14112 33928 14116
rect 33944 14172 34008 14176
rect 33944 14116 33948 14172
rect 33948 14116 34004 14172
rect 34004 14116 34008 14172
rect 33944 14112 34008 14116
rect 5046 13628 5110 13632
rect 5046 13572 5050 13628
rect 5050 13572 5106 13628
rect 5106 13572 5110 13628
rect 5046 13568 5110 13572
rect 5126 13628 5190 13632
rect 5126 13572 5130 13628
rect 5130 13572 5186 13628
rect 5186 13572 5190 13628
rect 5126 13568 5190 13572
rect 5206 13628 5270 13632
rect 5206 13572 5210 13628
rect 5210 13572 5266 13628
rect 5266 13572 5270 13628
rect 5206 13568 5270 13572
rect 5286 13628 5350 13632
rect 5286 13572 5290 13628
rect 5290 13572 5346 13628
rect 5346 13572 5350 13628
rect 5286 13568 5350 13572
rect 13234 13628 13298 13632
rect 13234 13572 13238 13628
rect 13238 13572 13294 13628
rect 13294 13572 13298 13628
rect 13234 13568 13298 13572
rect 13314 13628 13378 13632
rect 13314 13572 13318 13628
rect 13318 13572 13374 13628
rect 13374 13572 13378 13628
rect 13314 13568 13378 13572
rect 13394 13628 13458 13632
rect 13394 13572 13398 13628
rect 13398 13572 13454 13628
rect 13454 13572 13458 13628
rect 13394 13568 13458 13572
rect 13474 13628 13538 13632
rect 13474 13572 13478 13628
rect 13478 13572 13534 13628
rect 13534 13572 13538 13628
rect 13474 13568 13538 13572
rect 21422 13628 21486 13632
rect 21422 13572 21426 13628
rect 21426 13572 21482 13628
rect 21482 13572 21486 13628
rect 21422 13568 21486 13572
rect 21502 13628 21566 13632
rect 21502 13572 21506 13628
rect 21506 13572 21562 13628
rect 21562 13572 21566 13628
rect 21502 13568 21566 13572
rect 21582 13628 21646 13632
rect 21582 13572 21586 13628
rect 21586 13572 21642 13628
rect 21642 13572 21646 13628
rect 21582 13568 21646 13572
rect 21662 13628 21726 13632
rect 21662 13572 21666 13628
rect 21666 13572 21722 13628
rect 21722 13572 21726 13628
rect 21662 13568 21726 13572
rect 29610 13628 29674 13632
rect 29610 13572 29614 13628
rect 29614 13572 29670 13628
rect 29670 13572 29674 13628
rect 29610 13568 29674 13572
rect 29690 13628 29754 13632
rect 29690 13572 29694 13628
rect 29694 13572 29750 13628
rect 29750 13572 29754 13628
rect 29690 13568 29754 13572
rect 29770 13628 29834 13632
rect 29770 13572 29774 13628
rect 29774 13572 29830 13628
rect 29830 13572 29834 13628
rect 29770 13568 29834 13572
rect 29850 13628 29914 13632
rect 29850 13572 29854 13628
rect 29854 13572 29910 13628
rect 29910 13572 29914 13628
rect 29850 13568 29914 13572
rect 9140 13084 9204 13088
rect 9140 13028 9144 13084
rect 9144 13028 9200 13084
rect 9200 13028 9204 13084
rect 9140 13024 9204 13028
rect 9220 13084 9284 13088
rect 9220 13028 9224 13084
rect 9224 13028 9280 13084
rect 9280 13028 9284 13084
rect 9220 13024 9284 13028
rect 9300 13084 9364 13088
rect 9300 13028 9304 13084
rect 9304 13028 9360 13084
rect 9360 13028 9364 13084
rect 9300 13024 9364 13028
rect 9380 13084 9444 13088
rect 9380 13028 9384 13084
rect 9384 13028 9440 13084
rect 9440 13028 9444 13084
rect 9380 13024 9444 13028
rect 17328 13084 17392 13088
rect 17328 13028 17332 13084
rect 17332 13028 17388 13084
rect 17388 13028 17392 13084
rect 17328 13024 17392 13028
rect 17408 13084 17472 13088
rect 17408 13028 17412 13084
rect 17412 13028 17468 13084
rect 17468 13028 17472 13084
rect 17408 13024 17472 13028
rect 17488 13084 17552 13088
rect 17488 13028 17492 13084
rect 17492 13028 17548 13084
rect 17548 13028 17552 13084
rect 17488 13024 17552 13028
rect 17568 13084 17632 13088
rect 17568 13028 17572 13084
rect 17572 13028 17628 13084
rect 17628 13028 17632 13084
rect 17568 13024 17632 13028
rect 25516 13084 25580 13088
rect 25516 13028 25520 13084
rect 25520 13028 25576 13084
rect 25576 13028 25580 13084
rect 25516 13024 25580 13028
rect 25596 13084 25660 13088
rect 25596 13028 25600 13084
rect 25600 13028 25656 13084
rect 25656 13028 25660 13084
rect 25596 13024 25660 13028
rect 25676 13084 25740 13088
rect 25676 13028 25680 13084
rect 25680 13028 25736 13084
rect 25736 13028 25740 13084
rect 25676 13024 25740 13028
rect 25756 13084 25820 13088
rect 25756 13028 25760 13084
rect 25760 13028 25816 13084
rect 25816 13028 25820 13084
rect 25756 13024 25820 13028
rect 33704 13084 33768 13088
rect 33704 13028 33708 13084
rect 33708 13028 33764 13084
rect 33764 13028 33768 13084
rect 33704 13024 33768 13028
rect 33784 13084 33848 13088
rect 33784 13028 33788 13084
rect 33788 13028 33844 13084
rect 33844 13028 33848 13084
rect 33784 13024 33848 13028
rect 33864 13084 33928 13088
rect 33864 13028 33868 13084
rect 33868 13028 33924 13084
rect 33924 13028 33928 13084
rect 33864 13024 33928 13028
rect 33944 13084 34008 13088
rect 33944 13028 33948 13084
rect 33948 13028 34004 13084
rect 34004 13028 34008 13084
rect 33944 13024 34008 13028
rect 5046 12540 5110 12544
rect 5046 12484 5050 12540
rect 5050 12484 5106 12540
rect 5106 12484 5110 12540
rect 5046 12480 5110 12484
rect 5126 12540 5190 12544
rect 5126 12484 5130 12540
rect 5130 12484 5186 12540
rect 5186 12484 5190 12540
rect 5126 12480 5190 12484
rect 5206 12540 5270 12544
rect 5206 12484 5210 12540
rect 5210 12484 5266 12540
rect 5266 12484 5270 12540
rect 5206 12480 5270 12484
rect 5286 12540 5350 12544
rect 5286 12484 5290 12540
rect 5290 12484 5346 12540
rect 5346 12484 5350 12540
rect 5286 12480 5350 12484
rect 13234 12540 13298 12544
rect 13234 12484 13238 12540
rect 13238 12484 13294 12540
rect 13294 12484 13298 12540
rect 13234 12480 13298 12484
rect 13314 12540 13378 12544
rect 13314 12484 13318 12540
rect 13318 12484 13374 12540
rect 13374 12484 13378 12540
rect 13314 12480 13378 12484
rect 13394 12540 13458 12544
rect 13394 12484 13398 12540
rect 13398 12484 13454 12540
rect 13454 12484 13458 12540
rect 13394 12480 13458 12484
rect 13474 12540 13538 12544
rect 13474 12484 13478 12540
rect 13478 12484 13534 12540
rect 13534 12484 13538 12540
rect 13474 12480 13538 12484
rect 21422 12540 21486 12544
rect 21422 12484 21426 12540
rect 21426 12484 21482 12540
rect 21482 12484 21486 12540
rect 21422 12480 21486 12484
rect 21502 12540 21566 12544
rect 21502 12484 21506 12540
rect 21506 12484 21562 12540
rect 21562 12484 21566 12540
rect 21502 12480 21566 12484
rect 21582 12540 21646 12544
rect 21582 12484 21586 12540
rect 21586 12484 21642 12540
rect 21642 12484 21646 12540
rect 21582 12480 21646 12484
rect 21662 12540 21726 12544
rect 21662 12484 21666 12540
rect 21666 12484 21722 12540
rect 21722 12484 21726 12540
rect 21662 12480 21726 12484
rect 29610 12540 29674 12544
rect 29610 12484 29614 12540
rect 29614 12484 29670 12540
rect 29670 12484 29674 12540
rect 29610 12480 29674 12484
rect 29690 12540 29754 12544
rect 29690 12484 29694 12540
rect 29694 12484 29750 12540
rect 29750 12484 29754 12540
rect 29690 12480 29754 12484
rect 29770 12540 29834 12544
rect 29770 12484 29774 12540
rect 29774 12484 29830 12540
rect 29830 12484 29834 12540
rect 29770 12480 29834 12484
rect 29850 12540 29914 12544
rect 29850 12484 29854 12540
rect 29854 12484 29910 12540
rect 29910 12484 29914 12540
rect 29850 12480 29914 12484
rect 9140 11996 9204 12000
rect 9140 11940 9144 11996
rect 9144 11940 9200 11996
rect 9200 11940 9204 11996
rect 9140 11936 9204 11940
rect 9220 11996 9284 12000
rect 9220 11940 9224 11996
rect 9224 11940 9280 11996
rect 9280 11940 9284 11996
rect 9220 11936 9284 11940
rect 9300 11996 9364 12000
rect 9300 11940 9304 11996
rect 9304 11940 9360 11996
rect 9360 11940 9364 11996
rect 9300 11936 9364 11940
rect 9380 11996 9444 12000
rect 9380 11940 9384 11996
rect 9384 11940 9440 11996
rect 9440 11940 9444 11996
rect 9380 11936 9444 11940
rect 17328 11996 17392 12000
rect 17328 11940 17332 11996
rect 17332 11940 17388 11996
rect 17388 11940 17392 11996
rect 17328 11936 17392 11940
rect 17408 11996 17472 12000
rect 17408 11940 17412 11996
rect 17412 11940 17468 11996
rect 17468 11940 17472 11996
rect 17408 11936 17472 11940
rect 17488 11996 17552 12000
rect 17488 11940 17492 11996
rect 17492 11940 17548 11996
rect 17548 11940 17552 11996
rect 17488 11936 17552 11940
rect 17568 11996 17632 12000
rect 17568 11940 17572 11996
rect 17572 11940 17628 11996
rect 17628 11940 17632 11996
rect 17568 11936 17632 11940
rect 25516 11996 25580 12000
rect 25516 11940 25520 11996
rect 25520 11940 25576 11996
rect 25576 11940 25580 11996
rect 25516 11936 25580 11940
rect 25596 11996 25660 12000
rect 25596 11940 25600 11996
rect 25600 11940 25656 11996
rect 25656 11940 25660 11996
rect 25596 11936 25660 11940
rect 25676 11996 25740 12000
rect 25676 11940 25680 11996
rect 25680 11940 25736 11996
rect 25736 11940 25740 11996
rect 25676 11936 25740 11940
rect 25756 11996 25820 12000
rect 25756 11940 25760 11996
rect 25760 11940 25816 11996
rect 25816 11940 25820 11996
rect 25756 11936 25820 11940
rect 33704 11996 33768 12000
rect 33704 11940 33708 11996
rect 33708 11940 33764 11996
rect 33764 11940 33768 11996
rect 33704 11936 33768 11940
rect 33784 11996 33848 12000
rect 33784 11940 33788 11996
rect 33788 11940 33844 11996
rect 33844 11940 33848 11996
rect 33784 11936 33848 11940
rect 33864 11996 33928 12000
rect 33864 11940 33868 11996
rect 33868 11940 33924 11996
rect 33924 11940 33928 11996
rect 33864 11936 33928 11940
rect 33944 11996 34008 12000
rect 33944 11940 33948 11996
rect 33948 11940 34004 11996
rect 34004 11940 34008 11996
rect 33944 11936 34008 11940
rect 5046 11452 5110 11456
rect 5046 11396 5050 11452
rect 5050 11396 5106 11452
rect 5106 11396 5110 11452
rect 5046 11392 5110 11396
rect 5126 11452 5190 11456
rect 5126 11396 5130 11452
rect 5130 11396 5186 11452
rect 5186 11396 5190 11452
rect 5126 11392 5190 11396
rect 5206 11452 5270 11456
rect 5206 11396 5210 11452
rect 5210 11396 5266 11452
rect 5266 11396 5270 11452
rect 5206 11392 5270 11396
rect 5286 11452 5350 11456
rect 5286 11396 5290 11452
rect 5290 11396 5346 11452
rect 5346 11396 5350 11452
rect 5286 11392 5350 11396
rect 13234 11452 13298 11456
rect 13234 11396 13238 11452
rect 13238 11396 13294 11452
rect 13294 11396 13298 11452
rect 13234 11392 13298 11396
rect 13314 11452 13378 11456
rect 13314 11396 13318 11452
rect 13318 11396 13374 11452
rect 13374 11396 13378 11452
rect 13314 11392 13378 11396
rect 13394 11452 13458 11456
rect 13394 11396 13398 11452
rect 13398 11396 13454 11452
rect 13454 11396 13458 11452
rect 13394 11392 13458 11396
rect 13474 11452 13538 11456
rect 13474 11396 13478 11452
rect 13478 11396 13534 11452
rect 13534 11396 13538 11452
rect 13474 11392 13538 11396
rect 21422 11452 21486 11456
rect 21422 11396 21426 11452
rect 21426 11396 21482 11452
rect 21482 11396 21486 11452
rect 21422 11392 21486 11396
rect 21502 11452 21566 11456
rect 21502 11396 21506 11452
rect 21506 11396 21562 11452
rect 21562 11396 21566 11452
rect 21502 11392 21566 11396
rect 21582 11452 21646 11456
rect 21582 11396 21586 11452
rect 21586 11396 21642 11452
rect 21642 11396 21646 11452
rect 21582 11392 21646 11396
rect 21662 11452 21726 11456
rect 21662 11396 21666 11452
rect 21666 11396 21722 11452
rect 21722 11396 21726 11452
rect 21662 11392 21726 11396
rect 29610 11452 29674 11456
rect 29610 11396 29614 11452
rect 29614 11396 29670 11452
rect 29670 11396 29674 11452
rect 29610 11392 29674 11396
rect 29690 11452 29754 11456
rect 29690 11396 29694 11452
rect 29694 11396 29750 11452
rect 29750 11396 29754 11452
rect 29690 11392 29754 11396
rect 29770 11452 29834 11456
rect 29770 11396 29774 11452
rect 29774 11396 29830 11452
rect 29830 11396 29834 11452
rect 29770 11392 29834 11396
rect 29850 11452 29914 11456
rect 29850 11396 29854 11452
rect 29854 11396 29910 11452
rect 29910 11396 29914 11452
rect 29850 11392 29914 11396
rect 9140 10908 9204 10912
rect 9140 10852 9144 10908
rect 9144 10852 9200 10908
rect 9200 10852 9204 10908
rect 9140 10848 9204 10852
rect 9220 10908 9284 10912
rect 9220 10852 9224 10908
rect 9224 10852 9280 10908
rect 9280 10852 9284 10908
rect 9220 10848 9284 10852
rect 9300 10908 9364 10912
rect 9300 10852 9304 10908
rect 9304 10852 9360 10908
rect 9360 10852 9364 10908
rect 9300 10848 9364 10852
rect 9380 10908 9444 10912
rect 9380 10852 9384 10908
rect 9384 10852 9440 10908
rect 9440 10852 9444 10908
rect 9380 10848 9444 10852
rect 17328 10908 17392 10912
rect 17328 10852 17332 10908
rect 17332 10852 17388 10908
rect 17388 10852 17392 10908
rect 17328 10848 17392 10852
rect 17408 10908 17472 10912
rect 17408 10852 17412 10908
rect 17412 10852 17468 10908
rect 17468 10852 17472 10908
rect 17408 10848 17472 10852
rect 17488 10908 17552 10912
rect 17488 10852 17492 10908
rect 17492 10852 17548 10908
rect 17548 10852 17552 10908
rect 17488 10848 17552 10852
rect 17568 10908 17632 10912
rect 17568 10852 17572 10908
rect 17572 10852 17628 10908
rect 17628 10852 17632 10908
rect 17568 10848 17632 10852
rect 25516 10908 25580 10912
rect 25516 10852 25520 10908
rect 25520 10852 25576 10908
rect 25576 10852 25580 10908
rect 25516 10848 25580 10852
rect 25596 10908 25660 10912
rect 25596 10852 25600 10908
rect 25600 10852 25656 10908
rect 25656 10852 25660 10908
rect 25596 10848 25660 10852
rect 25676 10908 25740 10912
rect 25676 10852 25680 10908
rect 25680 10852 25736 10908
rect 25736 10852 25740 10908
rect 25676 10848 25740 10852
rect 25756 10908 25820 10912
rect 25756 10852 25760 10908
rect 25760 10852 25816 10908
rect 25816 10852 25820 10908
rect 25756 10848 25820 10852
rect 33704 10908 33768 10912
rect 33704 10852 33708 10908
rect 33708 10852 33764 10908
rect 33764 10852 33768 10908
rect 33704 10848 33768 10852
rect 33784 10908 33848 10912
rect 33784 10852 33788 10908
rect 33788 10852 33844 10908
rect 33844 10852 33848 10908
rect 33784 10848 33848 10852
rect 33864 10908 33928 10912
rect 33864 10852 33868 10908
rect 33868 10852 33924 10908
rect 33924 10852 33928 10908
rect 33864 10848 33928 10852
rect 33944 10908 34008 10912
rect 33944 10852 33948 10908
rect 33948 10852 34004 10908
rect 34004 10852 34008 10908
rect 33944 10848 34008 10852
rect 5046 10364 5110 10368
rect 5046 10308 5050 10364
rect 5050 10308 5106 10364
rect 5106 10308 5110 10364
rect 5046 10304 5110 10308
rect 5126 10364 5190 10368
rect 5126 10308 5130 10364
rect 5130 10308 5186 10364
rect 5186 10308 5190 10364
rect 5126 10304 5190 10308
rect 5206 10364 5270 10368
rect 5206 10308 5210 10364
rect 5210 10308 5266 10364
rect 5266 10308 5270 10364
rect 5206 10304 5270 10308
rect 5286 10364 5350 10368
rect 5286 10308 5290 10364
rect 5290 10308 5346 10364
rect 5346 10308 5350 10364
rect 5286 10304 5350 10308
rect 13234 10364 13298 10368
rect 13234 10308 13238 10364
rect 13238 10308 13294 10364
rect 13294 10308 13298 10364
rect 13234 10304 13298 10308
rect 13314 10364 13378 10368
rect 13314 10308 13318 10364
rect 13318 10308 13374 10364
rect 13374 10308 13378 10364
rect 13314 10304 13378 10308
rect 13394 10364 13458 10368
rect 13394 10308 13398 10364
rect 13398 10308 13454 10364
rect 13454 10308 13458 10364
rect 13394 10304 13458 10308
rect 13474 10364 13538 10368
rect 13474 10308 13478 10364
rect 13478 10308 13534 10364
rect 13534 10308 13538 10364
rect 13474 10304 13538 10308
rect 21422 10364 21486 10368
rect 21422 10308 21426 10364
rect 21426 10308 21482 10364
rect 21482 10308 21486 10364
rect 21422 10304 21486 10308
rect 21502 10364 21566 10368
rect 21502 10308 21506 10364
rect 21506 10308 21562 10364
rect 21562 10308 21566 10364
rect 21502 10304 21566 10308
rect 21582 10364 21646 10368
rect 21582 10308 21586 10364
rect 21586 10308 21642 10364
rect 21642 10308 21646 10364
rect 21582 10304 21646 10308
rect 21662 10364 21726 10368
rect 21662 10308 21666 10364
rect 21666 10308 21722 10364
rect 21722 10308 21726 10364
rect 21662 10304 21726 10308
rect 29610 10364 29674 10368
rect 29610 10308 29614 10364
rect 29614 10308 29670 10364
rect 29670 10308 29674 10364
rect 29610 10304 29674 10308
rect 29690 10364 29754 10368
rect 29690 10308 29694 10364
rect 29694 10308 29750 10364
rect 29750 10308 29754 10364
rect 29690 10304 29754 10308
rect 29770 10364 29834 10368
rect 29770 10308 29774 10364
rect 29774 10308 29830 10364
rect 29830 10308 29834 10364
rect 29770 10304 29834 10308
rect 29850 10364 29914 10368
rect 29850 10308 29854 10364
rect 29854 10308 29910 10364
rect 29910 10308 29914 10364
rect 29850 10304 29914 10308
rect 9140 9820 9204 9824
rect 9140 9764 9144 9820
rect 9144 9764 9200 9820
rect 9200 9764 9204 9820
rect 9140 9760 9204 9764
rect 9220 9820 9284 9824
rect 9220 9764 9224 9820
rect 9224 9764 9280 9820
rect 9280 9764 9284 9820
rect 9220 9760 9284 9764
rect 9300 9820 9364 9824
rect 9300 9764 9304 9820
rect 9304 9764 9360 9820
rect 9360 9764 9364 9820
rect 9300 9760 9364 9764
rect 9380 9820 9444 9824
rect 9380 9764 9384 9820
rect 9384 9764 9440 9820
rect 9440 9764 9444 9820
rect 9380 9760 9444 9764
rect 17328 9820 17392 9824
rect 17328 9764 17332 9820
rect 17332 9764 17388 9820
rect 17388 9764 17392 9820
rect 17328 9760 17392 9764
rect 17408 9820 17472 9824
rect 17408 9764 17412 9820
rect 17412 9764 17468 9820
rect 17468 9764 17472 9820
rect 17408 9760 17472 9764
rect 17488 9820 17552 9824
rect 17488 9764 17492 9820
rect 17492 9764 17548 9820
rect 17548 9764 17552 9820
rect 17488 9760 17552 9764
rect 17568 9820 17632 9824
rect 17568 9764 17572 9820
rect 17572 9764 17628 9820
rect 17628 9764 17632 9820
rect 17568 9760 17632 9764
rect 25516 9820 25580 9824
rect 25516 9764 25520 9820
rect 25520 9764 25576 9820
rect 25576 9764 25580 9820
rect 25516 9760 25580 9764
rect 25596 9820 25660 9824
rect 25596 9764 25600 9820
rect 25600 9764 25656 9820
rect 25656 9764 25660 9820
rect 25596 9760 25660 9764
rect 25676 9820 25740 9824
rect 25676 9764 25680 9820
rect 25680 9764 25736 9820
rect 25736 9764 25740 9820
rect 25676 9760 25740 9764
rect 25756 9820 25820 9824
rect 25756 9764 25760 9820
rect 25760 9764 25816 9820
rect 25816 9764 25820 9820
rect 25756 9760 25820 9764
rect 33704 9820 33768 9824
rect 33704 9764 33708 9820
rect 33708 9764 33764 9820
rect 33764 9764 33768 9820
rect 33704 9760 33768 9764
rect 33784 9820 33848 9824
rect 33784 9764 33788 9820
rect 33788 9764 33844 9820
rect 33844 9764 33848 9820
rect 33784 9760 33848 9764
rect 33864 9820 33928 9824
rect 33864 9764 33868 9820
rect 33868 9764 33924 9820
rect 33924 9764 33928 9820
rect 33864 9760 33928 9764
rect 33944 9820 34008 9824
rect 33944 9764 33948 9820
rect 33948 9764 34004 9820
rect 34004 9764 34008 9820
rect 33944 9760 34008 9764
rect 5046 9276 5110 9280
rect 5046 9220 5050 9276
rect 5050 9220 5106 9276
rect 5106 9220 5110 9276
rect 5046 9216 5110 9220
rect 5126 9276 5190 9280
rect 5126 9220 5130 9276
rect 5130 9220 5186 9276
rect 5186 9220 5190 9276
rect 5126 9216 5190 9220
rect 5206 9276 5270 9280
rect 5206 9220 5210 9276
rect 5210 9220 5266 9276
rect 5266 9220 5270 9276
rect 5206 9216 5270 9220
rect 5286 9276 5350 9280
rect 5286 9220 5290 9276
rect 5290 9220 5346 9276
rect 5346 9220 5350 9276
rect 5286 9216 5350 9220
rect 13234 9276 13298 9280
rect 13234 9220 13238 9276
rect 13238 9220 13294 9276
rect 13294 9220 13298 9276
rect 13234 9216 13298 9220
rect 13314 9276 13378 9280
rect 13314 9220 13318 9276
rect 13318 9220 13374 9276
rect 13374 9220 13378 9276
rect 13314 9216 13378 9220
rect 13394 9276 13458 9280
rect 13394 9220 13398 9276
rect 13398 9220 13454 9276
rect 13454 9220 13458 9276
rect 13394 9216 13458 9220
rect 13474 9276 13538 9280
rect 13474 9220 13478 9276
rect 13478 9220 13534 9276
rect 13534 9220 13538 9276
rect 13474 9216 13538 9220
rect 21422 9276 21486 9280
rect 21422 9220 21426 9276
rect 21426 9220 21482 9276
rect 21482 9220 21486 9276
rect 21422 9216 21486 9220
rect 21502 9276 21566 9280
rect 21502 9220 21506 9276
rect 21506 9220 21562 9276
rect 21562 9220 21566 9276
rect 21502 9216 21566 9220
rect 21582 9276 21646 9280
rect 21582 9220 21586 9276
rect 21586 9220 21642 9276
rect 21642 9220 21646 9276
rect 21582 9216 21646 9220
rect 21662 9276 21726 9280
rect 21662 9220 21666 9276
rect 21666 9220 21722 9276
rect 21722 9220 21726 9276
rect 21662 9216 21726 9220
rect 29610 9276 29674 9280
rect 29610 9220 29614 9276
rect 29614 9220 29670 9276
rect 29670 9220 29674 9276
rect 29610 9216 29674 9220
rect 29690 9276 29754 9280
rect 29690 9220 29694 9276
rect 29694 9220 29750 9276
rect 29750 9220 29754 9276
rect 29690 9216 29754 9220
rect 29770 9276 29834 9280
rect 29770 9220 29774 9276
rect 29774 9220 29830 9276
rect 29830 9220 29834 9276
rect 29770 9216 29834 9220
rect 29850 9276 29914 9280
rect 29850 9220 29854 9276
rect 29854 9220 29910 9276
rect 29910 9220 29914 9276
rect 29850 9216 29914 9220
rect 9140 8732 9204 8736
rect 9140 8676 9144 8732
rect 9144 8676 9200 8732
rect 9200 8676 9204 8732
rect 9140 8672 9204 8676
rect 9220 8732 9284 8736
rect 9220 8676 9224 8732
rect 9224 8676 9280 8732
rect 9280 8676 9284 8732
rect 9220 8672 9284 8676
rect 9300 8732 9364 8736
rect 9300 8676 9304 8732
rect 9304 8676 9360 8732
rect 9360 8676 9364 8732
rect 9300 8672 9364 8676
rect 9380 8732 9444 8736
rect 9380 8676 9384 8732
rect 9384 8676 9440 8732
rect 9440 8676 9444 8732
rect 9380 8672 9444 8676
rect 17328 8732 17392 8736
rect 17328 8676 17332 8732
rect 17332 8676 17388 8732
rect 17388 8676 17392 8732
rect 17328 8672 17392 8676
rect 17408 8732 17472 8736
rect 17408 8676 17412 8732
rect 17412 8676 17468 8732
rect 17468 8676 17472 8732
rect 17408 8672 17472 8676
rect 17488 8732 17552 8736
rect 17488 8676 17492 8732
rect 17492 8676 17548 8732
rect 17548 8676 17552 8732
rect 17488 8672 17552 8676
rect 17568 8732 17632 8736
rect 17568 8676 17572 8732
rect 17572 8676 17628 8732
rect 17628 8676 17632 8732
rect 17568 8672 17632 8676
rect 25516 8732 25580 8736
rect 25516 8676 25520 8732
rect 25520 8676 25576 8732
rect 25576 8676 25580 8732
rect 25516 8672 25580 8676
rect 25596 8732 25660 8736
rect 25596 8676 25600 8732
rect 25600 8676 25656 8732
rect 25656 8676 25660 8732
rect 25596 8672 25660 8676
rect 25676 8732 25740 8736
rect 25676 8676 25680 8732
rect 25680 8676 25736 8732
rect 25736 8676 25740 8732
rect 25676 8672 25740 8676
rect 25756 8732 25820 8736
rect 25756 8676 25760 8732
rect 25760 8676 25816 8732
rect 25816 8676 25820 8732
rect 25756 8672 25820 8676
rect 33704 8732 33768 8736
rect 33704 8676 33708 8732
rect 33708 8676 33764 8732
rect 33764 8676 33768 8732
rect 33704 8672 33768 8676
rect 33784 8732 33848 8736
rect 33784 8676 33788 8732
rect 33788 8676 33844 8732
rect 33844 8676 33848 8732
rect 33784 8672 33848 8676
rect 33864 8732 33928 8736
rect 33864 8676 33868 8732
rect 33868 8676 33924 8732
rect 33924 8676 33928 8732
rect 33864 8672 33928 8676
rect 33944 8732 34008 8736
rect 33944 8676 33948 8732
rect 33948 8676 34004 8732
rect 34004 8676 34008 8732
rect 33944 8672 34008 8676
rect 5046 8188 5110 8192
rect 5046 8132 5050 8188
rect 5050 8132 5106 8188
rect 5106 8132 5110 8188
rect 5046 8128 5110 8132
rect 5126 8188 5190 8192
rect 5126 8132 5130 8188
rect 5130 8132 5186 8188
rect 5186 8132 5190 8188
rect 5126 8128 5190 8132
rect 5206 8188 5270 8192
rect 5206 8132 5210 8188
rect 5210 8132 5266 8188
rect 5266 8132 5270 8188
rect 5206 8128 5270 8132
rect 5286 8188 5350 8192
rect 5286 8132 5290 8188
rect 5290 8132 5346 8188
rect 5346 8132 5350 8188
rect 5286 8128 5350 8132
rect 13234 8188 13298 8192
rect 13234 8132 13238 8188
rect 13238 8132 13294 8188
rect 13294 8132 13298 8188
rect 13234 8128 13298 8132
rect 13314 8188 13378 8192
rect 13314 8132 13318 8188
rect 13318 8132 13374 8188
rect 13374 8132 13378 8188
rect 13314 8128 13378 8132
rect 13394 8188 13458 8192
rect 13394 8132 13398 8188
rect 13398 8132 13454 8188
rect 13454 8132 13458 8188
rect 13394 8128 13458 8132
rect 13474 8188 13538 8192
rect 13474 8132 13478 8188
rect 13478 8132 13534 8188
rect 13534 8132 13538 8188
rect 13474 8128 13538 8132
rect 21422 8188 21486 8192
rect 21422 8132 21426 8188
rect 21426 8132 21482 8188
rect 21482 8132 21486 8188
rect 21422 8128 21486 8132
rect 21502 8188 21566 8192
rect 21502 8132 21506 8188
rect 21506 8132 21562 8188
rect 21562 8132 21566 8188
rect 21502 8128 21566 8132
rect 21582 8188 21646 8192
rect 21582 8132 21586 8188
rect 21586 8132 21642 8188
rect 21642 8132 21646 8188
rect 21582 8128 21646 8132
rect 21662 8188 21726 8192
rect 21662 8132 21666 8188
rect 21666 8132 21722 8188
rect 21722 8132 21726 8188
rect 21662 8128 21726 8132
rect 29610 8188 29674 8192
rect 29610 8132 29614 8188
rect 29614 8132 29670 8188
rect 29670 8132 29674 8188
rect 29610 8128 29674 8132
rect 29690 8188 29754 8192
rect 29690 8132 29694 8188
rect 29694 8132 29750 8188
rect 29750 8132 29754 8188
rect 29690 8128 29754 8132
rect 29770 8188 29834 8192
rect 29770 8132 29774 8188
rect 29774 8132 29830 8188
rect 29830 8132 29834 8188
rect 29770 8128 29834 8132
rect 29850 8188 29914 8192
rect 29850 8132 29854 8188
rect 29854 8132 29910 8188
rect 29910 8132 29914 8188
rect 29850 8128 29914 8132
rect 9140 7644 9204 7648
rect 9140 7588 9144 7644
rect 9144 7588 9200 7644
rect 9200 7588 9204 7644
rect 9140 7584 9204 7588
rect 9220 7644 9284 7648
rect 9220 7588 9224 7644
rect 9224 7588 9280 7644
rect 9280 7588 9284 7644
rect 9220 7584 9284 7588
rect 9300 7644 9364 7648
rect 9300 7588 9304 7644
rect 9304 7588 9360 7644
rect 9360 7588 9364 7644
rect 9300 7584 9364 7588
rect 9380 7644 9444 7648
rect 9380 7588 9384 7644
rect 9384 7588 9440 7644
rect 9440 7588 9444 7644
rect 9380 7584 9444 7588
rect 17328 7644 17392 7648
rect 17328 7588 17332 7644
rect 17332 7588 17388 7644
rect 17388 7588 17392 7644
rect 17328 7584 17392 7588
rect 17408 7644 17472 7648
rect 17408 7588 17412 7644
rect 17412 7588 17468 7644
rect 17468 7588 17472 7644
rect 17408 7584 17472 7588
rect 17488 7644 17552 7648
rect 17488 7588 17492 7644
rect 17492 7588 17548 7644
rect 17548 7588 17552 7644
rect 17488 7584 17552 7588
rect 17568 7644 17632 7648
rect 17568 7588 17572 7644
rect 17572 7588 17628 7644
rect 17628 7588 17632 7644
rect 17568 7584 17632 7588
rect 25516 7644 25580 7648
rect 25516 7588 25520 7644
rect 25520 7588 25576 7644
rect 25576 7588 25580 7644
rect 25516 7584 25580 7588
rect 25596 7644 25660 7648
rect 25596 7588 25600 7644
rect 25600 7588 25656 7644
rect 25656 7588 25660 7644
rect 25596 7584 25660 7588
rect 25676 7644 25740 7648
rect 25676 7588 25680 7644
rect 25680 7588 25736 7644
rect 25736 7588 25740 7644
rect 25676 7584 25740 7588
rect 25756 7644 25820 7648
rect 25756 7588 25760 7644
rect 25760 7588 25816 7644
rect 25816 7588 25820 7644
rect 25756 7584 25820 7588
rect 33704 7644 33768 7648
rect 33704 7588 33708 7644
rect 33708 7588 33764 7644
rect 33764 7588 33768 7644
rect 33704 7584 33768 7588
rect 33784 7644 33848 7648
rect 33784 7588 33788 7644
rect 33788 7588 33844 7644
rect 33844 7588 33848 7644
rect 33784 7584 33848 7588
rect 33864 7644 33928 7648
rect 33864 7588 33868 7644
rect 33868 7588 33924 7644
rect 33924 7588 33928 7644
rect 33864 7584 33928 7588
rect 33944 7644 34008 7648
rect 33944 7588 33948 7644
rect 33948 7588 34004 7644
rect 34004 7588 34008 7644
rect 33944 7584 34008 7588
rect 5046 7100 5110 7104
rect 5046 7044 5050 7100
rect 5050 7044 5106 7100
rect 5106 7044 5110 7100
rect 5046 7040 5110 7044
rect 5126 7100 5190 7104
rect 5126 7044 5130 7100
rect 5130 7044 5186 7100
rect 5186 7044 5190 7100
rect 5126 7040 5190 7044
rect 5206 7100 5270 7104
rect 5206 7044 5210 7100
rect 5210 7044 5266 7100
rect 5266 7044 5270 7100
rect 5206 7040 5270 7044
rect 5286 7100 5350 7104
rect 5286 7044 5290 7100
rect 5290 7044 5346 7100
rect 5346 7044 5350 7100
rect 5286 7040 5350 7044
rect 13234 7100 13298 7104
rect 13234 7044 13238 7100
rect 13238 7044 13294 7100
rect 13294 7044 13298 7100
rect 13234 7040 13298 7044
rect 13314 7100 13378 7104
rect 13314 7044 13318 7100
rect 13318 7044 13374 7100
rect 13374 7044 13378 7100
rect 13314 7040 13378 7044
rect 13394 7100 13458 7104
rect 13394 7044 13398 7100
rect 13398 7044 13454 7100
rect 13454 7044 13458 7100
rect 13394 7040 13458 7044
rect 13474 7100 13538 7104
rect 13474 7044 13478 7100
rect 13478 7044 13534 7100
rect 13534 7044 13538 7100
rect 13474 7040 13538 7044
rect 21422 7100 21486 7104
rect 21422 7044 21426 7100
rect 21426 7044 21482 7100
rect 21482 7044 21486 7100
rect 21422 7040 21486 7044
rect 21502 7100 21566 7104
rect 21502 7044 21506 7100
rect 21506 7044 21562 7100
rect 21562 7044 21566 7100
rect 21502 7040 21566 7044
rect 21582 7100 21646 7104
rect 21582 7044 21586 7100
rect 21586 7044 21642 7100
rect 21642 7044 21646 7100
rect 21582 7040 21646 7044
rect 21662 7100 21726 7104
rect 21662 7044 21666 7100
rect 21666 7044 21722 7100
rect 21722 7044 21726 7100
rect 21662 7040 21726 7044
rect 29610 7100 29674 7104
rect 29610 7044 29614 7100
rect 29614 7044 29670 7100
rect 29670 7044 29674 7100
rect 29610 7040 29674 7044
rect 29690 7100 29754 7104
rect 29690 7044 29694 7100
rect 29694 7044 29750 7100
rect 29750 7044 29754 7100
rect 29690 7040 29754 7044
rect 29770 7100 29834 7104
rect 29770 7044 29774 7100
rect 29774 7044 29830 7100
rect 29830 7044 29834 7100
rect 29770 7040 29834 7044
rect 29850 7100 29914 7104
rect 29850 7044 29854 7100
rect 29854 7044 29910 7100
rect 29910 7044 29914 7100
rect 29850 7040 29914 7044
rect 9140 6556 9204 6560
rect 9140 6500 9144 6556
rect 9144 6500 9200 6556
rect 9200 6500 9204 6556
rect 9140 6496 9204 6500
rect 9220 6556 9284 6560
rect 9220 6500 9224 6556
rect 9224 6500 9280 6556
rect 9280 6500 9284 6556
rect 9220 6496 9284 6500
rect 9300 6556 9364 6560
rect 9300 6500 9304 6556
rect 9304 6500 9360 6556
rect 9360 6500 9364 6556
rect 9300 6496 9364 6500
rect 9380 6556 9444 6560
rect 9380 6500 9384 6556
rect 9384 6500 9440 6556
rect 9440 6500 9444 6556
rect 9380 6496 9444 6500
rect 17328 6556 17392 6560
rect 17328 6500 17332 6556
rect 17332 6500 17388 6556
rect 17388 6500 17392 6556
rect 17328 6496 17392 6500
rect 17408 6556 17472 6560
rect 17408 6500 17412 6556
rect 17412 6500 17468 6556
rect 17468 6500 17472 6556
rect 17408 6496 17472 6500
rect 17488 6556 17552 6560
rect 17488 6500 17492 6556
rect 17492 6500 17548 6556
rect 17548 6500 17552 6556
rect 17488 6496 17552 6500
rect 17568 6556 17632 6560
rect 17568 6500 17572 6556
rect 17572 6500 17628 6556
rect 17628 6500 17632 6556
rect 17568 6496 17632 6500
rect 25516 6556 25580 6560
rect 25516 6500 25520 6556
rect 25520 6500 25576 6556
rect 25576 6500 25580 6556
rect 25516 6496 25580 6500
rect 25596 6556 25660 6560
rect 25596 6500 25600 6556
rect 25600 6500 25656 6556
rect 25656 6500 25660 6556
rect 25596 6496 25660 6500
rect 25676 6556 25740 6560
rect 25676 6500 25680 6556
rect 25680 6500 25736 6556
rect 25736 6500 25740 6556
rect 25676 6496 25740 6500
rect 25756 6556 25820 6560
rect 25756 6500 25760 6556
rect 25760 6500 25816 6556
rect 25816 6500 25820 6556
rect 25756 6496 25820 6500
rect 33704 6556 33768 6560
rect 33704 6500 33708 6556
rect 33708 6500 33764 6556
rect 33764 6500 33768 6556
rect 33704 6496 33768 6500
rect 33784 6556 33848 6560
rect 33784 6500 33788 6556
rect 33788 6500 33844 6556
rect 33844 6500 33848 6556
rect 33784 6496 33848 6500
rect 33864 6556 33928 6560
rect 33864 6500 33868 6556
rect 33868 6500 33924 6556
rect 33924 6500 33928 6556
rect 33864 6496 33928 6500
rect 33944 6556 34008 6560
rect 33944 6500 33948 6556
rect 33948 6500 34004 6556
rect 34004 6500 34008 6556
rect 33944 6496 34008 6500
rect 5046 6012 5110 6016
rect 5046 5956 5050 6012
rect 5050 5956 5106 6012
rect 5106 5956 5110 6012
rect 5046 5952 5110 5956
rect 5126 6012 5190 6016
rect 5126 5956 5130 6012
rect 5130 5956 5186 6012
rect 5186 5956 5190 6012
rect 5126 5952 5190 5956
rect 5206 6012 5270 6016
rect 5206 5956 5210 6012
rect 5210 5956 5266 6012
rect 5266 5956 5270 6012
rect 5206 5952 5270 5956
rect 5286 6012 5350 6016
rect 5286 5956 5290 6012
rect 5290 5956 5346 6012
rect 5346 5956 5350 6012
rect 5286 5952 5350 5956
rect 13234 6012 13298 6016
rect 13234 5956 13238 6012
rect 13238 5956 13294 6012
rect 13294 5956 13298 6012
rect 13234 5952 13298 5956
rect 13314 6012 13378 6016
rect 13314 5956 13318 6012
rect 13318 5956 13374 6012
rect 13374 5956 13378 6012
rect 13314 5952 13378 5956
rect 13394 6012 13458 6016
rect 13394 5956 13398 6012
rect 13398 5956 13454 6012
rect 13454 5956 13458 6012
rect 13394 5952 13458 5956
rect 13474 6012 13538 6016
rect 13474 5956 13478 6012
rect 13478 5956 13534 6012
rect 13534 5956 13538 6012
rect 13474 5952 13538 5956
rect 21422 6012 21486 6016
rect 21422 5956 21426 6012
rect 21426 5956 21482 6012
rect 21482 5956 21486 6012
rect 21422 5952 21486 5956
rect 21502 6012 21566 6016
rect 21502 5956 21506 6012
rect 21506 5956 21562 6012
rect 21562 5956 21566 6012
rect 21502 5952 21566 5956
rect 21582 6012 21646 6016
rect 21582 5956 21586 6012
rect 21586 5956 21642 6012
rect 21642 5956 21646 6012
rect 21582 5952 21646 5956
rect 21662 6012 21726 6016
rect 21662 5956 21666 6012
rect 21666 5956 21722 6012
rect 21722 5956 21726 6012
rect 21662 5952 21726 5956
rect 29610 6012 29674 6016
rect 29610 5956 29614 6012
rect 29614 5956 29670 6012
rect 29670 5956 29674 6012
rect 29610 5952 29674 5956
rect 29690 6012 29754 6016
rect 29690 5956 29694 6012
rect 29694 5956 29750 6012
rect 29750 5956 29754 6012
rect 29690 5952 29754 5956
rect 29770 6012 29834 6016
rect 29770 5956 29774 6012
rect 29774 5956 29830 6012
rect 29830 5956 29834 6012
rect 29770 5952 29834 5956
rect 29850 6012 29914 6016
rect 29850 5956 29854 6012
rect 29854 5956 29910 6012
rect 29910 5956 29914 6012
rect 29850 5952 29914 5956
rect 9140 5468 9204 5472
rect 9140 5412 9144 5468
rect 9144 5412 9200 5468
rect 9200 5412 9204 5468
rect 9140 5408 9204 5412
rect 9220 5468 9284 5472
rect 9220 5412 9224 5468
rect 9224 5412 9280 5468
rect 9280 5412 9284 5468
rect 9220 5408 9284 5412
rect 9300 5468 9364 5472
rect 9300 5412 9304 5468
rect 9304 5412 9360 5468
rect 9360 5412 9364 5468
rect 9300 5408 9364 5412
rect 9380 5468 9444 5472
rect 9380 5412 9384 5468
rect 9384 5412 9440 5468
rect 9440 5412 9444 5468
rect 9380 5408 9444 5412
rect 17328 5468 17392 5472
rect 17328 5412 17332 5468
rect 17332 5412 17388 5468
rect 17388 5412 17392 5468
rect 17328 5408 17392 5412
rect 17408 5468 17472 5472
rect 17408 5412 17412 5468
rect 17412 5412 17468 5468
rect 17468 5412 17472 5468
rect 17408 5408 17472 5412
rect 17488 5468 17552 5472
rect 17488 5412 17492 5468
rect 17492 5412 17548 5468
rect 17548 5412 17552 5468
rect 17488 5408 17552 5412
rect 17568 5468 17632 5472
rect 17568 5412 17572 5468
rect 17572 5412 17628 5468
rect 17628 5412 17632 5468
rect 17568 5408 17632 5412
rect 25516 5468 25580 5472
rect 25516 5412 25520 5468
rect 25520 5412 25576 5468
rect 25576 5412 25580 5468
rect 25516 5408 25580 5412
rect 25596 5468 25660 5472
rect 25596 5412 25600 5468
rect 25600 5412 25656 5468
rect 25656 5412 25660 5468
rect 25596 5408 25660 5412
rect 25676 5468 25740 5472
rect 25676 5412 25680 5468
rect 25680 5412 25736 5468
rect 25736 5412 25740 5468
rect 25676 5408 25740 5412
rect 25756 5468 25820 5472
rect 25756 5412 25760 5468
rect 25760 5412 25816 5468
rect 25816 5412 25820 5468
rect 25756 5408 25820 5412
rect 33704 5468 33768 5472
rect 33704 5412 33708 5468
rect 33708 5412 33764 5468
rect 33764 5412 33768 5468
rect 33704 5408 33768 5412
rect 33784 5468 33848 5472
rect 33784 5412 33788 5468
rect 33788 5412 33844 5468
rect 33844 5412 33848 5468
rect 33784 5408 33848 5412
rect 33864 5468 33928 5472
rect 33864 5412 33868 5468
rect 33868 5412 33924 5468
rect 33924 5412 33928 5468
rect 33864 5408 33928 5412
rect 33944 5468 34008 5472
rect 33944 5412 33948 5468
rect 33948 5412 34004 5468
rect 34004 5412 34008 5468
rect 33944 5408 34008 5412
rect 5046 4924 5110 4928
rect 5046 4868 5050 4924
rect 5050 4868 5106 4924
rect 5106 4868 5110 4924
rect 5046 4864 5110 4868
rect 5126 4924 5190 4928
rect 5126 4868 5130 4924
rect 5130 4868 5186 4924
rect 5186 4868 5190 4924
rect 5126 4864 5190 4868
rect 5206 4924 5270 4928
rect 5206 4868 5210 4924
rect 5210 4868 5266 4924
rect 5266 4868 5270 4924
rect 5206 4864 5270 4868
rect 5286 4924 5350 4928
rect 5286 4868 5290 4924
rect 5290 4868 5346 4924
rect 5346 4868 5350 4924
rect 5286 4864 5350 4868
rect 13234 4924 13298 4928
rect 13234 4868 13238 4924
rect 13238 4868 13294 4924
rect 13294 4868 13298 4924
rect 13234 4864 13298 4868
rect 13314 4924 13378 4928
rect 13314 4868 13318 4924
rect 13318 4868 13374 4924
rect 13374 4868 13378 4924
rect 13314 4864 13378 4868
rect 13394 4924 13458 4928
rect 13394 4868 13398 4924
rect 13398 4868 13454 4924
rect 13454 4868 13458 4924
rect 13394 4864 13458 4868
rect 13474 4924 13538 4928
rect 13474 4868 13478 4924
rect 13478 4868 13534 4924
rect 13534 4868 13538 4924
rect 13474 4864 13538 4868
rect 21422 4924 21486 4928
rect 21422 4868 21426 4924
rect 21426 4868 21482 4924
rect 21482 4868 21486 4924
rect 21422 4864 21486 4868
rect 21502 4924 21566 4928
rect 21502 4868 21506 4924
rect 21506 4868 21562 4924
rect 21562 4868 21566 4924
rect 21502 4864 21566 4868
rect 21582 4924 21646 4928
rect 21582 4868 21586 4924
rect 21586 4868 21642 4924
rect 21642 4868 21646 4924
rect 21582 4864 21646 4868
rect 21662 4924 21726 4928
rect 21662 4868 21666 4924
rect 21666 4868 21722 4924
rect 21722 4868 21726 4924
rect 21662 4864 21726 4868
rect 29610 4924 29674 4928
rect 29610 4868 29614 4924
rect 29614 4868 29670 4924
rect 29670 4868 29674 4924
rect 29610 4864 29674 4868
rect 29690 4924 29754 4928
rect 29690 4868 29694 4924
rect 29694 4868 29750 4924
rect 29750 4868 29754 4924
rect 29690 4864 29754 4868
rect 29770 4924 29834 4928
rect 29770 4868 29774 4924
rect 29774 4868 29830 4924
rect 29830 4868 29834 4924
rect 29770 4864 29834 4868
rect 29850 4924 29914 4928
rect 29850 4868 29854 4924
rect 29854 4868 29910 4924
rect 29910 4868 29914 4924
rect 29850 4864 29914 4868
rect 9140 4380 9204 4384
rect 9140 4324 9144 4380
rect 9144 4324 9200 4380
rect 9200 4324 9204 4380
rect 9140 4320 9204 4324
rect 9220 4380 9284 4384
rect 9220 4324 9224 4380
rect 9224 4324 9280 4380
rect 9280 4324 9284 4380
rect 9220 4320 9284 4324
rect 9300 4380 9364 4384
rect 9300 4324 9304 4380
rect 9304 4324 9360 4380
rect 9360 4324 9364 4380
rect 9300 4320 9364 4324
rect 9380 4380 9444 4384
rect 9380 4324 9384 4380
rect 9384 4324 9440 4380
rect 9440 4324 9444 4380
rect 9380 4320 9444 4324
rect 17328 4380 17392 4384
rect 17328 4324 17332 4380
rect 17332 4324 17388 4380
rect 17388 4324 17392 4380
rect 17328 4320 17392 4324
rect 17408 4380 17472 4384
rect 17408 4324 17412 4380
rect 17412 4324 17468 4380
rect 17468 4324 17472 4380
rect 17408 4320 17472 4324
rect 17488 4380 17552 4384
rect 17488 4324 17492 4380
rect 17492 4324 17548 4380
rect 17548 4324 17552 4380
rect 17488 4320 17552 4324
rect 17568 4380 17632 4384
rect 17568 4324 17572 4380
rect 17572 4324 17628 4380
rect 17628 4324 17632 4380
rect 17568 4320 17632 4324
rect 25516 4380 25580 4384
rect 25516 4324 25520 4380
rect 25520 4324 25576 4380
rect 25576 4324 25580 4380
rect 25516 4320 25580 4324
rect 25596 4380 25660 4384
rect 25596 4324 25600 4380
rect 25600 4324 25656 4380
rect 25656 4324 25660 4380
rect 25596 4320 25660 4324
rect 25676 4380 25740 4384
rect 25676 4324 25680 4380
rect 25680 4324 25736 4380
rect 25736 4324 25740 4380
rect 25676 4320 25740 4324
rect 25756 4380 25820 4384
rect 25756 4324 25760 4380
rect 25760 4324 25816 4380
rect 25816 4324 25820 4380
rect 25756 4320 25820 4324
rect 33704 4380 33768 4384
rect 33704 4324 33708 4380
rect 33708 4324 33764 4380
rect 33764 4324 33768 4380
rect 33704 4320 33768 4324
rect 33784 4380 33848 4384
rect 33784 4324 33788 4380
rect 33788 4324 33844 4380
rect 33844 4324 33848 4380
rect 33784 4320 33848 4324
rect 33864 4380 33928 4384
rect 33864 4324 33868 4380
rect 33868 4324 33924 4380
rect 33924 4324 33928 4380
rect 33864 4320 33928 4324
rect 33944 4380 34008 4384
rect 33944 4324 33948 4380
rect 33948 4324 34004 4380
rect 34004 4324 34008 4380
rect 33944 4320 34008 4324
rect 5046 3836 5110 3840
rect 5046 3780 5050 3836
rect 5050 3780 5106 3836
rect 5106 3780 5110 3836
rect 5046 3776 5110 3780
rect 5126 3836 5190 3840
rect 5126 3780 5130 3836
rect 5130 3780 5186 3836
rect 5186 3780 5190 3836
rect 5126 3776 5190 3780
rect 5206 3836 5270 3840
rect 5206 3780 5210 3836
rect 5210 3780 5266 3836
rect 5266 3780 5270 3836
rect 5206 3776 5270 3780
rect 5286 3836 5350 3840
rect 5286 3780 5290 3836
rect 5290 3780 5346 3836
rect 5346 3780 5350 3836
rect 5286 3776 5350 3780
rect 13234 3836 13298 3840
rect 13234 3780 13238 3836
rect 13238 3780 13294 3836
rect 13294 3780 13298 3836
rect 13234 3776 13298 3780
rect 13314 3836 13378 3840
rect 13314 3780 13318 3836
rect 13318 3780 13374 3836
rect 13374 3780 13378 3836
rect 13314 3776 13378 3780
rect 13394 3836 13458 3840
rect 13394 3780 13398 3836
rect 13398 3780 13454 3836
rect 13454 3780 13458 3836
rect 13394 3776 13458 3780
rect 13474 3836 13538 3840
rect 13474 3780 13478 3836
rect 13478 3780 13534 3836
rect 13534 3780 13538 3836
rect 13474 3776 13538 3780
rect 21422 3836 21486 3840
rect 21422 3780 21426 3836
rect 21426 3780 21482 3836
rect 21482 3780 21486 3836
rect 21422 3776 21486 3780
rect 21502 3836 21566 3840
rect 21502 3780 21506 3836
rect 21506 3780 21562 3836
rect 21562 3780 21566 3836
rect 21502 3776 21566 3780
rect 21582 3836 21646 3840
rect 21582 3780 21586 3836
rect 21586 3780 21642 3836
rect 21642 3780 21646 3836
rect 21582 3776 21646 3780
rect 21662 3836 21726 3840
rect 21662 3780 21666 3836
rect 21666 3780 21722 3836
rect 21722 3780 21726 3836
rect 21662 3776 21726 3780
rect 29610 3836 29674 3840
rect 29610 3780 29614 3836
rect 29614 3780 29670 3836
rect 29670 3780 29674 3836
rect 29610 3776 29674 3780
rect 29690 3836 29754 3840
rect 29690 3780 29694 3836
rect 29694 3780 29750 3836
rect 29750 3780 29754 3836
rect 29690 3776 29754 3780
rect 29770 3836 29834 3840
rect 29770 3780 29774 3836
rect 29774 3780 29830 3836
rect 29830 3780 29834 3836
rect 29770 3776 29834 3780
rect 29850 3836 29914 3840
rect 29850 3780 29854 3836
rect 29854 3780 29910 3836
rect 29910 3780 29914 3836
rect 29850 3776 29914 3780
rect 9140 3292 9204 3296
rect 9140 3236 9144 3292
rect 9144 3236 9200 3292
rect 9200 3236 9204 3292
rect 9140 3232 9204 3236
rect 9220 3292 9284 3296
rect 9220 3236 9224 3292
rect 9224 3236 9280 3292
rect 9280 3236 9284 3292
rect 9220 3232 9284 3236
rect 9300 3292 9364 3296
rect 9300 3236 9304 3292
rect 9304 3236 9360 3292
rect 9360 3236 9364 3292
rect 9300 3232 9364 3236
rect 9380 3292 9444 3296
rect 9380 3236 9384 3292
rect 9384 3236 9440 3292
rect 9440 3236 9444 3292
rect 9380 3232 9444 3236
rect 17328 3292 17392 3296
rect 17328 3236 17332 3292
rect 17332 3236 17388 3292
rect 17388 3236 17392 3292
rect 17328 3232 17392 3236
rect 17408 3292 17472 3296
rect 17408 3236 17412 3292
rect 17412 3236 17468 3292
rect 17468 3236 17472 3292
rect 17408 3232 17472 3236
rect 17488 3292 17552 3296
rect 17488 3236 17492 3292
rect 17492 3236 17548 3292
rect 17548 3236 17552 3292
rect 17488 3232 17552 3236
rect 17568 3292 17632 3296
rect 17568 3236 17572 3292
rect 17572 3236 17628 3292
rect 17628 3236 17632 3292
rect 17568 3232 17632 3236
rect 25516 3292 25580 3296
rect 25516 3236 25520 3292
rect 25520 3236 25576 3292
rect 25576 3236 25580 3292
rect 25516 3232 25580 3236
rect 25596 3292 25660 3296
rect 25596 3236 25600 3292
rect 25600 3236 25656 3292
rect 25656 3236 25660 3292
rect 25596 3232 25660 3236
rect 25676 3292 25740 3296
rect 25676 3236 25680 3292
rect 25680 3236 25736 3292
rect 25736 3236 25740 3292
rect 25676 3232 25740 3236
rect 25756 3292 25820 3296
rect 25756 3236 25760 3292
rect 25760 3236 25816 3292
rect 25816 3236 25820 3292
rect 25756 3232 25820 3236
rect 33704 3292 33768 3296
rect 33704 3236 33708 3292
rect 33708 3236 33764 3292
rect 33764 3236 33768 3292
rect 33704 3232 33768 3236
rect 33784 3292 33848 3296
rect 33784 3236 33788 3292
rect 33788 3236 33844 3292
rect 33844 3236 33848 3292
rect 33784 3232 33848 3236
rect 33864 3292 33928 3296
rect 33864 3236 33868 3292
rect 33868 3236 33924 3292
rect 33924 3236 33928 3292
rect 33864 3232 33928 3236
rect 33944 3292 34008 3296
rect 33944 3236 33948 3292
rect 33948 3236 34004 3292
rect 34004 3236 34008 3292
rect 33944 3232 34008 3236
rect 5046 2748 5110 2752
rect 5046 2692 5050 2748
rect 5050 2692 5106 2748
rect 5106 2692 5110 2748
rect 5046 2688 5110 2692
rect 5126 2748 5190 2752
rect 5126 2692 5130 2748
rect 5130 2692 5186 2748
rect 5186 2692 5190 2748
rect 5126 2688 5190 2692
rect 5206 2748 5270 2752
rect 5206 2692 5210 2748
rect 5210 2692 5266 2748
rect 5266 2692 5270 2748
rect 5206 2688 5270 2692
rect 5286 2748 5350 2752
rect 5286 2692 5290 2748
rect 5290 2692 5346 2748
rect 5346 2692 5350 2748
rect 5286 2688 5350 2692
rect 13234 2748 13298 2752
rect 13234 2692 13238 2748
rect 13238 2692 13294 2748
rect 13294 2692 13298 2748
rect 13234 2688 13298 2692
rect 13314 2748 13378 2752
rect 13314 2692 13318 2748
rect 13318 2692 13374 2748
rect 13374 2692 13378 2748
rect 13314 2688 13378 2692
rect 13394 2748 13458 2752
rect 13394 2692 13398 2748
rect 13398 2692 13454 2748
rect 13454 2692 13458 2748
rect 13394 2688 13458 2692
rect 13474 2748 13538 2752
rect 13474 2692 13478 2748
rect 13478 2692 13534 2748
rect 13534 2692 13538 2748
rect 13474 2688 13538 2692
rect 21422 2748 21486 2752
rect 21422 2692 21426 2748
rect 21426 2692 21482 2748
rect 21482 2692 21486 2748
rect 21422 2688 21486 2692
rect 21502 2748 21566 2752
rect 21502 2692 21506 2748
rect 21506 2692 21562 2748
rect 21562 2692 21566 2748
rect 21502 2688 21566 2692
rect 21582 2748 21646 2752
rect 21582 2692 21586 2748
rect 21586 2692 21642 2748
rect 21642 2692 21646 2748
rect 21582 2688 21646 2692
rect 21662 2748 21726 2752
rect 21662 2692 21666 2748
rect 21666 2692 21722 2748
rect 21722 2692 21726 2748
rect 21662 2688 21726 2692
rect 29610 2748 29674 2752
rect 29610 2692 29614 2748
rect 29614 2692 29670 2748
rect 29670 2692 29674 2748
rect 29610 2688 29674 2692
rect 29690 2748 29754 2752
rect 29690 2692 29694 2748
rect 29694 2692 29750 2748
rect 29750 2692 29754 2748
rect 29690 2688 29754 2692
rect 29770 2748 29834 2752
rect 29770 2692 29774 2748
rect 29774 2692 29830 2748
rect 29830 2692 29834 2748
rect 29770 2688 29834 2692
rect 29850 2748 29914 2752
rect 29850 2692 29854 2748
rect 29854 2692 29910 2748
rect 29910 2692 29914 2748
rect 29850 2688 29914 2692
rect 9140 2204 9204 2208
rect 9140 2148 9144 2204
rect 9144 2148 9200 2204
rect 9200 2148 9204 2204
rect 9140 2144 9204 2148
rect 9220 2204 9284 2208
rect 9220 2148 9224 2204
rect 9224 2148 9280 2204
rect 9280 2148 9284 2204
rect 9220 2144 9284 2148
rect 9300 2204 9364 2208
rect 9300 2148 9304 2204
rect 9304 2148 9360 2204
rect 9360 2148 9364 2204
rect 9300 2144 9364 2148
rect 9380 2204 9444 2208
rect 9380 2148 9384 2204
rect 9384 2148 9440 2204
rect 9440 2148 9444 2204
rect 9380 2144 9444 2148
rect 17328 2204 17392 2208
rect 17328 2148 17332 2204
rect 17332 2148 17388 2204
rect 17388 2148 17392 2204
rect 17328 2144 17392 2148
rect 17408 2204 17472 2208
rect 17408 2148 17412 2204
rect 17412 2148 17468 2204
rect 17468 2148 17472 2204
rect 17408 2144 17472 2148
rect 17488 2204 17552 2208
rect 17488 2148 17492 2204
rect 17492 2148 17548 2204
rect 17548 2148 17552 2204
rect 17488 2144 17552 2148
rect 17568 2204 17632 2208
rect 17568 2148 17572 2204
rect 17572 2148 17628 2204
rect 17628 2148 17632 2204
rect 17568 2144 17632 2148
rect 25516 2204 25580 2208
rect 25516 2148 25520 2204
rect 25520 2148 25576 2204
rect 25576 2148 25580 2204
rect 25516 2144 25580 2148
rect 25596 2204 25660 2208
rect 25596 2148 25600 2204
rect 25600 2148 25656 2204
rect 25656 2148 25660 2204
rect 25596 2144 25660 2148
rect 25676 2204 25740 2208
rect 25676 2148 25680 2204
rect 25680 2148 25736 2204
rect 25736 2148 25740 2204
rect 25676 2144 25740 2148
rect 25756 2204 25820 2208
rect 25756 2148 25760 2204
rect 25760 2148 25816 2204
rect 25816 2148 25820 2204
rect 25756 2144 25820 2148
rect 33704 2204 33768 2208
rect 33704 2148 33708 2204
rect 33708 2148 33764 2204
rect 33764 2148 33768 2204
rect 33704 2144 33768 2148
rect 33784 2204 33848 2208
rect 33784 2148 33788 2204
rect 33788 2148 33844 2204
rect 33844 2148 33848 2204
rect 33784 2144 33848 2148
rect 33864 2204 33928 2208
rect 33864 2148 33868 2204
rect 33868 2148 33924 2204
rect 33924 2148 33928 2204
rect 33864 2144 33928 2148
rect 33944 2204 34008 2208
rect 33944 2148 33948 2204
rect 33948 2148 34004 2204
rect 34004 2148 34008 2204
rect 33944 2144 34008 2148
<< metal4 >>
rect 5038 32128 5358 32688
rect 5038 32064 5046 32128
rect 5110 32064 5126 32128
rect 5190 32064 5206 32128
rect 5270 32064 5286 32128
rect 5350 32064 5358 32128
rect 5038 31040 5358 32064
rect 5038 30976 5046 31040
rect 5110 30976 5126 31040
rect 5190 30976 5206 31040
rect 5270 30976 5286 31040
rect 5350 30976 5358 31040
rect 5038 29952 5358 30976
rect 5038 29888 5046 29952
rect 5110 29888 5126 29952
rect 5190 29888 5206 29952
rect 5270 29888 5286 29952
rect 5350 29888 5358 29952
rect 5038 28864 5358 29888
rect 5038 28800 5046 28864
rect 5110 28800 5126 28864
rect 5190 28800 5206 28864
rect 5270 28800 5286 28864
rect 5350 28800 5358 28864
rect 5038 27776 5358 28800
rect 5038 27712 5046 27776
rect 5110 27712 5126 27776
rect 5190 27712 5206 27776
rect 5270 27712 5286 27776
rect 5350 27712 5358 27776
rect 5038 26688 5358 27712
rect 5038 26624 5046 26688
rect 5110 26624 5126 26688
rect 5190 26624 5206 26688
rect 5270 26624 5286 26688
rect 5350 26624 5358 26688
rect 5038 25600 5358 26624
rect 5038 25536 5046 25600
rect 5110 25536 5126 25600
rect 5190 25536 5206 25600
rect 5270 25536 5286 25600
rect 5350 25536 5358 25600
rect 5038 24512 5358 25536
rect 5038 24448 5046 24512
rect 5110 24448 5126 24512
rect 5190 24448 5206 24512
rect 5270 24448 5286 24512
rect 5350 24448 5358 24512
rect 5038 23424 5358 24448
rect 5038 23360 5046 23424
rect 5110 23360 5126 23424
rect 5190 23360 5206 23424
rect 5270 23360 5286 23424
rect 5350 23360 5358 23424
rect 5038 22336 5358 23360
rect 5038 22272 5046 22336
rect 5110 22272 5126 22336
rect 5190 22272 5206 22336
rect 5270 22272 5286 22336
rect 5350 22272 5358 22336
rect 5038 21248 5358 22272
rect 5038 21184 5046 21248
rect 5110 21184 5126 21248
rect 5190 21184 5206 21248
rect 5270 21184 5286 21248
rect 5350 21184 5358 21248
rect 5038 20160 5358 21184
rect 5038 20096 5046 20160
rect 5110 20096 5126 20160
rect 5190 20096 5206 20160
rect 5270 20096 5286 20160
rect 5350 20096 5358 20160
rect 5038 19072 5358 20096
rect 5038 19008 5046 19072
rect 5110 19008 5126 19072
rect 5190 19008 5206 19072
rect 5270 19008 5286 19072
rect 5350 19008 5358 19072
rect 5038 17984 5358 19008
rect 5038 17920 5046 17984
rect 5110 17920 5126 17984
rect 5190 17920 5206 17984
rect 5270 17920 5286 17984
rect 5350 17920 5358 17984
rect 5038 16896 5358 17920
rect 5038 16832 5046 16896
rect 5110 16832 5126 16896
rect 5190 16832 5206 16896
rect 5270 16832 5286 16896
rect 5350 16832 5358 16896
rect 5038 15808 5358 16832
rect 5038 15744 5046 15808
rect 5110 15744 5126 15808
rect 5190 15744 5206 15808
rect 5270 15744 5286 15808
rect 5350 15744 5358 15808
rect 5038 14720 5358 15744
rect 5038 14656 5046 14720
rect 5110 14656 5126 14720
rect 5190 14656 5206 14720
rect 5270 14656 5286 14720
rect 5350 14656 5358 14720
rect 5038 13632 5358 14656
rect 5038 13568 5046 13632
rect 5110 13568 5126 13632
rect 5190 13568 5206 13632
rect 5270 13568 5286 13632
rect 5350 13568 5358 13632
rect 5038 12544 5358 13568
rect 5038 12480 5046 12544
rect 5110 12480 5126 12544
rect 5190 12480 5206 12544
rect 5270 12480 5286 12544
rect 5350 12480 5358 12544
rect 5038 11456 5358 12480
rect 5038 11392 5046 11456
rect 5110 11392 5126 11456
rect 5190 11392 5206 11456
rect 5270 11392 5286 11456
rect 5350 11392 5358 11456
rect 5038 10368 5358 11392
rect 5038 10304 5046 10368
rect 5110 10304 5126 10368
rect 5190 10304 5206 10368
rect 5270 10304 5286 10368
rect 5350 10304 5358 10368
rect 5038 9280 5358 10304
rect 5038 9216 5046 9280
rect 5110 9216 5126 9280
rect 5190 9216 5206 9280
rect 5270 9216 5286 9280
rect 5350 9216 5358 9280
rect 5038 8192 5358 9216
rect 5038 8128 5046 8192
rect 5110 8128 5126 8192
rect 5190 8128 5206 8192
rect 5270 8128 5286 8192
rect 5350 8128 5358 8192
rect 5038 7104 5358 8128
rect 5038 7040 5046 7104
rect 5110 7040 5126 7104
rect 5190 7040 5206 7104
rect 5270 7040 5286 7104
rect 5350 7040 5358 7104
rect 5038 6016 5358 7040
rect 5038 5952 5046 6016
rect 5110 5952 5126 6016
rect 5190 5952 5206 6016
rect 5270 5952 5286 6016
rect 5350 5952 5358 6016
rect 5038 4928 5358 5952
rect 5038 4864 5046 4928
rect 5110 4864 5126 4928
rect 5190 4864 5206 4928
rect 5270 4864 5286 4928
rect 5350 4864 5358 4928
rect 5038 3840 5358 4864
rect 5038 3776 5046 3840
rect 5110 3776 5126 3840
rect 5190 3776 5206 3840
rect 5270 3776 5286 3840
rect 5350 3776 5358 3840
rect 5038 2752 5358 3776
rect 5038 2688 5046 2752
rect 5110 2688 5126 2752
rect 5190 2688 5206 2752
rect 5270 2688 5286 2752
rect 5350 2688 5358 2752
rect 5038 2128 5358 2688
rect 9132 32672 9452 32688
rect 9132 32608 9140 32672
rect 9204 32608 9220 32672
rect 9284 32608 9300 32672
rect 9364 32608 9380 32672
rect 9444 32608 9452 32672
rect 9132 31584 9452 32608
rect 9132 31520 9140 31584
rect 9204 31520 9220 31584
rect 9284 31520 9300 31584
rect 9364 31520 9380 31584
rect 9444 31520 9452 31584
rect 9132 30496 9452 31520
rect 9132 30432 9140 30496
rect 9204 30432 9220 30496
rect 9284 30432 9300 30496
rect 9364 30432 9380 30496
rect 9444 30432 9452 30496
rect 9132 29408 9452 30432
rect 9132 29344 9140 29408
rect 9204 29344 9220 29408
rect 9284 29344 9300 29408
rect 9364 29344 9380 29408
rect 9444 29344 9452 29408
rect 9132 28320 9452 29344
rect 9132 28256 9140 28320
rect 9204 28256 9220 28320
rect 9284 28256 9300 28320
rect 9364 28256 9380 28320
rect 9444 28256 9452 28320
rect 9132 27232 9452 28256
rect 9132 27168 9140 27232
rect 9204 27168 9220 27232
rect 9284 27168 9300 27232
rect 9364 27168 9380 27232
rect 9444 27168 9452 27232
rect 9132 26144 9452 27168
rect 9132 26080 9140 26144
rect 9204 26080 9220 26144
rect 9284 26080 9300 26144
rect 9364 26080 9380 26144
rect 9444 26080 9452 26144
rect 9132 25056 9452 26080
rect 9132 24992 9140 25056
rect 9204 24992 9220 25056
rect 9284 24992 9300 25056
rect 9364 24992 9380 25056
rect 9444 24992 9452 25056
rect 9132 23968 9452 24992
rect 9132 23904 9140 23968
rect 9204 23904 9220 23968
rect 9284 23904 9300 23968
rect 9364 23904 9380 23968
rect 9444 23904 9452 23968
rect 9132 22880 9452 23904
rect 9132 22816 9140 22880
rect 9204 22816 9220 22880
rect 9284 22816 9300 22880
rect 9364 22816 9380 22880
rect 9444 22816 9452 22880
rect 9132 21792 9452 22816
rect 9132 21728 9140 21792
rect 9204 21728 9220 21792
rect 9284 21728 9300 21792
rect 9364 21728 9380 21792
rect 9444 21728 9452 21792
rect 9132 20704 9452 21728
rect 9132 20640 9140 20704
rect 9204 20640 9220 20704
rect 9284 20640 9300 20704
rect 9364 20640 9380 20704
rect 9444 20640 9452 20704
rect 9132 19616 9452 20640
rect 9132 19552 9140 19616
rect 9204 19552 9220 19616
rect 9284 19552 9300 19616
rect 9364 19552 9380 19616
rect 9444 19552 9452 19616
rect 9132 18528 9452 19552
rect 9132 18464 9140 18528
rect 9204 18464 9220 18528
rect 9284 18464 9300 18528
rect 9364 18464 9380 18528
rect 9444 18464 9452 18528
rect 9132 17440 9452 18464
rect 9132 17376 9140 17440
rect 9204 17376 9220 17440
rect 9284 17376 9300 17440
rect 9364 17376 9380 17440
rect 9444 17376 9452 17440
rect 9132 16352 9452 17376
rect 9132 16288 9140 16352
rect 9204 16288 9220 16352
rect 9284 16288 9300 16352
rect 9364 16288 9380 16352
rect 9444 16288 9452 16352
rect 9132 15264 9452 16288
rect 9132 15200 9140 15264
rect 9204 15200 9220 15264
rect 9284 15200 9300 15264
rect 9364 15200 9380 15264
rect 9444 15200 9452 15264
rect 9132 14176 9452 15200
rect 9132 14112 9140 14176
rect 9204 14112 9220 14176
rect 9284 14112 9300 14176
rect 9364 14112 9380 14176
rect 9444 14112 9452 14176
rect 9132 13088 9452 14112
rect 9132 13024 9140 13088
rect 9204 13024 9220 13088
rect 9284 13024 9300 13088
rect 9364 13024 9380 13088
rect 9444 13024 9452 13088
rect 9132 12000 9452 13024
rect 9132 11936 9140 12000
rect 9204 11936 9220 12000
rect 9284 11936 9300 12000
rect 9364 11936 9380 12000
rect 9444 11936 9452 12000
rect 9132 10912 9452 11936
rect 9132 10848 9140 10912
rect 9204 10848 9220 10912
rect 9284 10848 9300 10912
rect 9364 10848 9380 10912
rect 9444 10848 9452 10912
rect 9132 9824 9452 10848
rect 9132 9760 9140 9824
rect 9204 9760 9220 9824
rect 9284 9760 9300 9824
rect 9364 9760 9380 9824
rect 9444 9760 9452 9824
rect 9132 8736 9452 9760
rect 9132 8672 9140 8736
rect 9204 8672 9220 8736
rect 9284 8672 9300 8736
rect 9364 8672 9380 8736
rect 9444 8672 9452 8736
rect 9132 7648 9452 8672
rect 9132 7584 9140 7648
rect 9204 7584 9220 7648
rect 9284 7584 9300 7648
rect 9364 7584 9380 7648
rect 9444 7584 9452 7648
rect 9132 6560 9452 7584
rect 9132 6496 9140 6560
rect 9204 6496 9220 6560
rect 9284 6496 9300 6560
rect 9364 6496 9380 6560
rect 9444 6496 9452 6560
rect 9132 5472 9452 6496
rect 9132 5408 9140 5472
rect 9204 5408 9220 5472
rect 9284 5408 9300 5472
rect 9364 5408 9380 5472
rect 9444 5408 9452 5472
rect 9132 4384 9452 5408
rect 9132 4320 9140 4384
rect 9204 4320 9220 4384
rect 9284 4320 9300 4384
rect 9364 4320 9380 4384
rect 9444 4320 9452 4384
rect 9132 3296 9452 4320
rect 9132 3232 9140 3296
rect 9204 3232 9220 3296
rect 9284 3232 9300 3296
rect 9364 3232 9380 3296
rect 9444 3232 9452 3296
rect 9132 2208 9452 3232
rect 9132 2144 9140 2208
rect 9204 2144 9220 2208
rect 9284 2144 9300 2208
rect 9364 2144 9380 2208
rect 9444 2144 9452 2208
rect 9132 2128 9452 2144
rect 13226 32128 13546 32688
rect 13226 32064 13234 32128
rect 13298 32064 13314 32128
rect 13378 32064 13394 32128
rect 13458 32064 13474 32128
rect 13538 32064 13546 32128
rect 13226 31040 13546 32064
rect 13226 30976 13234 31040
rect 13298 30976 13314 31040
rect 13378 30976 13394 31040
rect 13458 30976 13474 31040
rect 13538 30976 13546 31040
rect 13226 29952 13546 30976
rect 13226 29888 13234 29952
rect 13298 29888 13314 29952
rect 13378 29888 13394 29952
rect 13458 29888 13474 29952
rect 13538 29888 13546 29952
rect 13226 28864 13546 29888
rect 13226 28800 13234 28864
rect 13298 28800 13314 28864
rect 13378 28800 13394 28864
rect 13458 28800 13474 28864
rect 13538 28800 13546 28864
rect 13226 27776 13546 28800
rect 13226 27712 13234 27776
rect 13298 27712 13314 27776
rect 13378 27712 13394 27776
rect 13458 27712 13474 27776
rect 13538 27712 13546 27776
rect 13226 26688 13546 27712
rect 13226 26624 13234 26688
rect 13298 26624 13314 26688
rect 13378 26624 13394 26688
rect 13458 26624 13474 26688
rect 13538 26624 13546 26688
rect 13226 25600 13546 26624
rect 13226 25536 13234 25600
rect 13298 25536 13314 25600
rect 13378 25536 13394 25600
rect 13458 25536 13474 25600
rect 13538 25536 13546 25600
rect 13226 24512 13546 25536
rect 13226 24448 13234 24512
rect 13298 24448 13314 24512
rect 13378 24448 13394 24512
rect 13458 24448 13474 24512
rect 13538 24448 13546 24512
rect 13226 23424 13546 24448
rect 13226 23360 13234 23424
rect 13298 23360 13314 23424
rect 13378 23360 13394 23424
rect 13458 23360 13474 23424
rect 13538 23360 13546 23424
rect 13226 22336 13546 23360
rect 13226 22272 13234 22336
rect 13298 22272 13314 22336
rect 13378 22272 13394 22336
rect 13458 22272 13474 22336
rect 13538 22272 13546 22336
rect 13226 21248 13546 22272
rect 13226 21184 13234 21248
rect 13298 21184 13314 21248
rect 13378 21184 13394 21248
rect 13458 21184 13474 21248
rect 13538 21184 13546 21248
rect 13226 20160 13546 21184
rect 13226 20096 13234 20160
rect 13298 20096 13314 20160
rect 13378 20096 13394 20160
rect 13458 20096 13474 20160
rect 13538 20096 13546 20160
rect 13226 19072 13546 20096
rect 13226 19008 13234 19072
rect 13298 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13546 19072
rect 13226 17984 13546 19008
rect 13226 17920 13234 17984
rect 13298 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13546 17984
rect 13226 16896 13546 17920
rect 13226 16832 13234 16896
rect 13298 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13546 16896
rect 13226 15808 13546 16832
rect 13226 15744 13234 15808
rect 13298 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13546 15808
rect 13226 14720 13546 15744
rect 13226 14656 13234 14720
rect 13298 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13546 14720
rect 13226 13632 13546 14656
rect 13226 13568 13234 13632
rect 13298 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13546 13632
rect 13226 12544 13546 13568
rect 13226 12480 13234 12544
rect 13298 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13546 12544
rect 13226 11456 13546 12480
rect 13226 11392 13234 11456
rect 13298 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13546 11456
rect 13226 10368 13546 11392
rect 13226 10304 13234 10368
rect 13298 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13546 10368
rect 13226 9280 13546 10304
rect 13226 9216 13234 9280
rect 13298 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13546 9280
rect 13226 8192 13546 9216
rect 13226 8128 13234 8192
rect 13298 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13546 8192
rect 13226 7104 13546 8128
rect 13226 7040 13234 7104
rect 13298 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13546 7104
rect 13226 6016 13546 7040
rect 13226 5952 13234 6016
rect 13298 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13546 6016
rect 13226 4928 13546 5952
rect 13226 4864 13234 4928
rect 13298 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13546 4928
rect 13226 3840 13546 4864
rect 13226 3776 13234 3840
rect 13298 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13546 3840
rect 13226 2752 13546 3776
rect 13226 2688 13234 2752
rect 13298 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13546 2752
rect 13226 2128 13546 2688
rect 17320 32672 17640 32688
rect 17320 32608 17328 32672
rect 17392 32608 17408 32672
rect 17472 32608 17488 32672
rect 17552 32608 17568 32672
rect 17632 32608 17640 32672
rect 17320 31584 17640 32608
rect 17320 31520 17328 31584
rect 17392 31520 17408 31584
rect 17472 31520 17488 31584
rect 17552 31520 17568 31584
rect 17632 31520 17640 31584
rect 17320 30496 17640 31520
rect 17320 30432 17328 30496
rect 17392 30432 17408 30496
rect 17472 30432 17488 30496
rect 17552 30432 17568 30496
rect 17632 30432 17640 30496
rect 17320 29408 17640 30432
rect 17320 29344 17328 29408
rect 17392 29344 17408 29408
rect 17472 29344 17488 29408
rect 17552 29344 17568 29408
rect 17632 29344 17640 29408
rect 17320 28320 17640 29344
rect 17320 28256 17328 28320
rect 17392 28256 17408 28320
rect 17472 28256 17488 28320
rect 17552 28256 17568 28320
rect 17632 28256 17640 28320
rect 17320 27232 17640 28256
rect 17320 27168 17328 27232
rect 17392 27168 17408 27232
rect 17472 27168 17488 27232
rect 17552 27168 17568 27232
rect 17632 27168 17640 27232
rect 17320 26144 17640 27168
rect 17320 26080 17328 26144
rect 17392 26080 17408 26144
rect 17472 26080 17488 26144
rect 17552 26080 17568 26144
rect 17632 26080 17640 26144
rect 17320 25056 17640 26080
rect 17320 24992 17328 25056
rect 17392 24992 17408 25056
rect 17472 24992 17488 25056
rect 17552 24992 17568 25056
rect 17632 24992 17640 25056
rect 17320 23968 17640 24992
rect 17320 23904 17328 23968
rect 17392 23904 17408 23968
rect 17472 23904 17488 23968
rect 17552 23904 17568 23968
rect 17632 23904 17640 23968
rect 17320 22880 17640 23904
rect 17320 22816 17328 22880
rect 17392 22816 17408 22880
rect 17472 22816 17488 22880
rect 17552 22816 17568 22880
rect 17632 22816 17640 22880
rect 17320 21792 17640 22816
rect 17320 21728 17328 21792
rect 17392 21728 17408 21792
rect 17472 21728 17488 21792
rect 17552 21728 17568 21792
rect 17632 21728 17640 21792
rect 17320 20704 17640 21728
rect 17320 20640 17328 20704
rect 17392 20640 17408 20704
rect 17472 20640 17488 20704
rect 17552 20640 17568 20704
rect 17632 20640 17640 20704
rect 17320 19616 17640 20640
rect 17320 19552 17328 19616
rect 17392 19552 17408 19616
rect 17472 19552 17488 19616
rect 17552 19552 17568 19616
rect 17632 19552 17640 19616
rect 17320 18528 17640 19552
rect 17320 18464 17328 18528
rect 17392 18464 17408 18528
rect 17472 18464 17488 18528
rect 17552 18464 17568 18528
rect 17632 18464 17640 18528
rect 17320 17440 17640 18464
rect 17320 17376 17328 17440
rect 17392 17376 17408 17440
rect 17472 17376 17488 17440
rect 17552 17376 17568 17440
rect 17632 17376 17640 17440
rect 17320 16352 17640 17376
rect 17320 16288 17328 16352
rect 17392 16288 17408 16352
rect 17472 16288 17488 16352
rect 17552 16288 17568 16352
rect 17632 16288 17640 16352
rect 17320 15264 17640 16288
rect 17320 15200 17328 15264
rect 17392 15200 17408 15264
rect 17472 15200 17488 15264
rect 17552 15200 17568 15264
rect 17632 15200 17640 15264
rect 17320 14176 17640 15200
rect 17320 14112 17328 14176
rect 17392 14112 17408 14176
rect 17472 14112 17488 14176
rect 17552 14112 17568 14176
rect 17632 14112 17640 14176
rect 17320 13088 17640 14112
rect 17320 13024 17328 13088
rect 17392 13024 17408 13088
rect 17472 13024 17488 13088
rect 17552 13024 17568 13088
rect 17632 13024 17640 13088
rect 17320 12000 17640 13024
rect 17320 11936 17328 12000
rect 17392 11936 17408 12000
rect 17472 11936 17488 12000
rect 17552 11936 17568 12000
rect 17632 11936 17640 12000
rect 17320 10912 17640 11936
rect 17320 10848 17328 10912
rect 17392 10848 17408 10912
rect 17472 10848 17488 10912
rect 17552 10848 17568 10912
rect 17632 10848 17640 10912
rect 17320 9824 17640 10848
rect 17320 9760 17328 9824
rect 17392 9760 17408 9824
rect 17472 9760 17488 9824
rect 17552 9760 17568 9824
rect 17632 9760 17640 9824
rect 17320 8736 17640 9760
rect 17320 8672 17328 8736
rect 17392 8672 17408 8736
rect 17472 8672 17488 8736
rect 17552 8672 17568 8736
rect 17632 8672 17640 8736
rect 17320 7648 17640 8672
rect 17320 7584 17328 7648
rect 17392 7584 17408 7648
rect 17472 7584 17488 7648
rect 17552 7584 17568 7648
rect 17632 7584 17640 7648
rect 17320 6560 17640 7584
rect 17320 6496 17328 6560
rect 17392 6496 17408 6560
rect 17472 6496 17488 6560
rect 17552 6496 17568 6560
rect 17632 6496 17640 6560
rect 17320 5472 17640 6496
rect 17320 5408 17328 5472
rect 17392 5408 17408 5472
rect 17472 5408 17488 5472
rect 17552 5408 17568 5472
rect 17632 5408 17640 5472
rect 17320 4384 17640 5408
rect 17320 4320 17328 4384
rect 17392 4320 17408 4384
rect 17472 4320 17488 4384
rect 17552 4320 17568 4384
rect 17632 4320 17640 4384
rect 17320 3296 17640 4320
rect 17320 3232 17328 3296
rect 17392 3232 17408 3296
rect 17472 3232 17488 3296
rect 17552 3232 17568 3296
rect 17632 3232 17640 3296
rect 17320 2208 17640 3232
rect 17320 2144 17328 2208
rect 17392 2144 17408 2208
rect 17472 2144 17488 2208
rect 17552 2144 17568 2208
rect 17632 2144 17640 2208
rect 17320 2128 17640 2144
rect 21414 32128 21734 32688
rect 21414 32064 21422 32128
rect 21486 32064 21502 32128
rect 21566 32064 21582 32128
rect 21646 32064 21662 32128
rect 21726 32064 21734 32128
rect 21414 31040 21734 32064
rect 21414 30976 21422 31040
rect 21486 30976 21502 31040
rect 21566 30976 21582 31040
rect 21646 30976 21662 31040
rect 21726 30976 21734 31040
rect 21414 29952 21734 30976
rect 21414 29888 21422 29952
rect 21486 29888 21502 29952
rect 21566 29888 21582 29952
rect 21646 29888 21662 29952
rect 21726 29888 21734 29952
rect 21414 28864 21734 29888
rect 21414 28800 21422 28864
rect 21486 28800 21502 28864
rect 21566 28800 21582 28864
rect 21646 28800 21662 28864
rect 21726 28800 21734 28864
rect 21414 27776 21734 28800
rect 21414 27712 21422 27776
rect 21486 27712 21502 27776
rect 21566 27712 21582 27776
rect 21646 27712 21662 27776
rect 21726 27712 21734 27776
rect 21414 26688 21734 27712
rect 21414 26624 21422 26688
rect 21486 26624 21502 26688
rect 21566 26624 21582 26688
rect 21646 26624 21662 26688
rect 21726 26624 21734 26688
rect 21414 25600 21734 26624
rect 21414 25536 21422 25600
rect 21486 25536 21502 25600
rect 21566 25536 21582 25600
rect 21646 25536 21662 25600
rect 21726 25536 21734 25600
rect 21414 24512 21734 25536
rect 21414 24448 21422 24512
rect 21486 24448 21502 24512
rect 21566 24448 21582 24512
rect 21646 24448 21662 24512
rect 21726 24448 21734 24512
rect 21414 23424 21734 24448
rect 21414 23360 21422 23424
rect 21486 23360 21502 23424
rect 21566 23360 21582 23424
rect 21646 23360 21662 23424
rect 21726 23360 21734 23424
rect 21414 22336 21734 23360
rect 21414 22272 21422 22336
rect 21486 22272 21502 22336
rect 21566 22272 21582 22336
rect 21646 22272 21662 22336
rect 21726 22272 21734 22336
rect 21414 21248 21734 22272
rect 21414 21184 21422 21248
rect 21486 21184 21502 21248
rect 21566 21184 21582 21248
rect 21646 21184 21662 21248
rect 21726 21184 21734 21248
rect 21414 20160 21734 21184
rect 21414 20096 21422 20160
rect 21486 20096 21502 20160
rect 21566 20096 21582 20160
rect 21646 20096 21662 20160
rect 21726 20096 21734 20160
rect 21414 19072 21734 20096
rect 21414 19008 21422 19072
rect 21486 19008 21502 19072
rect 21566 19008 21582 19072
rect 21646 19008 21662 19072
rect 21726 19008 21734 19072
rect 21414 17984 21734 19008
rect 21414 17920 21422 17984
rect 21486 17920 21502 17984
rect 21566 17920 21582 17984
rect 21646 17920 21662 17984
rect 21726 17920 21734 17984
rect 21414 16896 21734 17920
rect 21414 16832 21422 16896
rect 21486 16832 21502 16896
rect 21566 16832 21582 16896
rect 21646 16832 21662 16896
rect 21726 16832 21734 16896
rect 21414 15808 21734 16832
rect 21414 15744 21422 15808
rect 21486 15744 21502 15808
rect 21566 15744 21582 15808
rect 21646 15744 21662 15808
rect 21726 15744 21734 15808
rect 21414 14720 21734 15744
rect 21414 14656 21422 14720
rect 21486 14656 21502 14720
rect 21566 14656 21582 14720
rect 21646 14656 21662 14720
rect 21726 14656 21734 14720
rect 21414 13632 21734 14656
rect 21414 13568 21422 13632
rect 21486 13568 21502 13632
rect 21566 13568 21582 13632
rect 21646 13568 21662 13632
rect 21726 13568 21734 13632
rect 21414 12544 21734 13568
rect 21414 12480 21422 12544
rect 21486 12480 21502 12544
rect 21566 12480 21582 12544
rect 21646 12480 21662 12544
rect 21726 12480 21734 12544
rect 21414 11456 21734 12480
rect 21414 11392 21422 11456
rect 21486 11392 21502 11456
rect 21566 11392 21582 11456
rect 21646 11392 21662 11456
rect 21726 11392 21734 11456
rect 21414 10368 21734 11392
rect 21414 10304 21422 10368
rect 21486 10304 21502 10368
rect 21566 10304 21582 10368
rect 21646 10304 21662 10368
rect 21726 10304 21734 10368
rect 21414 9280 21734 10304
rect 21414 9216 21422 9280
rect 21486 9216 21502 9280
rect 21566 9216 21582 9280
rect 21646 9216 21662 9280
rect 21726 9216 21734 9280
rect 21414 8192 21734 9216
rect 21414 8128 21422 8192
rect 21486 8128 21502 8192
rect 21566 8128 21582 8192
rect 21646 8128 21662 8192
rect 21726 8128 21734 8192
rect 21414 7104 21734 8128
rect 21414 7040 21422 7104
rect 21486 7040 21502 7104
rect 21566 7040 21582 7104
rect 21646 7040 21662 7104
rect 21726 7040 21734 7104
rect 21414 6016 21734 7040
rect 21414 5952 21422 6016
rect 21486 5952 21502 6016
rect 21566 5952 21582 6016
rect 21646 5952 21662 6016
rect 21726 5952 21734 6016
rect 21414 4928 21734 5952
rect 21414 4864 21422 4928
rect 21486 4864 21502 4928
rect 21566 4864 21582 4928
rect 21646 4864 21662 4928
rect 21726 4864 21734 4928
rect 21414 3840 21734 4864
rect 21414 3776 21422 3840
rect 21486 3776 21502 3840
rect 21566 3776 21582 3840
rect 21646 3776 21662 3840
rect 21726 3776 21734 3840
rect 21414 2752 21734 3776
rect 21414 2688 21422 2752
rect 21486 2688 21502 2752
rect 21566 2688 21582 2752
rect 21646 2688 21662 2752
rect 21726 2688 21734 2752
rect 21414 2128 21734 2688
rect 25508 32672 25828 32688
rect 25508 32608 25516 32672
rect 25580 32608 25596 32672
rect 25660 32608 25676 32672
rect 25740 32608 25756 32672
rect 25820 32608 25828 32672
rect 25508 31584 25828 32608
rect 25508 31520 25516 31584
rect 25580 31520 25596 31584
rect 25660 31520 25676 31584
rect 25740 31520 25756 31584
rect 25820 31520 25828 31584
rect 25508 30496 25828 31520
rect 25508 30432 25516 30496
rect 25580 30432 25596 30496
rect 25660 30432 25676 30496
rect 25740 30432 25756 30496
rect 25820 30432 25828 30496
rect 25508 29408 25828 30432
rect 25508 29344 25516 29408
rect 25580 29344 25596 29408
rect 25660 29344 25676 29408
rect 25740 29344 25756 29408
rect 25820 29344 25828 29408
rect 25508 28320 25828 29344
rect 25508 28256 25516 28320
rect 25580 28256 25596 28320
rect 25660 28256 25676 28320
rect 25740 28256 25756 28320
rect 25820 28256 25828 28320
rect 25508 27232 25828 28256
rect 25508 27168 25516 27232
rect 25580 27168 25596 27232
rect 25660 27168 25676 27232
rect 25740 27168 25756 27232
rect 25820 27168 25828 27232
rect 25508 26144 25828 27168
rect 25508 26080 25516 26144
rect 25580 26080 25596 26144
rect 25660 26080 25676 26144
rect 25740 26080 25756 26144
rect 25820 26080 25828 26144
rect 25508 25056 25828 26080
rect 25508 24992 25516 25056
rect 25580 24992 25596 25056
rect 25660 24992 25676 25056
rect 25740 24992 25756 25056
rect 25820 24992 25828 25056
rect 25508 23968 25828 24992
rect 25508 23904 25516 23968
rect 25580 23904 25596 23968
rect 25660 23904 25676 23968
rect 25740 23904 25756 23968
rect 25820 23904 25828 23968
rect 25508 22880 25828 23904
rect 25508 22816 25516 22880
rect 25580 22816 25596 22880
rect 25660 22816 25676 22880
rect 25740 22816 25756 22880
rect 25820 22816 25828 22880
rect 25508 21792 25828 22816
rect 25508 21728 25516 21792
rect 25580 21728 25596 21792
rect 25660 21728 25676 21792
rect 25740 21728 25756 21792
rect 25820 21728 25828 21792
rect 25508 20704 25828 21728
rect 25508 20640 25516 20704
rect 25580 20640 25596 20704
rect 25660 20640 25676 20704
rect 25740 20640 25756 20704
rect 25820 20640 25828 20704
rect 25508 19616 25828 20640
rect 25508 19552 25516 19616
rect 25580 19552 25596 19616
rect 25660 19552 25676 19616
rect 25740 19552 25756 19616
rect 25820 19552 25828 19616
rect 25508 18528 25828 19552
rect 25508 18464 25516 18528
rect 25580 18464 25596 18528
rect 25660 18464 25676 18528
rect 25740 18464 25756 18528
rect 25820 18464 25828 18528
rect 25508 17440 25828 18464
rect 25508 17376 25516 17440
rect 25580 17376 25596 17440
rect 25660 17376 25676 17440
rect 25740 17376 25756 17440
rect 25820 17376 25828 17440
rect 25508 16352 25828 17376
rect 25508 16288 25516 16352
rect 25580 16288 25596 16352
rect 25660 16288 25676 16352
rect 25740 16288 25756 16352
rect 25820 16288 25828 16352
rect 25508 15264 25828 16288
rect 25508 15200 25516 15264
rect 25580 15200 25596 15264
rect 25660 15200 25676 15264
rect 25740 15200 25756 15264
rect 25820 15200 25828 15264
rect 25508 14176 25828 15200
rect 25508 14112 25516 14176
rect 25580 14112 25596 14176
rect 25660 14112 25676 14176
rect 25740 14112 25756 14176
rect 25820 14112 25828 14176
rect 25508 13088 25828 14112
rect 25508 13024 25516 13088
rect 25580 13024 25596 13088
rect 25660 13024 25676 13088
rect 25740 13024 25756 13088
rect 25820 13024 25828 13088
rect 25508 12000 25828 13024
rect 25508 11936 25516 12000
rect 25580 11936 25596 12000
rect 25660 11936 25676 12000
rect 25740 11936 25756 12000
rect 25820 11936 25828 12000
rect 25508 10912 25828 11936
rect 25508 10848 25516 10912
rect 25580 10848 25596 10912
rect 25660 10848 25676 10912
rect 25740 10848 25756 10912
rect 25820 10848 25828 10912
rect 25508 9824 25828 10848
rect 25508 9760 25516 9824
rect 25580 9760 25596 9824
rect 25660 9760 25676 9824
rect 25740 9760 25756 9824
rect 25820 9760 25828 9824
rect 25508 8736 25828 9760
rect 25508 8672 25516 8736
rect 25580 8672 25596 8736
rect 25660 8672 25676 8736
rect 25740 8672 25756 8736
rect 25820 8672 25828 8736
rect 25508 7648 25828 8672
rect 25508 7584 25516 7648
rect 25580 7584 25596 7648
rect 25660 7584 25676 7648
rect 25740 7584 25756 7648
rect 25820 7584 25828 7648
rect 25508 6560 25828 7584
rect 25508 6496 25516 6560
rect 25580 6496 25596 6560
rect 25660 6496 25676 6560
rect 25740 6496 25756 6560
rect 25820 6496 25828 6560
rect 25508 5472 25828 6496
rect 25508 5408 25516 5472
rect 25580 5408 25596 5472
rect 25660 5408 25676 5472
rect 25740 5408 25756 5472
rect 25820 5408 25828 5472
rect 25508 4384 25828 5408
rect 25508 4320 25516 4384
rect 25580 4320 25596 4384
rect 25660 4320 25676 4384
rect 25740 4320 25756 4384
rect 25820 4320 25828 4384
rect 25508 3296 25828 4320
rect 25508 3232 25516 3296
rect 25580 3232 25596 3296
rect 25660 3232 25676 3296
rect 25740 3232 25756 3296
rect 25820 3232 25828 3296
rect 25508 2208 25828 3232
rect 25508 2144 25516 2208
rect 25580 2144 25596 2208
rect 25660 2144 25676 2208
rect 25740 2144 25756 2208
rect 25820 2144 25828 2208
rect 25508 2128 25828 2144
rect 29602 32128 29922 32688
rect 29602 32064 29610 32128
rect 29674 32064 29690 32128
rect 29754 32064 29770 32128
rect 29834 32064 29850 32128
rect 29914 32064 29922 32128
rect 29602 31040 29922 32064
rect 29602 30976 29610 31040
rect 29674 30976 29690 31040
rect 29754 30976 29770 31040
rect 29834 30976 29850 31040
rect 29914 30976 29922 31040
rect 29602 29952 29922 30976
rect 29602 29888 29610 29952
rect 29674 29888 29690 29952
rect 29754 29888 29770 29952
rect 29834 29888 29850 29952
rect 29914 29888 29922 29952
rect 29602 28864 29922 29888
rect 29602 28800 29610 28864
rect 29674 28800 29690 28864
rect 29754 28800 29770 28864
rect 29834 28800 29850 28864
rect 29914 28800 29922 28864
rect 29602 27776 29922 28800
rect 29602 27712 29610 27776
rect 29674 27712 29690 27776
rect 29754 27712 29770 27776
rect 29834 27712 29850 27776
rect 29914 27712 29922 27776
rect 29602 26688 29922 27712
rect 29602 26624 29610 26688
rect 29674 26624 29690 26688
rect 29754 26624 29770 26688
rect 29834 26624 29850 26688
rect 29914 26624 29922 26688
rect 29602 25600 29922 26624
rect 29602 25536 29610 25600
rect 29674 25536 29690 25600
rect 29754 25536 29770 25600
rect 29834 25536 29850 25600
rect 29914 25536 29922 25600
rect 29602 24512 29922 25536
rect 29602 24448 29610 24512
rect 29674 24448 29690 24512
rect 29754 24448 29770 24512
rect 29834 24448 29850 24512
rect 29914 24448 29922 24512
rect 29602 23424 29922 24448
rect 29602 23360 29610 23424
rect 29674 23360 29690 23424
rect 29754 23360 29770 23424
rect 29834 23360 29850 23424
rect 29914 23360 29922 23424
rect 29602 22336 29922 23360
rect 29602 22272 29610 22336
rect 29674 22272 29690 22336
rect 29754 22272 29770 22336
rect 29834 22272 29850 22336
rect 29914 22272 29922 22336
rect 29602 21248 29922 22272
rect 29602 21184 29610 21248
rect 29674 21184 29690 21248
rect 29754 21184 29770 21248
rect 29834 21184 29850 21248
rect 29914 21184 29922 21248
rect 29602 20160 29922 21184
rect 29602 20096 29610 20160
rect 29674 20096 29690 20160
rect 29754 20096 29770 20160
rect 29834 20096 29850 20160
rect 29914 20096 29922 20160
rect 29602 19072 29922 20096
rect 29602 19008 29610 19072
rect 29674 19008 29690 19072
rect 29754 19008 29770 19072
rect 29834 19008 29850 19072
rect 29914 19008 29922 19072
rect 29602 17984 29922 19008
rect 29602 17920 29610 17984
rect 29674 17920 29690 17984
rect 29754 17920 29770 17984
rect 29834 17920 29850 17984
rect 29914 17920 29922 17984
rect 29602 16896 29922 17920
rect 29602 16832 29610 16896
rect 29674 16832 29690 16896
rect 29754 16832 29770 16896
rect 29834 16832 29850 16896
rect 29914 16832 29922 16896
rect 29602 15808 29922 16832
rect 29602 15744 29610 15808
rect 29674 15744 29690 15808
rect 29754 15744 29770 15808
rect 29834 15744 29850 15808
rect 29914 15744 29922 15808
rect 29602 14720 29922 15744
rect 29602 14656 29610 14720
rect 29674 14656 29690 14720
rect 29754 14656 29770 14720
rect 29834 14656 29850 14720
rect 29914 14656 29922 14720
rect 29602 13632 29922 14656
rect 29602 13568 29610 13632
rect 29674 13568 29690 13632
rect 29754 13568 29770 13632
rect 29834 13568 29850 13632
rect 29914 13568 29922 13632
rect 29602 12544 29922 13568
rect 29602 12480 29610 12544
rect 29674 12480 29690 12544
rect 29754 12480 29770 12544
rect 29834 12480 29850 12544
rect 29914 12480 29922 12544
rect 29602 11456 29922 12480
rect 29602 11392 29610 11456
rect 29674 11392 29690 11456
rect 29754 11392 29770 11456
rect 29834 11392 29850 11456
rect 29914 11392 29922 11456
rect 29602 10368 29922 11392
rect 29602 10304 29610 10368
rect 29674 10304 29690 10368
rect 29754 10304 29770 10368
rect 29834 10304 29850 10368
rect 29914 10304 29922 10368
rect 29602 9280 29922 10304
rect 29602 9216 29610 9280
rect 29674 9216 29690 9280
rect 29754 9216 29770 9280
rect 29834 9216 29850 9280
rect 29914 9216 29922 9280
rect 29602 8192 29922 9216
rect 29602 8128 29610 8192
rect 29674 8128 29690 8192
rect 29754 8128 29770 8192
rect 29834 8128 29850 8192
rect 29914 8128 29922 8192
rect 29602 7104 29922 8128
rect 29602 7040 29610 7104
rect 29674 7040 29690 7104
rect 29754 7040 29770 7104
rect 29834 7040 29850 7104
rect 29914 7040 29922 7104
rect 29602 6016 29922 7040
rect 29602 5952 29610 6016
rect 29674 5952 29690 6016
rect 29754 5952 29770 6016
rect 29834 5952 29850 6016
rect 29914 5952 29922 6016
rect 29602 4928 29922 5952
rect 29602 4864 29610 4928
rect 29674 4864 29690 4928
rect 29754 4864 29770 4928
rect 29834 4864 29850 4928
rect 29914 4864 29922 4928
rect 29602 3840 29922 4864
rect 29602 3776 29610 3840
rect 29674 3776 29690 3840
rect 29754 3776 29770 3840
rect 29834 3776 29850 3840
rect 29914 3776 29922 3840
rect 29602 2752 29922 3776
rect 29602 2688 29610 2752
rect 29674 2688 29690 2752
rect 29754 2688 29770 2752
rect 29834 2688 29850 2752
rect 29914 2688 29922 2752
rect 29602 2128 29922 2688
rect 33696 32672 34016 32688
rect 33696 32608 33704 32672
rect 33768 32608 33784 32672
rect 33848 32608 33864 32672
rect 33928 32608 33944 32672
rect 34008 32608 34016 32672
rect 33696 31584 34016 32608
rect 33696 31520 33704 31584
rect 33768 31520 33784 31584
rect 33848 31520 33864 31584
rect 33928 31520 33944 31584
rect 34008 31520 34016 31584
rect 33696 30496 34016 31520
rect 33696 30432 33704 30496
rect 33768 30432 33784 30496
rect 33848 30432 33864 30496
rect 33928 30432 33944 30496
rect 34008 30432 34016 30496
rect 33696 29408 34016 30432
rect 33696 29344 33704 29408
rect 33768 29344 33784 29408
rect 33848 29344 33864 29408
rect 33928 29344 33944 29408
rect 34008 29344 34016 29408
rect 33696 28320 34016 29344
rect 33696 28256 33704 28320
rect 33768 28256 33784 28320
rect 33848 28256 33864 28320
rect 33928 28256 33944 28320
rect 34008 28256 34016 28320
rect 33696 27232 34016 28256
rect 33696 27168 33704 27232
rect 33768 27168 33784 27232
rect 33848 27168 33864 27232
rect 33928 27168 33944 27232
rect 34008 27168 34016 27232
rect 33696 26144 34016 27168
rect 33696 26080 33704 26144
rect 33768 26080 33784 26144
rect 33848 26080 33864 26144
rect 33928 26080 33944 26144
rect 34008 26080 34016 26144
rect 33696 25056 34016 26080
rect 33696 24992 33704 25056
rect 33768 24992 33784 25056
rect 33848 24992 33864 25056
rect 33928 24992 33944 25056
rect 34008 24992 34016 25056
rect 33696 23968 34016 24992
rect 33696 23904 33704 23968
rect 33768 23904 33784 23968
rect 33848 23904 33864 23968
rect 33928 23904 33944 23968
rect 34008 23904 34016 23968
rect 33696 22880 34016 23904
rect 33696 22816 33704 22880
rect 33768 22816 33784 22880
rect 33848 22816 33864 22880
rect 33928 22816 33944 22880
rect 34008 22816 34016 22880
rect 33696 21792 34016 22816
rect 33696 21728 33704 21792
rect 33768 21728 33784 21792
rect 33848 21728 33864 21792
rect 33928 21728 33944 21792
rect 34008 21728 34016 21792
rect 33696 20704 34016 21728
rect 33696 20640 33704 20704
rect 33768 20640 33784 20704
rect 33848 20640 33864 20704
rect 33928 20640 33944 20704
rect 34008 20640 34016 20704
rect 33696 19616 34016 20640
rect 33696 19552 33704 19616
rect 33768 19552 33784 19616
rect 33848 19552 33864 19616
rect 33928 19552 33944 19616
rect 34008 19552 34016 19616
rect 33696 18528 34016 19552
rect 33696 18464 33704 18528
rect 33768 18464 33784 18528
rect 33848 18464 33864 18528
rect 33928 18464 33944 18528
rect 34008 18464 34016 18528
rect 33696 17440 34016 18464
rect 33696 17376 33704 17440
rect 33768 17376 33784 17440
rect 33848 17376 33864 17440
rect 33928 17376 33944 17440
rect 34008 17376 34016 17440
rect 33696 16352 34016 17376
rect 33696 16288 33704 16352
rect 33768 16288 33784 16352
rect 33848 16288 33864 16352
rect 33928 16288 33944 16352
rect 34008 16288 34016 16352
rect 33696 15264 34016 16288
rect 33696 15200 33704 15264
rect 33768 15200 33784 15264
rect 33848 15200 33864 15264
rect 33928 15200 33944 15264
rect 34008 15200 34016 15264
rect 33696 14176 34016 15200
rect 33696 14112 33704 14176
rect 33768 14112 33784 14176
rect 33848 14112 33864 14176
rect 33928 14112 33944 14176
rect 34008 14112 34016 14176
rect 33696 13088 34016 14112
rect 33696 13024 33704 13088
rect 33768 13024 33784 13088
rect 33848 13024 33864 13088
rect 33928 13024 33944 13088
rect 34008 13024 34016 13088
rect 33696 12000 34016 13024
rect 33696 11936 33704 12000
rect 33768 11936 33784 12000
rect 33848 11936 33864 12000
rect 33928 11936 33944 12000
rect 34008 11936 34016 12000
rect 33696 10912 34016 11936
rect 33696 10848 33704 10912
rect 33768 10848 33784 10912
rect 33848 10848 33864 10912
rect 33928 10848 33944 10912
rect 34008 10848 34016 10912
rect 33696 9824 34016 10848
rect 33696 9760 33704 9824
rect 33768 9760 33784 9824
rect 33848 9760 33864 9824
rect 33928 9760 33944 9824
rect 34008 9760 34016 9824
rect 33696 8736 34016 9760
rect 33696 8672 33704 8736
rect 33768 8672 33784 8736
rect 33848 8672 33864 8736
rect 33928 8672 33944 8736
rect 34008 8672 34016 8736
rect 33696 7648 34016 8672
rect 33696 7584 33704 7648
rect 33768 7584 33784 7648
rect 33848 7584 33864 7648
rect 33928 7584 33944 7648
rect 34008 7584 34016 7648
rect 33696 6560 34016 7584
rect 33696 6496 33704 6560
rect 33768 6496 33784 6560
rect 33848 6496 33864 6560
rect 33928 6496 33944 6560
rect 34008 6496 34016 6560
rect 33696 5472 34016 6496
rect 33696 5408 33704 5472
rect 33768 5408 33784 5472
rect 33848 5408 33864 5472
rect 33928 5408 33944 5472
rect 34008 5408 34016 5472
rect 33696 4384 34016 5408
rect 33696 4320 33704 4384
rect 33768 4320 33784 4384
rect 33848 4320 33864 4384
rect 33928 4320 33944 4384
rect 34008 4320 34016 4384
rect 33696 3296 34016 4320
rect 33696 3232 33704 3296
rect 33768 3232 33784 3296
rect 33848 3232 33864 3296
rect 33928 3232 33944 3296
rect 34008 3232 34016 3296
rect 33696 2208 34016 3232
rect 33696 2144 33704 2208
rect 33768 2144 33784 2208
rect 33848 2144 33864 2208
rect 33928 2144 33944 2208
rect 34008 2144 34016 2208
rect 33696 2128 34016 2144
use sky130_fd_sc_hd__and2b_1  _088_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _089_
timestamp 1688980957
transform -1 0 14996 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _090_
timestamp 1688980957
transform 1 0 15824 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _091_
timestamp 1688980957
transform -1 0 18676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _092_
timestamp 1688980957
transform -1 0 20884 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _093_
timestamp 1688980957
transform -1 0 21712 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _094_
timestamp 1688980957
transform -1 0 23460 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _095_
timestamp 1688980957
transform -1 0 26404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _096_
timestamp 1688980957
transform -1 0 27508 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _097_
timestamp 1688980957
transform -1 0 30084 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _098_
timestamp 1688980957
transform 1 0 23552 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _099_
timestamp 1688980957
transform 1 0 27416 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _100_
timestamp 1688980957
transform -1 0 31924 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _101_
timestamp 1688980957
transform 1 0 24564 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _102_
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _103_
timestamp 1688980957
transform -1 0 23276 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _104_
timestamp 1688980957
transform -1 0 24932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _105_
timestamp 1688980957
transform -1 0 26864 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _106_
timestamp 1688980957
transform -1 0 27968 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _107_
timestamp 1688980957
transform -1 0 29440 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _108_
timestamp 1688980957
transform -1 0 31924 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _109_
timestamp 1688980957
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _110_
timestamp 1688980957
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _111_
timestamp 1688980957
transform 1 0 25576 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _112_
timestamp 1688980957
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _113_
timestamp 1688980957
transform 1 0 29624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _114_
timestamp 1688980957
transform 1 0 29992 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _115_
timestamp 1688980957
transform 1 0 30728 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _116_
timestamp 1688980957
transform 1 0 30820 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _117_
timestamp 1688980957
transform 1 0 29992 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _118_
timestamp 1688980957
transform 1 0 29992 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _119_
timestamp 1688980957
transform 1 0 30728 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _120_
timestamp 1688980957
transform 1 0 30268 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _121_
timestamp 1688980957
transform 1 0 31556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _122_
timestamp 1688980957
transform 1 0 30728 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _123_
timestamp 1688980957
transform 1 0 30820 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _124_
timestamp 1688980957
transform 1 0 30820 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _125_
timestamp 1688980957
transform 1 0 29256 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _126_
timestamp 1688980957
transform 1 0 29624 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _127_
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _128_
timestamp 1688980957
transform 1 0 28888 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _129_
timestamp 1688980957
transform 1 0 26864 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _130_
timestamp 1688980957
transform 1 0 27784 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _131_
timestamp 1688980957
transform 1 0 18584 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _132_
timestamp 1688980957
transform 1 0 9568 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _133_
timestamp 1688980957
transform 1 0 7544 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _134_
timestamp 1688980957
transform 1 0 8096 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _135_
timestamp 1688980957
transform -1 0 12052 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _136_
timestamp 1688980957
transform 1 0 10856 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _137_
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _138_
timestamp 1688980957
transform -1 0 16008 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _139_
timestamp 1688980957
transform -1 0 17388 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _140_
timestamp 1688980957
transform 1 0 15180 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _141_
timestamp 1688980957
transform -1 0 11040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _142_
timestamp 1688980957
transform -1 0 5060 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _143_
timestamp 1688980957
transform -1 0 4876 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _144_
timestamp 1688980957
transform -1 0 4876 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _145_
timestamp 1688980957
transform -1 0 4876 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _146_
timestamp 1688980957
transform -1 0 5244 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _147_
timestamp 1688980957
transform -1 0 4140 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _148_
timestamp 1688980957
transform -1 0 5244 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _149_
timestamp 1688980957
transform -1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _150_
timestamp 1688980957
transform -1 0 5796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _151_
timestamp 1688980957
transform -1 0 5060 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _152_
timestamp 1688980957
transform -1 0 4140 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _153_
timestamp 1688980957
transform -1 0 5060 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _154_
timestamp 1688980957
transform -1 0 4508 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _155_
timestamp 1688980957
transform -1 0 4140 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _156_
timestamp 1688980957
transform -1 0 4232 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _157_
timestamp 1688980957
transform -1 0 5060 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _158_
timestamp 1688980957
transform -1 0 4876 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _159_
timestamp 1688980957
transform -1 0 5796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _160_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3680 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _161_
timestamp 1688980957
transform -1 0 15640 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _162_
timestamp 1688980957
transform -1 0 18584 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _163_
timestamp 1688980957
transform 1 0 19320 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _164_
timestamp 1688980957
transform 1 0 18124 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _165_
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _166_
timestamp 1688980957
transform -1 0 4324 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _167_
timestamp 1688980957
transform -1 0 4876 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _168_
timestamp 1688980957
transform -1 0 5060 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _169_
timestamp 1688980957
transform -1 0 6532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _170_
timestamp 1688980957
transform -1 0 4324 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _171_
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _172_
timestamp 1688980957
transform -1 0 6256 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _173_
timestamp 1688980957
transform -1 0 8832 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _174_
timestamp 1688980957
transform -1 0 10856 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _175_
timestamp 1688980957
transform 1 0 9016 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _176_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13156 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _177_
timestamp 1688980957
transform -1 0 14628 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _178_
timestamp 1688980957
transform -1 0 16468 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _179_
timestamp 1688980957
transform -1 0 18124 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _180_
timestamp 1688980957
transform -1 0 20332 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _181_
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _182_
timestamp 1688980957
transform -1 0 23552 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _183_
timestamp 1688980957
transform -1 0 25116 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _184_
timestamp 1688980957
transform 1 0 25300 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _185_
timestamp 1688980957
transform -1 0 28428 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _186_
timestamp 1688980957
transform -1 0 31372 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _187_
timestamp 1688980957
transform -1 0 31004 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _188_
timestamp 1688980957
transform -1 0 32476 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _189_
timestamp 1688980957
transform 1 0 25392 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _190_
timestamp 1688980957
transform -1 0 26220 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _191_
timestamp 1688980957
transform 1 0 22172 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _192_
timestamp 1688980957
transform 1 0 23368 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _193_
timestamp 1688980957
transform -1 0 26404 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _194_
timestamp 1688980957
transform -1 0 28428 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _195_
timestamp 1688980957
transform -1 0 29348 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _196_
timestamp 1688980957
transform -1 0 31004 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _197_
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _198_
timestamp 1688980957
transform 1 0 28704 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _199_
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _200_
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _201_
timestamp 1688980957
transform 1 0 31648 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _202_
timestamp 1688980957
transform 1 0 31648 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _203_
timestamp 1688980957
transform 1 0 31648 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _204_
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _205_
timestamp 1688980957
transform 1 0 31648 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _206_
timestamp 1688980957
transform 1 0 31648 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _207_
timestamp 1688980957
transform 1 0 31648 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _208_
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _209_
timestamp 1688980957
transform 1 0 31648 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _210_
timestamp 1688980957
transform 1 0 31648 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _211_
timestamp 1688980957
transform 1 0 31648 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _212_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _213_
timestamp 1688980957
transform 1 0 31648 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _214_
timestamp 1688980957
transform 1 0 31648 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _215_
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _216_
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _217_
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _218_
timestamp 1688980957
transform 1 0 31648 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _219_
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _220_
timestamp 1688980957
transform 1 0 10120 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _221_
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _222_
timestamp 1688980957
transform 1 0 9108 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _223_
timestamp 1688980957
transform 1 0 8464 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _224_
timestamp 1688980957
transform -1 0 13064 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _225_
timestamp 1688980957
transform -1 0 14628 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _226_
timestamp 1688980957
transform -1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _227_
timestamp 1688980957
transform 1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _228_
timestamp 1688980957
transform 1 0 17020 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _229_
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _230_
timestamp 1688980957
transform 1 0 2116 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _231_
timestamp 1688980957
transform 1 0 1748 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _233_
timestamp 1688980957
transform 1 0 1748 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1688980957
transform 1 0 1748 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _235_
timestamp 1688980957
transform 1 0 2852 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _236_
timestamp 1688980957
transform 1 0 1748 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _237_
timestamp 1688980957
transform 1 0 1748 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _238_
timestamp 1688980957
transform 1 0 2852 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _240_
timestamp 1688980957
transform -1 0 4324 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _241_
timestamp 1688980957
transform 1 0 1748 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _242_
timestamp 1688980957
transform 1 0 1748 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _243_
timestamp 1688980957
transform 1 0 1748 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _244_
timestamp 1688980957
transform 1 0 1748 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _245_
timestamp 1688980957
transform 1 0 1748 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _246_
timestamp 1688980957
transform 1 0 1748 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _247_
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _248_
timestamp 1688980957
transform -1 0 3220 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _249_
timestamp 1688980957
transform -1 0 13524 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _250_
timestamp 1688980957
transform -1 0 18676 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _251_
timestamp 1688980957
transform -1 0 20332 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _252_
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _253_
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _254_
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _255_
timestamp 1688980957
transform 1 0 1932 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _256_
timestamp 1688980957
transform 1 0 1748 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _257_
timestamp 1688980957
transform 1 0 1748 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _258_
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _259_
timestamp 1688980957
transform -1 0 5704 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _260_
timestamp 1688980957
transform 1 0 5520 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _261_
timestamp 1688980957
transform -1 0 8280 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _262_
timestamp 1688980957
transform -1 0 10304 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _263_
timestamp 1688980957
transform -1 0 12328 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A_N dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A_N
timestamp 1688980957
transform 1 0 15180 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A_N
timestamp 1688980957
transform 1 0 15640 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A_N
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A_N
timestamp 1688980957
transform -1 0 21436 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A_N
timestamp 1688980957
transform 1 0 21988 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A_N
timestamp 1688980957
transform 1 0 23460 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A_N
timestamp 1688980957
transform -1 0 27232 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A_N
timestamp 1688980957
transform 1 0 28152 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A_N
timestamp 1688980957
transform 1 0 30084 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A_N
timestamp 1688980957
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A_N
timestamp 1688980957
transform 1 0 27968 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A_N
timestamp 1688980957
transform -1 0 31372 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A_N
timestamp 1688980957
transform -1 0 25484 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A_N
timestamp 1688980957
transform 1 0 25392 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A_N
timestamp 1688980957
transform 1 0 23276 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A_N
timestamp 1688980957
transform 1 0 25208 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A_N
timestamp 1688980957
transform 1 0 29256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A_N
timestamp 1688980957
transform 1 0 28888 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A_N
timestamp 1688980957
transform 1 0 29716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A_N
timestamp 1688980957
transform 1 0 31188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A_N
timestamp 1688980957
transform 1 0 30544 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A_N
timestamp 1688980957
transform 1 0 20976 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A_N
timestamp 1688980957
transform 1 0 25760 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A_N
timestamp 1688980957
transform 1 0 28704 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A_N
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A_N
timestamp 1688980957
transform 1 0 29808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A_N
timestamp 1688980957
transform 1 0 30544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A_N
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A_N
timestamp 1688980957
transform 1 0 29808 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A_N
timestamp 1688980957
transform 1 0 29808 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A_N
timestamp 1688980957
transform 1 0 30544 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A_N
timestamp 1688980957
transform 1 0 31004 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A_N
timestamp 1688980957
transform 1 0 31372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A_N
timestamp 1688980957
transform 1 0 30544 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A_N
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A_N
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A_N
timestamp 1688980957
transform 1 0 29072 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A_N
timestamp 1688980957
transform 1 0 28704 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A_N
timestamp 1688980957
transform -1 0 26864 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A_N
timestamp 1688980957
transform 1 0 28704 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A_N
timestamp 1688980957
transform 1 0 27416 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A_N
timestamp 1688980957
transform 1 0 28336 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A_N
timestamp 1688980957
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A_N
timestamp 1688980957
transform 1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A_N
timestamp 1688980957
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A_N
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A_N
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A_N
timestamp 1688980957
transform -1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A_N
timestamp 1688980957
transform -1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A_N
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A_N
timestamp 1688980957
transform 1 0 17572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A_N
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A_N
timestamp 1688980957
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A_N
timestamp 1688980957
transform -1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A_N
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A_N
timestamp 1688980957
transform 1 0 5244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A_N
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A_N
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A_N
timestamp 1688980957
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A_N
timestamp 1688980957
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A_N
timestamp 1688980957
transform 1 0 5060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A_N
timestamp 1688980957
transform 1 0 15640 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A_N
timestamp 1688980957
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A_N
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A_N
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A_N
timestamp 1688980957
transform 1 0 11868 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A_N
timestamp 1688980957
transform 1 0 5428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A_N
timestamp 1688980957
transform 1 0 5060 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A_N
timestamp 1688980957
transform 1 0 9108 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A_N
timestamp 1688980957
transform 1 0 11040 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A_N
timestamp 1688980957
transform -1 0 9936 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__CLK
timestamp 1688980957
transform -1 0 18308 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__CLK
timestamp 1688980957
transform -1 0 21068 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__181__CLK
timestamp 1688980957
transform 1 0 22356 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__CLK
timestamp 1688980957
transform -1 0 22448 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__183__CLK
timestamp 1688980957
transform -1 0 25760 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__CLK
timestamp 1688980957
transform -1 0 28704 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__CLK
timestamp 1688980957
transform -1 0 27324 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__CLK
timestamp 1688980957
transform 1 0 22264 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__CLK
timestamp 1688980957
transform 1 0 21988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__CLK
timestamp 1688980957
transform 1 0 24840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__CLK
timestamp 1688980957
transform -1 0 28152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__CLK
timestamp 1688980957
transform -1 0 30728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__CLK
timestamp 1688980957
transform 1 0 31096 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__CLK
timestamp 1688980957
transform 1 0 29992 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__CLK
timestamp 1688980957
transform -1 0 23276 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__CLK
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__CLK
timestamp 1688980957
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__CLK
timestamp 1688980957
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 9844 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 7268 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 9844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 25852 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 28428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 25852 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_wb_clk_i_A
timestamp 1688980957
transform 1 0 28428 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_A
timestamp 1688980957
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout91_A
timestamp 1688980957
transform 1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout92_A
timestamp 1688980957
transform 1 0 16192 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout93_A
timestamp 1688980957
transform -1 0 26864 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout94_A
timestamp 1688980957
transform 1 0 30636 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout95_A
timestamp 1688980957
transform 1 0 27968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19136 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_wb_clk_i
timestamp 1688980957
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_wb_clk_i
timestamp 1688980957
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_wb_clk_i
timestamp 1688980957
transform -1 0 7084 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_wb_clk_i
timestamp 1688980957
transform -1 0 9660 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_wb_clk_i
timestamp 1688980957
transform -1 0 27876 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_wb_clk_i
timestamp 1688980957
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_wb_clk_i
timestamp 1688980957
transform 1 0 26036 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_wb_clk_i
timestamp 1688980957
transform 1 0 28612 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout90 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout91
timestamp 1688980957
transform -1 0 1932 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout92 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16008 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout93
timestamp 1688980957
transform 1 0 27048 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout94 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30820 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout95
timestamp 1688980957
transform 1 0 27416 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout96
timestamp 1688980957
transform -1 0 32016 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_32 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_44
timestamp 1688980957
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_69 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_206 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_214 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_262
timestamp 1688980957
transform 1 0 25208 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_266
timestamp 1688980957
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_290
timestamp 1688980957
transform 1 0 27784 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_294
timestamp 1688980957
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_318
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_322
timestamp 1688980957
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_19
timestamp 1688980957
transform 1 0 2852 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_31
timestamp 1688980957
transform 1 0 3956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_63
timestamp 1688980957
transform 1 0 6900 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_121
timestamp 1688980957
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_147 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_151
timestamp 1688980957
transform 1 0 14996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_177
timestamp 1688980957
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_187
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_199
timestamp 1688980957
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_216
timestamp 1688980957
transform 1 0 20976 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_229
timestamp 1688980957
transform 1 0 22172 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 1688980957
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_52
timestamp 1688980957
transform 1 0 5888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_58
timestamp 1688980957
transform 1 0 6440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_68
timestamp 1688980957
transform 1 0 7360 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_74
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_89
timestamp 1688980957
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_138
timestamp 1688980957
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_205
timestamp 1688980957
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_217
timestamp 1688980957
transform 1 0 21068 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_225
timestamp 1688980957
transform 1 0 21804 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_300
timestamp 1688980957
transform 1 0 28704 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_304
timestamp 1688980957
transform 1 0 29072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_318
timestamp 1688980957
transform 1 0 30360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_322
timestamp 1688980957
transform 1 0 30728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_326
timestamp 1688980957
transform 1 0 31096 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_329
timestamp 1688980957
transform 1 0 31372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_341
timestamp 1688980957
transform 1 0 32476 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_9
timestamp 1688980957
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_19
timestamp 1688980957
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_31
timestamp 1688980957
transform 1 0 3956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_43
timestamp 1688980957
transform 1 0 5060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_117
timestamp 1688980957
transform 1 0 11868 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_121
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_139
timestamp 1688980957
transform 1 0 13892 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_148
timestamp 1688980957
transform 1 0 14720 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_154
timestamp 1688980957
transform 1 0 15272 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_164
timestamp 1688980957
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_178
timestamp 1688980957
transform 1 0 17480 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_184
timestamp 1688980957
transform 1 0 18032 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_201
timestamp 1688980957
transform 1 0 19596 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_213
timestamp 1688980957
transform 1 0 20700 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_221
timestamp 1688980957
transform 1 0 21436 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_233
timestamp 1688980957
transform 1 0 22540 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_289
timestamp 1688980957
transform 1 0 27692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_307
timestamp 1688980957
transform 1 0 29348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_333
timestamp 1688980957
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_346
timestamp 1688980957
transform 1 0 32936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_352
timestamp 1688980957
transform 1 0 33488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 1688980957
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_103
timestamp 1688980957
transform 1 0 10580 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_120
timestamp 1688980957
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1688980957
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_147
timestamp 1688980957
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_162
timestamp 1688980957
transform 1 0 16008 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1688980957
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_241
timestamp 1688980957
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_317
timestamp 1688980957
transform 1 0 30268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_329
timestamp 1688980957
transform 1 0 31372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_336
timestamp 1688980957
transform 1 0 32016 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_346
timestamp 1688980957
transform 1 0 32936 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_352
timestamp 1688980957
transform 1 0 33488 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_33
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_37
timestamp 1688980957
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_49
timestamp 1688980957
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_75
timestamp 1688980957
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_98
timestamp 1688980957
transform 1 0 10120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1688980957
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_121
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_130
timestamp 1688980957
transform 1 0 13064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_140
timestamp 1688980957
transform 1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_144
timestamp 1688980957
transform 1 0 14352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_148
timestamp 1688980957
transform 1 0 14720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_152
timestamp 1688980957
transform 1 0 15088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_159
timestamp 1688980957
transform 1 0 15732 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_163
timestamp 1688980957
transform 1 0 16100 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_189
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_201
timestamp 1688980957
transform 1 0 19596 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_213
timestamp 1688980957
transform 1 0 20700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_221
timestamp 1688980957
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_243
timestamp 1688980957
transform 1 0 23460 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_265
timestamp 1688980957
transform 1 0 25484 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_297
timestamp 1688980957
transform 1 0 28428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_332
timestamp 1688980957
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_37
timestamp 1688980957
transform 1 0 4508 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_49
timestamp 1688980957
transform 1 0 5612 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_61
timestamp 1688980957
transform 1 0 6716 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_73
timestamp 1688980957
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_81
timestamp 1688980957
transform 1 0 8556 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_102
timestamp 1688980957
transform 1 0 10488 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_110
timestamp 1688980957
transform 1 0 11224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_119
timestamp 1688980957
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_123
timestamp 1688980957
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_135
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_257
timestamp 1688980957
transform 1 0 24748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_260
timestamp 1688980957
transform 1 0 25024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_264
timestamp 1688980957
transform 1 0 25392 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_337
timestamp 1688980957
transform 1 0 32108 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_343
timestamp 1688980957
transform 1 0 32660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_47
timestamp 1688980957
transform 1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_89
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_102
timestamp 1688980957
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_277
timestamp 1688980957
transform 1 0 26588 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_23
timestamp 1688980957
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_45
timestamp 1688980957
transform 1 0 5244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_57
timestamp 1688980957
transform 1 0 6348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_69
timestamp 1688980957
transform 1 0 7452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_81
timestamp 1688980957
transform 1 0 8556 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_285
timestamp 1688980957
transform 1 0 27324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_330
timestamp 1688980957
transform 1 0 31464 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_336
timestamp 1688980957
transform 1 0 32016 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_43
timestamp 1688980957
transform 1 0 5060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_178
timestamp 1688980957
transform 1 0 17480 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_190
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_202
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_214
timestamp 1688980957
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1688980957
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_289
timestamp 1688980957
transform 1 0 27692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_294
timestamp 1688980957
transform 1 0 28152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_346
timestamp 1688980957
transform 1 0 32936 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_352
timestamp 1688980957
transform 1 0 33488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_43
timestamp 1688980957
transform 1 0 5060 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_47
timestamp 1688980957
transform 1 0 5428 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_59
timestamp 1688980957
transform 1 0 6532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_71
timestamp 1688980957
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_297
timestamp 1688980957
transform 1 0 28428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_348
timestamp 1688980957
transform 1 0 33120 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_352
timestamp 1688980957
transform 1 0 33488 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_37
timestamp 1688980957
transform 1 0 4508 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_41
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1688980957
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_310
timestamp 1688980957
transform 1 0 29624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_346
timestamp 1688980957
transform 1 0 32936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_352
timestamp 1688980957
transform 1 0 33488 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_37
timestamp 1688980957
transform 1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_45
timestamp 1688980957
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_56
timestamp 1688980957
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_68
timestamp 1688980957
transform 1 0 7360 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1688980957
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_201
timestamp 1688980957
transform 1 0 19596 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_210
timestamp 1688980957
transform 1 0 20424 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_222
timestamp 1688980957
transform 1 0 21528 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_234
timestamp 1688980957
transform 1 0 22632 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_246
timestamp 1688980957
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_315
timestamp 1688980957
transform 1 0 30084 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_348
timestamp 1688980957
transform 1 0 33120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_352
timestamp 1688980957
transform 1 0 33488 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_37
timestamp 1688980957
transform 1 0 4508 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_49
timestamp 1688980957
transform 1 0 5612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_155
timestamp 1688980957
transform 1 0 15364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_260
timestamp 1688980957
transform 1 0 25024 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_272
timestamp 1688980957
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_289
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_301
timestamp 1688980957
transform 1 0 28796 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_346
timestamp 1688980957
transform 1 0 32936 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_352
timestamp 1688980957
transform 1 0 33488 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1688980957
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_69
timestamp 1688980957
transform 1 0 7452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_164
timestamp 1688980957
transform 1 0 16192 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_176
timestamp 1688980957
transform 1 0 17296 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_188
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_291
timestamp 1688980957
transform 1 0 27876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_303
timestamp 1688980957
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_315
timestamp 1688980957
transform 1 0 30084 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_348
timestamp 1688980957
transform 1 0 33120 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_352
timestamp 1688980957
transform 1 0 33488 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_19
timestamp 1688980957
transform 1 0 2852 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_34
timestamp 1688980957
transform 1 0 4232 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_38
timestamp 1688980957
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_50
timestamp 1688980957
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_97
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1688980957
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_319
timestamp 1688980957
transform 1 0 30452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_23
timestamp 1688980957
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_37
timestamp 1688980957
transform 1 0 4508 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_49
timestamp 1688980957
transform 1 0 5612 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_61
timestamp 1688980957
transform 1 0 6716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_73
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_317
timestamp 1688980957
transform 1 0 30268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_322
timestamp 1688980957
transform 1 0 30728 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_328
timestamp 1688980957
transform 1 0 31280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_346
timestamp 1688980957
transform 1 0 32936 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_352
timestamp 1688980957
transform 1 0 33488 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_43
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_141
timestamp 1688980957
transform 1 0 14076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_153
timestamp 1688980957
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 1688980957
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_197
timestamp 1688980957
transform 1 0 19228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_206
timestamp 1688980957
transform 1 0 20056 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_218
timestamp 1688980957
transform 1 0 21160 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_317
timestamp 1688980957
transform 1 0 30268 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_9
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_43
timestamp 1688980957
transform 1 0 5060 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_54
timestamp 1688980957
transform 1 0 6072 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_66
timestamp 1688980957
transform 1 0 7176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_78
timestamp 1688980957
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_105
timestamp 1688980957
transform 1 0 10764 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_117
timestamp 1688980957
transform 1 0 11868 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_129
timestamp 1688980957
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_137
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_261
timestamp 1688980957
transform 1 0 25116 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_273
timestamp 1688980957
transform 1 0 26220 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_285
timestamp 1688980957
transform 1 0 27324 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_297
timestamp 1688980957
transform 1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_53
timestamp 1688980957
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_246
timestamp 1688980957
transform 1 0 23736 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_258
timestamp 1688980957
transform 1 0 24840 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_270
timestamp 1688980957
transform 1 0 25944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_278
timestamp 1688980957
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_325
timestamp 1688980957
transform 1 0 31004 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_346
timestamp 1688980957
transform 1 0 32936 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_352
timestamp 1688980957
transform 1 0 33488 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_37
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_49
timestamp 1688980957
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_61
timestamp 1688980957
transform 1 0 6716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_73
timestamp 1688980957
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1688980957
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_101
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_108
timestamp 1688980957
transform 1 0 11040 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_112
timestamp 1688980957
transform 1 0 11408 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_124
timestamp 1688980957
transform 1 0 12512 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_136
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_206
timestamp 1688980957
transform 1 0 20056 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_218
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_230
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_242
timestamp 1688980957
transform 1 0 23368 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1688980957
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_315
timestamp 1688980957
transform 1 0 30084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_348
timestamp 1688980957
transform 1 0 33120 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_352
timestamp 1688980957
transform 1 0 33488 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_9
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_41
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_45
timestamp 1688980957
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_53
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_209
timestamp 1688980957
transform 1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_213
timestamp 1688980957
transform 1 0 20700 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 1688980957
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_311
timestamp 1688980957
transform 1 0 29716 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_346
timestamp 1688980957
transform 1 0 32936 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_352
timestamp 1688980957
transform 1 0 33488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_45
timestamp 1688980957
transform 1 0 5244 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_49
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_61
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_73
timestamp 1688980957
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1688980957
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_115
timestamp 1688980957
transform 1 0 11684 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_119
timestamp 1688980957
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_131
timestamp 1688980957
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_177
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_185
timestamp 1688980957
transform 1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_213
timestamp 1688980957
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_217
timestamp 1688980957
transform 1 0 21068 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_229
timestamp 1688980957
transform 1 0 22172 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_241
timestamp 1688980957
transform 1 0 23276 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_315
timestamp 1688980957
transform 1 0 30084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_348
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_352
timestamp 1688980957
transform 1 0 33488 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_25
timestamp 1688980957
transform 1 0 3404 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_43
timestamp 1688980957
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_153
timestamp 1688980957
transform 1 0 15180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_165
timestamp 1688980957
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_191
timestamp 1688980957
transform 1 0 18676 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_195
timestamp 1688980957
transform 1 0 19044 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_204
timestamp 1688980957
transform 1 0 19872 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_208
timestamp 1688980957
transform 1 0 20240 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_220
timestamp 1688980957
transform 1 0 21344 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_311
timestamp 1688980957
transform 1 0 29716 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_346
timestamp 1688980957
transform 1 0 32936 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_352
timestamp 1688980957
transform 1 0 33488 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_19
timestamp 1688980957
transform 1 0 2852 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_45
timestamp 1688980957
transform 1 0 5244 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_57
timestamp 1688980957
transform 1 0 6348 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_71
timestamp 1688980957
transform 1 0 7636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_261
timestamp 1688980957
transform 1 0 25116 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_315
timestamp 1688980957
transform 1 0 30084 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_348
timestamp 1688980957
transform 1 0 33120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_352
timestamp 1688980957
transform 1 0 33488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_33
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_43
timestamp 1688980957
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1688980957
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_23
timestamp 1688980957
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_43
timestamp 1688980957
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_47
timestamp 1688980957
transform 1 0 5428 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_59
timestamp 1688980957
transform 1 0 6532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_71
timestamp 1688980957
transform 1 0 7636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_208
timestamp 1688980957
transform 1 0 20240 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_220
timestamp 1688980957
transform 1 0 21344 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_224
timestamp 1688980957
transform 1 0 21712 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_236
timestamp 1688980957
transform 1 0 22816 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_248
timestamp 1688980957
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_346
timestamp 1688980957
transform 1 0 32936 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_352
timestamp 1688980957
transform 1 0 33488 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_23
timestamp 1688980957
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_43
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_55
timestamp 1688980957
transform 1 0 6164 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_67
timestamp 1688980957
transform 1 0 7268 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_79
timestamp 1688980957
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_173
timestamp 1688980957
transform 1 0 17020 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_237
timestamp 1688980957
transform 1 0 22908 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_241
timestamp 1688980957
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1688980957
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_261
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_273
timestamp 1688980957
transform 1 0 26220 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_285
timestamp 1688980957
transform 1 0 27324 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_297
timestamp 1688980957
transform 1 0 28428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_305
timestamp 1688980957
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_9
timestamp 1688980957
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_41
timestamp 1688980957
transform 1 0 4876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_53
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1688980957
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_323
timestamp 1688980957
transform 1 0 30820 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_327
timestamp 1688980957
transform 1 0 31188 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_346
timestamp 1688980957
transform 1 0 32936 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_352
timestamp 1688980957
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_7
timestamp 1688980957
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_51
timestamp 1688980957
transform 1 0 5796 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_63
timestamp 1688980957
transform 1 0 6900 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_75
timestamp 1688980957
transform 1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_183
timestamp 1688980957
transform 1 0 17940 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_190
timestamp 1688980957
transform 1 0 18584 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1688980957
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_348
timestamp 1688980957
transform 1 0 33120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_352
timestamp 1688980957
transform 1 0 33488 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_41
timestamp 1688980957
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_285
timestamp 1688980957
transform 1 0 27324 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_297
timestamp 1688980957
transform 1 0 28428 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_309
timestamp 1688980957
transform 1 0 29532 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_321
timestamp 1688980957
transform 1 0 30636 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_327
timestamp 1688980957
transform 1 0 31188 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_23
timestamp 1688980957
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_37
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_49
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_61
timestamp 1688980957
transform 1 0 6716 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_73
timestamp 1688980957
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_173
timestamp 1688980957
transform 1 0 17020 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_191
timestamp 1688980957
transform 1 0 18676 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_346
timestamp 1688980957
transform 1 0 32936 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_352
timestamp 1688980957
transform 1 0 33488 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_9
timestamp 1688980957
transform 1 0 1932 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_19
timestamp 1688980957
transform 1 0 2852 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_28
timestamp 1688980957
transform 1 0 3680 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_40
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_52
timestamp 1688980957
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_325
timestamp 1688980957
transform 1 0 31004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_346
timestamp 1688980957
transform 1 0 32936 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_352
timestamp 1688980957
transform 1 0 33488 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_23
timestamp 1688980957
transform 1 0 3220 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_37
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_69
timestamp 1688980957
transform 1 0 7452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_81
timestamp 1688980957
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1688980957
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_348
timestamp 1688980957
transform 1 0 33120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_352
timestamp 1688980957
transform 1 0 33488 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_41
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_317
timestamp 1688980957
transform 1 0 30268 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_23
timestamp 1688980957
transform 1 0 3220 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_37
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_49
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_61
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_73
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_348
timestamp 1688980957
transform 1 0 33120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_352
timestamp 1688980957
transform 1 0 33488 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_45
timestamp 1688980957
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 1688980957
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_289
timestamp 1688980957
transform 1 0 27692 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_299
timestamp 1688980957
transform 1 0 28612 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_311
timestamp 1688980957
transform 1 0 29716 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_319
timestamp 1688980957
transform 1 0 30452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_346
timestamp 1688980957
transform 1 0 32936 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_352
timestamp 1688980957
transform 1 0 33488 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_9
timestamp 1688980957
transform 1 0 1932 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_19
timestamp 1688980957
transform 1 0 2852 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_43
timestamp 1688980957
transform 1 0 5060 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_55
timestamp 1688980957
transform 1 0 6164 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_67
timestamp 1688980957
transform 1 0 7268 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_79
timestamp 1688980957
transform 1 0 8372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_186
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_194
timestamp 1688980957
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_291
timestamp 1688980957
transform 1 0 27876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_303
timestamp 1688980957
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_346
timestamp 1688980957
transform 1 0 32936 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_352
timestamp 1688980957
transform 1 0 33488 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_35
timestamp 1688980957
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_47
timestamp 1688980957
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_97
timestamp 1688980957
transform 1 0 10028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_109
timestamp 1688980957
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_289
timestamp 1688980957
transform 1 0 27692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_319
timestamp 1688980957
transform 1 0 30452 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_9
timestamp 1688980957
transform 1 0 1932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_19
timestamp 1688980957
transform 1 0 2852 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_37
timestamp 1688980957
transform 1 0 4508 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_49
timestamp 1688980957
transform 1 0 5612 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_61
timestamp 1688980957
transform 1 0 6716 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_73
timestamp 1688980957
transform 1 0 7820 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_81
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_157
timestamp 1688980957
transform 1 0 15548 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_160
timestamp 1688980957
transform 1 0 15824 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_172
timestamp 1688980957
transform 1 0 16928 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_184
timestamp 1688980957
transform 1 0 18032 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_33
timestamp 1688980957
transform 1 0 4140 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_45
timestamp 1688980957
transform 1 0 5244 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_135
timestamp 1688980957
transform 1 0 13524 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_147
timestamp 1688980957
transform 1 0 14628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_151
timestamp 1688980957
transform 1 0 14996 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_162
timestamp 1688980957
transform 1 0 16008 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_166
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_346
timestamp 1688980957
transform 1 0 32936 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_352
timestamp 1688980957
transform 1 0 33488 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_37
timestamp 1688980957
transform 1 0 4508 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_49
timestamp 1688980957
transform 1 0 5612 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_61
timestamp 1688980957
transform 1 0 6716 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_73
timestamp 1688980957
transform 1 0 7820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_81
timestamp 1688980957
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_297
timestamp 1688980957
transform 1 0 28428 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_313
timestamp 1688980957
transform 1 0 29900 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_348
timestamp 1688980957
transform 1 0 33120 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_352
timestamp 1688980957
transform 1 0 33488 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_45
timestamp 1688980957
transform 1 0 5244 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_53
timestamp 1688980957
transform 1 0 5980 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_178
timestamp 1688980957
transform 1 0 17480 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_190
timestamp 1688980957
transform 1 0 18584 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_202
timestamp 1688980957
transform 1 0 19688 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_214
timestamp 1688980957
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1688980957
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_299
timestamp 1688980957
transform 1 0 28612 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_302
timestamp 1688980957
transform 1 0 28888 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_346
timestamp 1688980957
transform 1 0 32936 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_352
timestamp 1688980957
transform 1 0 33488 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_51
timestamp 1688980957
transform 1 0 5796 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_63
timestamp 1688980957
transform 1 0 6900 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_75
timestamp 1688980957
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_187
timestamp 1688980957
transform 1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_294
timestamp 1688980957
transform 1 0 28152 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_298
timestamp 1688980957
transform 1 0 28520 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_348
timestamp 1688980957
transform 1 0 33120 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_352
timestamp 1688980957
transform 1 0 33488 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_9
timestamp 1688980957
transform 1 0 1932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_49
timestamp 1688980957
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_66
timestamp 1688980957
transform 1 0 7176 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_78
timestamp 1688980957
transform 1 0 8280 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_90
timestamp 1688980957
transform 1 0 9384 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_98
timestamp 1688980957
transform 1 0 10120 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_109
timestamp 1688980957
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_285
timestamp 1688980957
transform 1 0 27324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_288
timestamp 1688980957
transform 1 0 27600 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_23
timestamp 1688980957
transform 1 0 3220 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1688980957
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_317
timestamp 1688980957
transform 1 0 30268 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_346
timestamp 1688980957
transform 1 0 32936 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_352
timestamp 1688980957
transform 1 0 33488 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_19
timestamp 1688980957
transform 1 0 2852 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_25
timestamp 1688980957
transform 1 0 3404 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_273
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_277
timestamp 1688980957
transform 1 0 26588 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_311
timestamp 1688980957
transform 1 0 29716 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_9
timestamp 1688980957
transform 1 0 1932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_38
timestamp 1688980957
transform 1 0 4600 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_44
timestamp 1688980957
transform 1 0 5152 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_69
timestamp 1688980957
transform 1 0 7452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_81
timestamp 1688980957
transform 1 0 8556 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_93
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_105
timestamp 1688980957
transform 1 0 10764 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_117
timestamp 1688980957
transform 1 0 11868 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_129
timestamp 1688980957
transform 1 0 12972 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_137
timestamp 1688980957
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1688980957
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_346
timestamp 1688980957
transform 1 0 32936 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_352
timestamp 1688980957
transform 1 0 33488 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_63
timestamp 1688980957
transform 1 0 6900 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_72
timestamp 1688980957
transform 1 0 7728 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_84
timestamp 1688980957
transform 1 0 8832 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_96
timestamp 1688980957
transform 1 0 9936 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_108
timestamp 1688980957
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_292
timestamp 1688980957
transform 1 0 27968 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_9
timestamp 1688980957
transform 1 0 1932 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_35
timestamp 1688980957
transform 1 0 4324 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_75
timestamp 1688980957
transform 1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_106
timestamp 1688980957
transform 1 0 10856 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_118
timestamp 1688980957
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_130
timestamp 1688980957
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_241
timestamp 1688980957
transform 1 0 23276 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_249
timestamp 1688980957
transform 1 0 24012 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_281
timestamp 1688980957
transform 1 0 26956 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_315
timestamp 1688980957
transform 1 0 30084 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_325
timestamp 1688980957
transform 1 0 31004 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_331
timestamp 1688980957
transform 1 0 31556 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_348
timestamp 1688980957
transform 1 0 33120 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_352
timestamp 1688980957
transform 1 0 33488 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_9
timestamp 1688980957
transform 1 0 1932 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_63
timestamp 1688980957
transform 1 0 6900 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_80
timestamp 1688980957
transform 1 0 8464 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_86
timestamp 1688980957
transform 1 0 9016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_103
timestamp 1688980957
transform 1 0 10580 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_131
timestamp 1688980957
transform 1 0 13156 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_135
timestamp 1688980957
transform 1 0 13524 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_151
timestamp 1688980957
transform 1 0 14996 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_155
timestamp 1688980957
transform 1 0 15364 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_166
timestamp 1688980957
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_191
timestamp 1688980957
transform 1 0 18676 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_195
timestamp 1688980957
transform 1 0 19044 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_207
timestamp 1688980957
transform 1 0 20148 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_215
timestamp 1688980957
transform 1 0 20884 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_229
timestamp 1688980957
transform 1 0 22172 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_233
timestamp 1688980957
transform 1 0 22540 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_243
timestamp 1688980957
transform 1 0 23460 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_266
timestamp 1688980957
transform 1 0 25576 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_277
timestamp 1688980957
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_287
timestamp 1688980957
transform 1 0 27508 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_313
timestamp 1688980957
transform 1 0 29900 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_23
timestamp 1688980957
transform 1 0 3220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_35
timestamp 1688980957
transform 1 0 4324 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_45
timestamp 1688980957
transform 1 0 5244 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_64
timestamp 1688980957
transform 1 0 6992 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_89
timestamp 1688980957
transform 1 0 9292 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_130
timestamp 1688980957
transform 1 0 13064 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_150
timestamp 1688980957
transform 1 0 14904 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_156
timestamp 1688980957
transform 1 0 15456 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_191
timestamp 1688980957
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_205
timestamp 1688980957
transform 1 0 19964 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_225
timestamp 1688980957
transform 1 0 21804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_234
timestamp 1688980957
transform 1 0 22632 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_275
timestamp 1688980957
transform 1 0 26404 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_349
timestamp 1688980957
transform 1 0 33212 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_31
timestamp 1688980957
transform 1 0 3956 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_61
timestamp 1688980957
transform 1 0 6716 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_100
timestamp 1688980957
transform 1 0 10304 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_147
timestamp 1688980957
transform 1 0 14628 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_215
timestamp 1688980957
transform 1 0 20884 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_244
timestamp 1688980957
transform 1 0 23552 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_306
timestamp 1688980957
transform 1 0 29256 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_312
timestamp 1688980957
transform 1 0 29808 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_346
timestamp 1688980957
transform 1 0 32936 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_352
timestamp 1688980957
transform 1 0 33488 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_19
timestamp 1688980957
transform 1 0 2852 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_51
timestamp 1688980957
transform 1 0 5796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_57
timestamp 1688980957
transform 1 0 6348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_67
timestamp 1688980957
transform 1 0 7268 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_92
timestamp 1688980957
transform 1 0 9568 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_96
timestamp 1688980957
transform 1 0 9936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_108
timestamp 1688980957
transform 1 0 11040 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_114
timestamp 1688980957
transform 1 0 11592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_161
timestamp 1688980957
transform 1 0 15916 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_169
timestamp 1688980957
transform 1 0 16652 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_179
timestamp 1688980957
transform 1 0 17572 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_187
timestamp 1688980957
transform 1 0 18308 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_203
timestamp 1688980957
transform 1 0 19780 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_213
timestamp 1688980957
transform 1 0 20700 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_217
timestamp 1688980957
transform 1 0 21068 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_229
timestamp 1688980957
transform 1 0 22172 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_249
timestamp 1688980957
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_264
timestamp 1688980957
transform 1 0 25392 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_268
timestamp 1688980957
transform 1 0 25760 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_280
timestamp 1688980957
transform 1 0 26864 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_284
timestamp 1688980957
transform 1 0 27232 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_296
timestamp 1688980957
transform 1 0 28336 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_300
timestamp 1688980957
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_325
timestamp 1688980957
transform 1 0 31004 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_329
timestamp 1688980957
transform 1 0 31372 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_349
timestamp 1688980957
transform 1 0 33212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_21
timestamp 1688980957
transform 1 0 3036 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_29
timestamp 1688980957
transform 1 0 3772 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_68
timestamp 1688980957
transform 1 0 7360 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_74
timestamp 1688980957
transform 1 0 7912 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_85
timestamp 1688980957
transform 1 0 8924 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_141
timestamp 1688980957
transform 1 0 14076 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_179
timestamp 1688980957
transform 1 0 17572 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_189
timestamp 1688980957
transform 1 0 18492 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_195
timestamp 1688980957
transform 1 0 19044 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_221
timestamp 1688980957
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_277
timestamp 1688980957
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_333
timestamp 1688980957
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5060 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold2 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 5244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold4
timestamp 1688980957
transform -1 0 2852 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 2852 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold6
timestamp 1688980957
transform -1 0 2852 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold8
timestamp 1688980957
transform -1 0 2852 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform 1 0 3956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold10
timestamp 1688980957
transform -1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold12
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold14
timestamp 1688980957
transform -1 0 2852 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 6624 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold16
timestamp 1688980957
transform 1 0 9384 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 2852 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold18
timestamp 1688980957
transform -1 0 2852 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 9936 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold20
timestamp 1688980957
transform 1 0 12512 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform 1 0 30544 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold22
timestamp 1688980957
transform -1 0 31648 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 11408 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold24
timestamp 1688980957
transform -1 0 11408 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold26
timestamp 1688980957
transform 1 0 15088 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 4048 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold28
timestamp 1688980957
transform 1 0 7360 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 14444 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold30
timestamp 1688980957
transform -1 0 13984 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 32016 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold32
timestamp 1688980957
transform 1 0 32108 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 18860 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold34
timestamp 1688980957
transform 1 0 17204 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 32016 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold36
timestamp 1688980957
transform 1 0 32108 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform 1 0 30176 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold38
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 32108 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold40
timestamp 1688980957
transform -1 0 32016 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 26588 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold42
timestamp 1688980957
transform -1 0 26312 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform 1 0 30544 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold44
timestamp 1688980957
transform -1 0 31648 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 12236 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold46
timestamp 1688980957
transform 1 0 9936 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 28428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold48
timestamp 1688980957
transform 1 0 29900 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 30912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold50
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 30912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold52
timestamp 1688980957
transform 1 0 32108 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 30912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold54
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 30544 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold56
timestamp 1688980957
transform 1 0 32108 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 25576 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold58
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 24748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold60
timestamp 1688980957
transform 1 0 26404 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform -1 0 13800 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold62
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform 1 0 30912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold64
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 28980 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold66
timestamp 1688980957
transform -1 0 32016 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 13064 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold68
timestamp 1688980957
transform -1 0 11408 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 30544 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold70
timestamp 1688980957
transform -1 0 32016 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 32108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold72
timestamp 1688980957
transform -1 0 32016 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform -1 0 15088 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold74
timestamp 1688980957
transform -1 0 16560 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 32108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold76
timestamp 1688980957
transform -1 0 32016 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 10212 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold78
timestamp 1688980957
transform -1 0 8464 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 21436 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold80
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 31280 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold82
timestamp 1688980957
transform -1 0 31648 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 30636 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold84
timestamp 1688980957
transform -1 0 32016 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform -1 0 17388 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold86
timestamp 1688980957
transform -1 0 16560 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 21712 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold88
timestamp 1688980957
transform 1 0 24380 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 31740 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold90
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform -1 0 29072 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold92
timestamp 1688980957
transform -1 0 29440 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 26864 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold94
timestamp 1688980957
transform -1 0 27968 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 31740 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold96
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 29440 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold98
timestamp 1688980957
transform -1 0 32108 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 29164 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold100
timestamp 1688980957
transform -1 0 29900 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform -1 0 26956 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold102
timestamp 1688980957
transform 1 0 29532 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 26496 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold104
timestamp 1688980957
transform 1 0 29072 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold106
timestamp 1688980957
transform 1 0 7820 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 19596 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold108
timestamp 1688980957
transform 1 0 17664 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform -1 0 7452 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold110
timestamp 1688980957
transform -1 0 4324 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 29072 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold112
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 32476 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold114
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 1472 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold116
timestamp 1688980957
transform 1 0 4324 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform -1 0 26588 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold118
timestamp 1688980957
transform -1 0 25852 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold120
timestamp 1688980957
transform -1 0 2852 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold122
timestamp 1688980957
transform -1 0 2852 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform 1 0 3220 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold124
timestamp 1688980957
transform -1 0 2852 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 29808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold126
timestamp 1688980957
transform -1 0 30544 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform 1 0 2852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold128
timestamp 1688980957
transform -1 0 2852 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 27600 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold130
timestamp 1688980957
transform -1 0 31648 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform 1 0 4324 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold132
timestamp 1688980957
transform -1 0 2852 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 26128 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold134
timestamp 1688980957
transform 1 0 30544 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold136
timestamp 1688980957
transform 1 0 2852 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform 1 0 4324 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold138
timestamp 1688980957
transform -1 0 2852 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform -1 0 8464 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold140
timestamp 1688980957
transform -1 0 6256 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold142
timestamp 1688980957
transform 1 0 2852 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold144
timestamp 1688980957
transform -1 0 2852 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 5428 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold146
timestamp 1688980957
transform -1 0 2852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold148
timestamp 1688980957
transform -1 0 29072 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold150
timestamp 1688980957
transform -1 0 2852 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform -1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold152
timestamp 1688980957
transform 1 0 4324 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform -1 0 9660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold154
timestamp 1688980957
transform -1 0 5796 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform -1 0 18308 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold156
timestamp 1688980957
transform 1 0 19228 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold158
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform -1 0 17480 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold160
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold162
timestamp 1688980957
transform 1 0 2852 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform 1 0 28704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold164
timestamp 1688980957
transform 1 0 30544 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 5520 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold166
timestamp 1688980957
transform -1 0 6256 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform -1 0 20424 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold168
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform 1 0 3220 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold170
timestamp 1688980957
transform -1 0 2852 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform -1 0 25116 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold172
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform -1 0 27692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_12  hold174
timestamp 1688980957
transform -1 0 32108 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  hold175 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  hold176
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform -1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform -1 0 3680 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 8004 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform 1 0 6992 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform 1 0 30912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform 1 0 30176 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform -1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform 1 0 30912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform 1 0 31280 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform -1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform -1 0 30544 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform 1 0 30912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform 1 0 16468 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform -1 0 17572 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform 1 0 27232 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform 1 0 27232 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform 1 0 24748 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform 1 0 28152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform -1 0 4692 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 3956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform -1 0 3680 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform -1 0 4508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform -1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform -1 0 9844 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform -1 0 4508 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform -1 0 3956 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform 1 0 2852 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform -1 0 3588 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 31648 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform 1 0 29808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform 1 0 10672 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform -1 0 11960 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 32016 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform 1 0 30912 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform -1 0 32016 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform 1 0 30912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform -1 0 5796 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform 1 0 25116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform 1 0 24748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform -1 0 30544 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform 1 0 25944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform 1 0 11776 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform -1 0 32016 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform 1 0 30912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform 1 0 2852 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform -1 0 5244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform 1 0 14352 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform 1 0 14352 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform 1 0 16100 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform -1 0 5244 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform -1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 31280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform 1 0 31280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 2484 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform -1 0 3680 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform 1 0 24104 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform 1 0 27232 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform 1 0 27968 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform -1 0 12604 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform -1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform 1 0 13156 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform -1 0 13800 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform 1 0 26680 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform -1 0 32016 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform -1 0 32108 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1688980957
transform -1 0 32108 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform 1 0 31280 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold261
timestamp 1688980957
transform -1 0 30636 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform 1 0 29808 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold263
timestamp 1688980957
transform 1 0 13984 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform 1 0 14720 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1688980957
transform -1 0 22632 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1688980957
transform -1 0 24012 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 1688980957
transform -1 0 32016 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1688980957
transform 1 0 31372 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1688980957
transform -1 0 25116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold270
timestamp 1688980957
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1688980957
transform -1 0 4508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold274
timestamp 1688980957
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform -1 0 4324 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 1688980957
transform -1 0 3680 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 1688980957
transform 1 0 12328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform -1 0 30636 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform -1 0 33580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1688980957
transform 1 0 6992 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1688980957
transform 1 0 6532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1688980957
transform -1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1688980957
transform -1 0 3588 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold286
timestamp 1688980957
transform -1 0 4508 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform 1 0 11408 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1688980957
transform -1 0 9936 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1688980957
transform 1 0 25760 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform 1 0 29072 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 1688980957
transform -1 0 10948 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform -1 0 10120 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform 1 0 9384 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1688980957
transform -1 0 9384 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform -1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold296
timestamp 1688980957
transform -1 0 5244 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1688980957
transform -1 0 18860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform -1 0 4692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform -1 0 4508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1688980957
transform 1 0 26680 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1688980957
transform 1 0 27968 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1688980957
transform 1 0 25852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform -1 0 28244 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1688980957
transform 1 0 25392 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1688980957
transform -1 0 29164 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1688980957
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1688980957
transform 1 0 28336 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform -1 0 33212 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform -1 0 3588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform -1 0 4508 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 1688980957
transform -1 0 29440 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform 1 0 28336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1688980957
transform -1 0 28704 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1688980957
transform 1 0 24748 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1688980957
transform -1 0 28152 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform 1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 1688980957
transform 1 0 22816 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1688980957
transform 1 0 23276 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1688980957
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1688980957
transform -1 0 3680 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1688980957
transform -1 0 5244 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform -1 0 3680 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 1688980957
transform -1 0 4508 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 1688980957
transform -1 0 7636 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1688980957
transform -1 0 11132 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold328
timestamp 1688980957
transform -1 0 7176 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1688980957
transform 1 0 27876 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 1688980957
transform 1 0 28980 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 1688980957
transform 1 0 5244 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1688980957
transform -1 0 4508 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold334
timestamp 1688980957
transform 1 0 16744 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold335
timestamp 1688980957
transform 1 0 19320 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1688980957
transform 1 0 19320 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold337
timestamp 1688980957
transform 1 0 5336 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1688980957
transform -1 0 9660 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1688980957
transform 1 0 22632 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1688980957
transform -1 0 25024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1688980957
transform -1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 1688980957
transform -1 0 4508 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1688980957
transform 1 0 15456 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold344
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1688980957
transform 1 0 19504 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold346
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1688980957
transform -1 0 4508 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1688980957
transform -1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1688980957
transform -1 0 11408 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1688980957
transform -1 0 15364 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold352
timestamp 1688980957
transform 1 0 23460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  output2 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2852 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output3
timestamp 1688980957
transform -1 0 5244 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output4
timestamp 1688980957
transform -1 0 3036 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output5
timestamp 1688980957
transform -1 0 7268 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output6
timestamp 1688980957
transform -1 0 8188 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output7
timestamp 1688980957
transform -1 0 8832 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output8
timestamp 1688980957
transform -1 0 11040 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output9
timestamp 1688980957
transform -1 0 12512 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output10
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output11
timestamp 1688980957
transform 1 0 15088 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output12
timestamp 1688980957
transform 1 0 16744 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output13
timestamp 1688980957
transform -1 0 5244 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output14
timestamp 1688980957
transform 1 0 19872 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output15
timestamp 1688980957
transform -1 0 23276 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output16
timestamp 1688980957
transform 1 0 26036 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output17
timestamp 1688980957
transform 1 0 24564 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output18
timestamp 1688980957
transform 1 0 27508 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output19
timestamp 1688980957
transform 1 0 28428 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output20
timestamp 1688980957
transform -1 0 32476 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output21
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output22
timestamp 1688980957
transform 1 0 27968 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output23
timestamp 1688980957
transform 1 0 30544 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output24
timestamp 1688980957
transform 1 0 17664 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output25
timestamp 1688980957
transform -1 0 23276 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output26
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output27
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output28
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output29
timestamp 1688980957
transform 1 0 27876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output30
timestamp 1688980957
transform -1 0 30360 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output31
timestamp 1688980957
transform 1 0 31648 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output32
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output33
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output34
timestamp 1688980957
transform 1 0 30544 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output35
timestamp 1688980957
transform 1 0 20240 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output36
timestamp 1688980957
transform 1 0 32752 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output37
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output38
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output39
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output40
timestamp 1688980957
transform 1 0 32108 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output41
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output42
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output43
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output44
timestamp 1688980957
transform 1 0 32108 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output45
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output46
timestamp 1688980957
transform 1 0 32108 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output47
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output48
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output49
timestamp 1688980957
transform 1 0 32108 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output50
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output51
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output52
timestamp 1688980957
transform 1 0 32108 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output53
timestamp 1688980957
transform 1 0 32108 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output54
timestamp 1688980957
transform -1 0 29900 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output55
timestamp 1688980957
transform 1 0 27968 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output56
timestamp 1688980957
transform 1 0 30176 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output57
timestamp 1688980957
transform 1 0 32108 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output58
timestamp 1688980957
transform -1 0 7360 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output59
timestamp 1688980957
transform -1 0 6256 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output60
timestamp 1688980957
transform -1 0 8832 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output61
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output62
timestamp 1688980957
transform -1 0 13156 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output63
timestamp 1688980957
transform -1 0 13156 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output64
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output65
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output66
timestamp 1688980957
transform -1 0 18308 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output67
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output68
timestamp 1688980957
transform -1 0 5888 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output69
timestamp 1688980957
transform -1 0 5060 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output70
timestamp 1688980957
transform -1 0 2852 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output71
timestamp 1688980957
transform -1 0 2852 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output72
timestamp 1688980957
transform -1 0 2852 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output73
timestamp 1688980957
transform -1 0 2852 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output74
timestamp 1688980957
transform -1 0 2852 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output75
timestamp 1688980957
transform -1 0 2852 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output76
timestamp 1688980957
transform -1 0 2852 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output77
timestamp 1688980957
transform -1 0 4324 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output78
timestamp 1688980957
transform -1 0 2852 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output79
timestamp 1688980957
transform -1 0 2852 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output80
timestamp 1688980957
transform -1 0 2852 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output81
timestamp 1688980957
transform -1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output82
timestamp 1688980957
transform -1 0 2852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output83
timestamp 1688980957
transform -1 0 2852 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output84
timestamp 1688980957
transform -1 0 2852 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output85
timestamp 1688980957
transform -1 0 2852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output86
timestamp 1688980957
transform -1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output87
timestamp 1688980957
transform -1 0 2852 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output88
timestamp 1688980957
transform -1 0 2852 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  output89
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 33856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 33856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 33856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 33856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 33856 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 33856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 33856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 33856 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 33856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 33856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 33856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 33856 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 33856 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 33856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 33856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 33856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 33856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 33856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 33856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 33856 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 33856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 33856 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 33856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 33856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 33856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 33856 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 33856 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 33856 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 33856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 33856 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 33856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 33856 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 33856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 33856 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 33856 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 33856 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 33856 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 33856 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 33856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 33856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 33856 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 33856 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 33856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 33856 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 33856 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 33856 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 33856 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 33856 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 33856 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 33856 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 33856 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 33856 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 33856 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 33856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 33856 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 3680 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 8832 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 13984 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 19136 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 24288 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 29440 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  unused_tie_97 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  unused_tie_98
timestamp 1688980957
transform -1 0 3128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  unused_tie_99
timestamp 1688980957
transform -1 0 4048 0 1 2176
box -38 -48 314 592
<< labels >>
flabel metal2 s 846 0 902 800 0 FreeSans 224 90 0 0 irq[0]
port 0 nsew signal tristate
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 irq[1]
port 1 nsew signal tristate
flabel metal2 s 3606 0 3662 800 0 FreeSans 224 90 0 0 irq[2]
port 2 nsew signal tristate
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 la_data_out[0]
port 3 nsew signal tristate
flabel metal2 s 2594 34200 2650 35000 0 FreeSans 224 90 0 0 la_data_out[10]
port 4 nsew signal tristate
flabel metal2 s 4158 34200 4214 35000 0 FreeSans 224 90 0 0 la_data_out[11]
port 5 nsew signal tristate
flabel metal2 s 5722 34200 5778 35000 0 FreeSans 224 90 0 0 la_data_out[12]
port 6 nsew signal tristate
flabel metal2 s 7286 34200 7342 35000 0 FreeSans 224 90 0 0 la_data_out[13]
port 7 nsew signal tristate
flabel metal2 s 8850 34200 8906 35000 0 FreeSans 224 90 0 0 la_data_out[14]
port 8 nsew signal tristate
flabel metal2 s 10414 34200 10470 35000 0 FreeSans 224 90 0 0 la_data_out[15]
port 9 nsew signal tristate
flabel metal2 s 11978 34200 12034 35000 0 FreeSans 224 90 0 0 la_data_out[16]
port 10 nsew signal tristate
flabel metal2 s 13542 34200 13598 35000 0 FreeSans 224 90 0 0 la_data_out[17]
port 11 nsew signal tristate
flabel metal2 s 15106 34200 15162 35000 0 FreeSans 224 90 0 0 la_data_out[18]
port 12 nsew signal tristate
flabel metal2 s 16670 34200 16726 35000 0 FreeSans 224 90 0 0 la_data_out[19]
port 13 nsew signal tristate
flabel metal2 s 1030 34200 1086 35000 0 FreeSans 224 90 0 0 la_data_out[1]
port 14 nsew signal tristate
flabel metal2 s 19798 34200 19854 35000 0 FreeSans 224 90 0 0 la_data_out[20]
port 15 nsew signal tristate
flabel metal2 s 21362 34200 21418 35000 0 FreeSans 224 90 0 0 la_data_out[21]
port 16 nsew signal tristate
flabel metal2 s 22926 34200 22982 35000 0 FreeSans 224 90 0 0 la_data_out[22]
port 17 nsew signal tristate
flabel metal2 s 24490 34200 24546 35000 0 FreeSans 224 90 0 0 la_data_out[23]
port 18 nsew signal tristate
flabel metal2 s 26054 34200 26110 35000 0 FreeSans 224 90 0 0 la_data_out[24]
port 19 nsew signal tristate
flabel metal2 s 27618 34200 27674 35000 0 FreeSans 224 90 0 0 la_data_out[25]
port 20 nsew signal tristate
flabel metal2 s 29182 34200 29238 35000 0 FreeSans 224 90 0 0 la_data_out[26]
port 21 nsew signal tristate
flabel metal2 s 30746 34200 30802 35000 0 FreeSans 224 90 0 0 la_data_out[27]
port 22 nsew signal tristate
flabel metal2 s 32310 34200 32366 35000 0 FreeSans 224 90 0 0 la_data_out[28]
port 23 nsew signal tristate
flabel metal2 s 33874 34200 33930 35000 0 FreeSans 224 90 0 0 la_data_out[29]
port 24 nsew signal tristate
flabel metal2 s 18234 34200 18290 35000 0 FreeSans 224 90 0 0 la_data_out[2]
port 25 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 26 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 27 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 28 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 29 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 30 nsew signal tristate
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 31 nsew signal tristate
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 32 nsew signal tristate
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 33 nsew signal tristate
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 34 nsew signal tristate
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 35 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 36 nsew signal tristate
flabel metal3 s 34200 5720 35000 5840 0 FreeSans 480 0 0 0 la_data_out[40]
port 37 nsew signal tristate
flabel metal3 s 34200 7080 35000 7200 0 FreeSans 480 0 0 0 la_data_out[41]
port 38 nsew signal tristate
flabel metal3 s 34200 8440 35000 8560 0 FreeSans 480 0 0 0 la_data_out[42]
port 39 nsew signal tristate
flabel metal3 s 34200 9800 35000 9920 0 FreeSans 480 0 0 0 la_data_out[43]
port 40 nsew signal tristate
flabel metal3 s 34200 11160 35000 11280 0 FreeSans 480 0 0 0 la_data_out[44]
port 41 nsew signal tristate
flabel metal3 s 34200 12520 35000 12640 0 FreeSans 480 0 0 0 la_data_out[45]
port 42 nsew signal tristate
flabel metal3 s 34200 13880 35000 14000 0 FreeSans 480 0 0 0 la_data_out[46]
port 43 nsew signal tristate
flabel metal3 s 34200 15240 35000 15360 0 FreeSans 480 0 0 0 la_data_out[47]
port 44 nsew signal tristate
flabel metal3 s 34200 16600 35000 16720 0 FreeSans 480 0 0 0 la_data_out[48]
port 45 nsew signal tristate
flabel metal3 s 34200 17960 35000 18080 0 FreeSans 480 0 0 0 la_data_out[49]
port 46 nsew signal tristate
flabel metal3 s 34200 4360 35000 4480 0 FreeSans 480 0 0 0 la_data_out[4]
port 47 nsew signal tristate
flabel metal3 s 34200 20680 35000 20800 0 FreeSans 480 0 0 0 la_data_out[50]
port 48 nsew signal tristate
flabel metal3 s 34200 22040 35000 22160 0 FreeSans 480 0 0 0 la_data_out[51]
port 49 nsew signal tristate
flabel metal3 s 34200 23400 35000 23520 0 FreeSans 480 0 0 0 la_data_out[52]
port 50 nsew signal tristate
flabel metal3 s 34200 24760 35000 24880 0 FreeSans 480 0 0 0 la_data_out[53]
port 51 nsew signal tristate
flabel metal3 s 34200 26120 35000 26240 0 FreeSans 480 0 0 0 la_data_out[54]
port 52 nsew signal tristate
flabel metal3 s 34200 27480 35000 27600 0 FreeSans 480 0 0 0 la_data_out[55]
port 53 nsew signal tristate
flabel metal3 s 34200 28840 35000 28960 0 FreeSans 480 0 0 0 la_data_out[56]
port 54 nsew signal tristate
flabel metal3 s 34200 30200 35000 30320 0 FreeSans 480 0 0 0 la_data_out[57]
port 55 nsew signal tristate
flabel metal3 s 34200 31560 35000 31680 0 FreeSans 480 0 0 0 la_data_out[58]
port 56 nsew signal tristate
flabel metal3 s 34200 32920 35000 33040 0 FreeSans 480 0 0 0 la_data_out[59]
port 57 nsew signal tristate
flabel metal3 s 34200 19320 35000 19440 0 FreeSans 480 0 0 0 la_data_out[5]
port 58 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 59 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 60 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 61 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 62 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 63 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 64 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 65 nsew signal tristate
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 66 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 67 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 68 nsew signal tristate
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 69 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 la_data_out[70]
port 70 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 la_data_out[71]
port 71 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 la_data_out[72]
port 72 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 la_data_out[73]
port 73 nsew signal tristate
flabel metal3 s 0 22040 800 22160 0 FreeSans 480 0 0 0 la_data_out[74]
port 74 nsew signal tristate
flabel metal3 s 0 23400 800 23520 0 FreeSans 480 0 0 0 la_data_out[75]
port 75 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 la_data_out[76]
port 76 nsew signal tristate
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 la_data_out[77]
port 77 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 la_data_out[78]
port 78 nsew signal tristate
flabel metal3 s 0 28840 800 28960 0 FreeSans 480 0 0 0 la_data_out[79]
port 79 nsew signal tristate
flabel metal3 s 0 15240 800 15360 0 FreeSans 480 0 0 0 la_data_out[7]
port 80 nsew signal tristate
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 la_data_out[80]
port 81 nsew signal tristate
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 la_data_out[81]
port 82 nsew signal tristate
flabel metal3 s 0 7080 800 7200 0 FreeSans 480 0 0 0 la_data_out[82]
port 83 nsew signal tristate
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 la_data_out[83]
port 84 nsew signal tristate
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 la_data_out[84]
port 85 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 la_data_out[85]
port 86 nsew signal tristate
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 la_data_out[86]
port 87 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 la_data_out[87]
port 88 nsew signal tristate
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 la_data_out[8]
port 89 nsew signal tristate
flabel metal3 s 0 31560 800 31680 0 FreeSans 480 0 0 0 la_data_out[9]
port 90 nsew signal tristate
flabel metal4 s 5038 2128 5358 32688 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 13226 2128 13546 32688 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 21414 2128 21734 32688 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 29602 2128 29922 32688 0 FreeSans 1920 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal4 s 9132 2128 9452 32688 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew ground bidirectional
flabel metal4 s 17320 2128 17640 32688 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew ground bidirectional
flabel metal4 s 25508 2128 25828 32688 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew ground bidirectional
flabel metal4 s 33696 2128 34016 32688 0 FreeSans 1920 90 0 0 vssd1
port 92 nsew ground bidirectional
flabel metal3 s 34200 1640 35000 1760 0 FreeSans 480 0 0 0 wb_clk_i
port 93 nsew signal input
flabel metal3 s 34200 3000 35000 3120 0 FreeSans 480 0 0 0 wb_rst_i
port 94 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 35000 35000
<< end >>
