// This is the unpowered netlist.
module execution_unit (busy,
    dest_pred_val,
    int_return,
    is_load,
    is_store,
    pred_val,
    rst,
    sign_extend,
    take_branch,
    wb_clk_i,
    curr_PC,
    dest_idx,
    dest_mask,
    dest_pred,
    dest_val,
    instruction,
    loadstore_address,
    loadstore_size,
    new_PC,
    pred_idx,
    reg1_idx,
    reg1_val,
    reg2_idx,
    reg2_val);
 output busy;
 output dest_pred_val;
 output int_return;
 output is_load;
 output is_store;
 input pred_val;
 input rst;
 output sign_extend;
 output take_branch;
 input wb_clk_i;
 input [27:0] curr_PC;
 output [5:0] dest_idx;
 output [1:0] dest_mask;
 output [2:0] dest_pred;
 output [31:0] dest_val;
 input [41:0] instruction;
 output [31:0] loadstore_address;
 output [1:0] loadstore_size;
 output [27:0] new_PC;
 output [2:0] pred_idx;
 output [5:0] reg1_idx;
 input [31:0] reg1_val;
 output [5:0] reg2_idx;
 input [31:0] reg2_val;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire busy_l;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire div_complete;
 wire \div_counter[0] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_res[0] ;
 wire \div_res[10] ;
 wire \div_res[11] ;
 wire \div_res[12] ;
 wire \div_res[13] ;
 wire \div_res[14] ;
 wire \div_res[15] ;
 wire \div_res[16] ;
 wire \div_res[17] ;
 wire \div_res[18] ;
 wire \div_res[19] ;
 wire \div_res[1] ;
 wire \div_res[20] ;
 wire \div_res[21] ;
 wire \div_res[22] ;
 wire \div_res[23] ;
 wire \div_res[24] ;
 wire \div_res[25] ;
 wire \div_res[26] ;
 wire \div_res[27] ;
 wire \div_res[28] ;
 wire \div_res[29] ;
 wire \div_res[2] ;
 wire \div_res[30] ;
 wire \div_res[31] ;
 wire \div_res[3] ;
 wire \div_res[4] ;
 wire \div_res[5] ;
 wire \div_res[6] ;
 wire \div_res[7] ;
 wire \div_res[8] ;
 wire \div_res[9] ;
 wire \div_shifter[0] ;
 wire \div_shifter[10] ;
 wire \div_shifter[11] ;
 wire \div_shifter[12] ;
 wire \div_shifter[13] ;
 wire \div_shifter[14] ;
 wire \div_shifter[15] ;
 wire \div_shifter[16] ;
 wire \div_shifter[17] ;
 wire \div_shifter[18] ;
 wire \div_shifter[19] ;
 wire \div_shifter[1] ;
 wire \div_shifter[20] ;
 wire \div_shifter[21] ;
 wire \div_shifter[22] ;
 wire \div_shifter[23] ;
 wire \div_shifter[24] ;
 wire \div_shifter[25] ;
 wire \div_shifter[26] ;
 wire \div_shifter[27] ;
 wire \div_shifter[28] ;
 wire \div_shifter[29] ;
 wire \div_shifter[2] ;
 wire \div_shifter[30] ;
 wire \div_shifter[31] ;
 wire \div_shifter[32] ;
 wire \div_shifter[33] ;
 wire \div_shifter[34] ;
 wire \div_shifter[35] ;
 wire \div_shifter[36] ;
 wire \div_shifter[37] ;
 wire \div_shifter[38] ;
 wire \div_shifter[39] ;
 wire \div_shifter[3] ;
 wire \div_shifter[40] ;
 wire \div_shifter[41] ;
 wire \div_shifter[42] ;
 wire \div_shifter[43] ;
 wire \div_shifter[44] ;
 wire \div_shifter[45] ;
 wire \div_shifter[46] ;
 wire \div_shifter[47] ;
 wire \div_shifter[48] ;
 wire \div_shifter[49] ;
 wire \div_shifter[4] ;
 wire \div_shifter[50] ;
 wire \div_shifter[51] ;
 wire \div_shifter[52] ;
 wire \div_shifter[53] ;
 wire \div_shifter[54] ;
 wire \div_shifter[55] ;
 wire \div_shifter[56] ;
 wire \div_shifter[57] ;
 wire \div_shifter[58] ;
 wire \div_shifter[59] ;
 wire \div_shifter[5] ;
 wire \div_shifter[60] ;
 wire \div_shifter[61] ;
 wire \div_shifter[62] ;
 wire \div_shifter[63] ;
 wire \div_shifter[6] ;
 wire \div_shifter[7] ;
 wire \div_shifter[8] ;
 wire \div_shifter[9] ;
 wire divi1_sign;
 wire \divi2_l[0] ;
 wire \divi2_l[10] ;
 wire \divi2_l[11] ;
 wire \divi2_l[12] ;
 wire \divi2_l[13] ;
 wire \divi2_l[14] ;
 wire \divi2_l[15] ;
 wire \divi2_l[16] ;
 wire \divi2_l[17] ;
 wire \divi2_l[18] ;
 wire \divi2_l[19] ;
 wire \divi2_l[1] ;
 wire \divi2_l[20] ;
 wire \divi2_l[21] ;
 wire \divi2_l[22] ;
 wire \divi2_l[23] ;
 wire \divi2_l[24] ;
 wire \divi2_l[25] ;
 wire \divi2_l[26] ;
 wire \divi2_l[27] ;
 wire \divi2_l[28] ;
 wire \divi2_l[29] ;
 wire \divi2_l[2] ;
 wire \divi2_l[30] ;
 wire \divi2_l[31] ;
 wire \divi2_l[3] ;
 wire \divi2_l[4] ;
 wire \divi2_l[5] ;
 wire \divi2_l[6] ;
 wire \divi2_l[7] ;
 wire \divi2_l[8] ;
 wire \divi2_l[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00468_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(instruction[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(instruction[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(instruction[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(instruction[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(instruction[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(instruction[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(instruction[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(instruction[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(instruction[37]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(instruction[38]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(instruction[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(instruction[40]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(reg1_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(reg1_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(reg1_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(reg1_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(reg1_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(reg1_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(reg1_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(reg1_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_03086_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(reg1_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(reg1_val[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(reg1_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(reg1_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(reg1_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(reg1_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(reg1_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_03378_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(reg1_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(reg2_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(reg2_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(reg2_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(reg2_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(reg2_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(reg2_val[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(reg2_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_06537_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(reg2_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(reg2_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(reg2_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(reg2_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(reg2_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(reg2_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(reg2_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(reg2_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(reg2_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(reg2_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(reg2_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(reg2_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(reg2_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(reg2_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(reg2_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(rst));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(instruction[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_03663_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_04701_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(reg1_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(reg1_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(reg1_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(reg1_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(reg1_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(reg1_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(reg1_val[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(instruction[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(reg1_val[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(reg1_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(reg1_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(reg1_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(reg1_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(reg1_val[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(reg1_val[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(instruction[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__06748__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__06749__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06750__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06770__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__A2 (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__B (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__B (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__B (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06803__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__B (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06806__A (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__B (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__B (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__A (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__B (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__B (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__B (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__B (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__B1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__B (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06841__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__B (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__B (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__A2_N (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06854__B (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06855__B (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06857__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__B (.DIODE(_05634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__B (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__B (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__B (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__B (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__A2_N (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__B (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__B (.DIODE(_05807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06878__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__B (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__B (.DIODE(_05874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__B (.DIODE(_05874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__A_N (.DIODE(_05874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__B (.DIODE(_05921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__A2_N (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__B (.DIODE(_06004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A2_N (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__B (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06903__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__B (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__B (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__B1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__A2_N (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A2 (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A3 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__A_N (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__B (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__B (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__B (.DIODE(_04764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A3 (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__C (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__B (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__C (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__A3 (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A3 (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__A3 (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A3 (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A3 (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A_N (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__B (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__B (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A3 (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A3 (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__A3 (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__A_N (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__B (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__B (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__B (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A3 (.DIODE(_05634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__A (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__B (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__B (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__B (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__C1 (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__D1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__C_N (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A3 (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A3 (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__A3 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A3 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__B (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07011__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__A3 (.DIODE(_05921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A3 (.DIODE(_05921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__B (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__D1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__B (.DIODE(_06567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__B (.DIODE(_06567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__B (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__A2 (.DIODE(_06567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__B (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__C (.DIODE(_06567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__A3 (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__A3 (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__B2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__B (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__B (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__B (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__S (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__A1 (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__D (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__B (.DIODE(_06661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__B (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__B (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__B (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__B (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__B (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__B (.DIODE(_06664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07131__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__S (.DIODE(_04652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__C (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__A2 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__B1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__A2 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__C (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A1 (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A2 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B1 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07165__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__S (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__A (.DIODE(_06694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A (.DIODE(_06694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__A (.DIODE(_06694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__B (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__B (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__B (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__C (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__D (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A_N (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__B_N (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__D (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__A (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__C (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__A (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__A (.DIODE(_05874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__C (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A1 (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A2 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__C1 (.DIODE(_05807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__C1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A1 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__B1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A2 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__A (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__A1 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A1 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A2 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A2 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__A (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07232__A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__S (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__B (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__A2 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__A0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__S (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__B1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__B1 (.DIODE(_05874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__A (.DIODE(_05874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A2 (.DIODE(_06719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B1 (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__S (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__B (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__A (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A1 (.DIODE(_00220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__B1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__C (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__C (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__C (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__B (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__C (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__B (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__C (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07349__C (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__S (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__C_N (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__B1 (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07374__C (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__A (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__C (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__D (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A3 (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A4 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__C (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__A3 (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__S (.DIODE(_00302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07398__B (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07398__C (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__B1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07403__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__C1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__S (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A2 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A3 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__B1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__A (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__C (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A3 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__B (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A2 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__S (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07451__A (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__A (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__S (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__S (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__A1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__B (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__S (.DIODE(_00274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__A2 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__A3 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__A (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A2 (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__S (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A2 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__B (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__B1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__B (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__A (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A1 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A2 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__B1 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__B1 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__A (.DIODE(_06529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A1 (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__S (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__C (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B1 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B2 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__A1 (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__B (.DIODE(_06703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__A (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__B (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__B (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__B1 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A2 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__B2 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A1 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__B2 (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__B2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__A2 (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__B2 (.DIODE(_00477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__C (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__D (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__B (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A1 (.DIODE(_00371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A1 (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__B2 (.DIODE(_00477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A2 (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__B2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07692__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__B1 (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__B2 (.DIODE(_00327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B2 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__A1 (.DIODE(_00220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__B2 (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__B1 (.DIODE(_00477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B1 (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A2 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B2 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__B1 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__B (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__S (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A2 (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__B2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B1 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__C1 (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__C1 (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__B (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__C (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__B2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A2 (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B1 (.DIODE(_00477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__A1 (.DIODE(_00220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__A2 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__B2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__B1 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__A1 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__A2 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__B1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__B2 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__A2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__B2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__A1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A2 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__B1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__B2 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__A (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__B (.DIODE(_00991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__B2 (.DIODE(_00326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A1 (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A (.DIODE(_00991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__B (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A1 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A2 (.DIODE(_00220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__B2 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A1 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A2 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__B1 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__B2 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A0 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A2 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B1 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B2 (.DIODE(_00372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A1 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__B1 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__A1 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__A2 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__B2 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A1 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__A (.DIODE(_06694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__B1 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__A (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A1 (.DIODE(_00320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08264__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08269__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__B1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__B (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__B (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A1 (.DIODE(_01190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A1 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A2 (.DIODE(_00220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__B2 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A2 (.DIODE(_00372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__A1 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__A2 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__B1 (.DIODE(_00476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__B2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__B2 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__A2 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A2 (.DIODE(_00220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__B2 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A1 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__B1 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__B2 (.DIODE(_00476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__B (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__A2 (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__B2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A2 (.DIODE(_00372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08432__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A2 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A1 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B2 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08490__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08491__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__B1 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__B2 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08527__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__B2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08537__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A2 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__B1 (.DIODE(_00476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A1 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__B1 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__B (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__B1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__B2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__B1 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__B1 (.DIODE(_00476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08624__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08626__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08626__A2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08626__B1 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08626__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A1 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A2 (.DIODE(_00372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__B2 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A2 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__B2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08639__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08640__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A1 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A2 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__B2 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__B1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08666__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08668__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08676__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08680__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08680__A2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08680__B1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08680__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08682__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__A1 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__A2 (.DIODE(_00372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__B2 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08709__B2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__B1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08745__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08746__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__A2 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08748__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__B2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A2 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__B2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08768__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08772__B2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08778__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08778__B (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__B1_N (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08794__B2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__A2 (.DIODE(_00372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08796__B2 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08800__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08800__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08800__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08800__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08801__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__B2 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A2 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08826__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08832__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__08834__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__B (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__A2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__B1 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__B2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__B (.DIODE(_01754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__B2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__A1 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__B1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__B2 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__A1 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__B (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__A1 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__A2 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__B2 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__B1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08904__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__A2 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__B1 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__B2 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__A2 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08922__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__B2 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__08924__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__08932__B (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__B (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08934__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A2 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__B1 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__B2 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08940__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__B1 (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__B2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A2 (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__B2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__A1_N (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__B1 (.DIODE(_00320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__B2 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__09007__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A1 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__B1 (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09107__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__B2 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A1 (.DIODE(_00220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A2 (.DIODE(_00461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__B1 (.DIODE(_00465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__B2 (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__09137__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A1 (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__B1 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__B2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__09141__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__A (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__A2 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09147__B2 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__B (.DIODE(_02071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__B (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__B1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__09159__B1 (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09161__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09163__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09171__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A2 (.DIODE(_00371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__A1 (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09216__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A1 (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__B2 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09234__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09236__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__A1 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09244__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A2 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__B1 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__A (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09254__B (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__09258__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__B1 (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__B1 (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__C1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__D1 (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__B2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09274__A (.DIODE(_02191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A (.DIODE(_02191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__09282__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A1 (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__B2 (.DIODE(_00477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__A1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09334__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__B2 (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09351__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09355__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09361__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09363__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A2 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A2 (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A3 (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A1 (.DIODE(_00138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09385__A_N (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__A1 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A2 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A2 (.DIODE(_00371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__B (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__B (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__D_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09436__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__A0 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__A1 (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A1 (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__C1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__C1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09468__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__A0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09484__S (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__S (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__S (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__S (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__C1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__C1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__A_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A_N (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__D_N (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A1 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__B1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__A1 (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__B1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__A1_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__A2_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__B1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__B1 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__B (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__A (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__B1 (.DIODE(_00477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A1 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A1 (.DIODE(_00158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__B2 (.DIODE(_00159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__B (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__C (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__B1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__09590__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09618__B2 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__B1 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__B (.DIODE(_02568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09652__B2 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09658__A (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__C1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__S (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09674__S (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__S (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__S (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__09686__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09694__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__C1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__09702__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09704__B1 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__B (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A3 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A2_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__A1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09712__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09718__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09728__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__B2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09730__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__B1 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A (.DIODE(_00327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A1 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__B2 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A2 (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A3 (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A1 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__A2 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__B2 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__A3 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A2 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__B2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09792__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__B2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A2 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__B1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__A (.DIODE(_02642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__B (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__A (.DIODE(_02642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__B (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__A2 (.DIODE(_02344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__B1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__B2 (.DIODE(_02568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A2 (.DIODE(_02568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__09834__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A2 (.DIODE(_02776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__B1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__09865__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__B1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09871__C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__B2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__C1 (.DIODE(_02789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A1 (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__B2 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A2 (.DIODE(_00371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__A2 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__B1 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09891__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A2 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__B1 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A1 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__B2 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09927__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09928__B (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__B (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09930__B1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09931__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A1 (.DIODE(_06702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__B2 (.DIODE(_06726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A1 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__B2 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A2 (.DIODE(_02568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__B1 (.DIODE(_02642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__B2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09988__A1 (.DIODE(_02642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09988__A2 (.DIODE(_02740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__B1 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A3 (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__S (.DIODE(_06569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__S (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__A2 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__C1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__A2 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__C1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10029__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__A2_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__C1 (.DIODE(_02951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10038__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10039__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__B2 (.DIODE(_02957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10044__B (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__A2 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__B1 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10075__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__A2 (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__A3 (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10077__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__B2 (.DIODE(_00230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10087__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__10095__A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__B2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10119__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__A (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__D (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__A3 (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__B1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__B1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__S (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__S (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__A2_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__C1 (.DIODE(_03105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10191__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__B2 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10197__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__S (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__A2 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__B1 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__B1 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__B (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__A1_N (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__A2_N (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__B1 (.DIODE(_00797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__B2 (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__B2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__A2 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__B1 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__B1 (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10266__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__A1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__A (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__B (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__C (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__D (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__B1_N (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__A (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__A2 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__B1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__A2 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10309__B1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__S (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A2_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B1 (.DIODE(_03241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__B2 (.DIODE(_03242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__A1 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__B2 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10343__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__B (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__C1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__B1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A2 (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__A3 (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__A2 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__A1 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__B1 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A1 (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10388__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A2 (.DIODE(_00463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10401__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A1 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A2 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__B1 (.DIODE(_00446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__B2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__B (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__C (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__D (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__C1 (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__D1 (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__B1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__C1 (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__S (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__S (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10464__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__A2_N (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__B2 (.DIODE(_03379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__A2 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__B2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A1 (.DIODE(_00230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__A (.DIODE(_00274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A1 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__B1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__B (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__A2 (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__B1 (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A (.DIODE(_00302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__B1 (.DIODE(_00463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A1_N (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A2_N (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__B1 (.DIODE(_00797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__B (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__C (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__B1_N (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__A_N (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__B1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__B (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__A (.DIODE(_02902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__B (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__C (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__D (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__A1 (.DIODE(_03215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__B1 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A2 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__B1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A2 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__A1 (.DIODE(_06553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__S (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__A1 (.DIODE(_06523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__A2 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__B1_N (.DIODE(_03522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10617__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__A (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__B (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__B1 (.DIODE(_03540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__A (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__B (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__C (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__D (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__A1 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A1 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__B2 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__A1 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A2 (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__A3 (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__B (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__C (.DIODE(_02908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__A (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10727__B (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__B1 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__B (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__B (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__S (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__B (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__B1 (.DIODE(_03665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10755__B2 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10757__A1 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10758__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__10760__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__A (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__A (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__B (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__C (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10788__B1 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__B1 (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A1 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__B2 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__A1 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10802__B2 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__B1 (.DIODE(_00463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10810__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__A1 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__A (.DIODE(_00273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__A (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__B (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__A1 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__B1 (.DIODE(_03765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__A (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__B (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__C (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__D (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A (.DIODE(_03764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__B1 (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__C (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__B (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__C1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__C1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10884__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__A (.DIODE(_06509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__B (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10890__A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__10890__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__B1 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10893__D (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__B (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__A2 (.DIODE(_00463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__B1 (.DIODE(_00468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__A (.DIODE(_00302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__A (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__A1 (.DIODE(_00446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__B2 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__A1 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10912__B2 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A (.DIODE(_00273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A1 (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10921__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__B1 (.DIODE(_03845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__C (.DIODE(_03845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__B2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__B2 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__B (.DIODE(_03764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A1 (.DIODE(_03540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__B1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__A (.DIODE(_03346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__B (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__C (.DIODE(_03635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__D (.DIODE(_03764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__B (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__B1 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__A3 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__B1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__C1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__B1 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11014__C (.DIODE(_03923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__B2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11023__A2 (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__A (.DIODE(_03845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__A (.DIODE(_03845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__B2 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11032__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A1 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A1 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__B2 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A1_N (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A2_N (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__B1 (.DIODE(_00797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__11046__A (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11047__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__11047__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11052__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__B2 (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__A2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__B1 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11075__A_N (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__11076__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A (.DIODE(_03764_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__B (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__A1 (.DIODE(_03765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11110__B1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11112__B1 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__B (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__A2 (.DIODE(_04023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11116__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__B2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__B2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__A2 (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__B2 (.DIODE(_04046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__C1 (.DIODE(_04032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__B2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11149__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__B1_N (.DIODE(_03894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__A (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__C_N (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A1 (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__A2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A1 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__B2 (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B2 (.DIODE(_00230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A2 (.DIODE(_00513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A3 (.DIODE(_00515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A1 (.DIODE(_00446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__B2 (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__B1 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__C1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A1 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A (.DIODE(_03887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__B (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A1 (.DIODE(_03888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__B1 (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__A (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A2 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__B1 (.DIODE(_04137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__B (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__C (.DIODE(_04137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__A1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__B1 (.DIODE(_04165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__B (.DIODE(_04137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__A1_N (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__A2_N (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__B1 (.DIODE(_00797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__B2 (.DIODE(_00468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__A1 (.DIODE(_00230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__B2 (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11277__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__B (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__B1 (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__A (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__B1 (.DIODE(_00431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A (.DIODE(_00274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__B1 (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11304__B2 (.DIODE(_00446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__A2 (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__B (.DIODE(_04066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__A (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__B (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__A1 (.DIODE(_04018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__A (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__C (.DIODE(_04254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11349__B1 (.DIODE(_04254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__B1 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11357__B1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__C (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__B1 (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__C1 (.DIODE(_04282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__B2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__A2 (.DIODE(_04254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__A (.DIODE(_00274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__B2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__A1 (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__B1 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__B (.DIODE(_04317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11420__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__A (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__A1 (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A1 (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A (.DIODE(_04362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__B (.DIODE(_04362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__A2 (.DIODE(_04362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11479__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A1 (.DIODE(_00433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__B1 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__C1 (.DIODE(_04387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__A1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__B2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11490__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11491__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__A2 (.DIODE(_04254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__A1 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__A1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__A2 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__B1 (.DIODE(_02176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__A2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__B1 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11512__A (.DIODE(_00273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__A (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A_N (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__B (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__B1 (.DIODE(_04464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__B (.DIODE(_04471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__B (.DIODE(_04471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__11585__B (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__B1 (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__11593__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11594__A1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11595__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__B1 (.DIODE(_06165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__B2 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__A (.DIODE(_04137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__B (.DIODE(_04254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__C_N (.DIODE(_04362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__D_N (.DIODE(_04471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__B2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__B1 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11612__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11614__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11614__B1 (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A1 (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A3 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11620__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__A1 (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__B2 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11624__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__B2 (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__11634__A1 (.DIODE(_00381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__A2 (.DIODE(_02080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A1 (.DIODE(_00467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__A2 (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__B1 (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__B1 (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A3 (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__C1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__B1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__B (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__11689__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11693__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__11695__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__C (.DIODE(_04614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__B1 (.DIODE(_04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__B2 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11699__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11701__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__11703__A2 (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11703__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A2 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__B1 (.DIODE(_02176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__A2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__B1 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__A (.DIODE(_00359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11709__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__A1 (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__B2 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A1 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__B2 (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11731__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__B (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A1 (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A1 (.DIODE(_04464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__A2 (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__B1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A2 (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__11783__A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__C1 (.DIODE(_04710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__A1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__B2 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__B1 (.DIODE(_04701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__B2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__A (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__B (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__B (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11801__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11801__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__B (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__A (.DIODE(_04728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__A (.DIODE(_04728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__B1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__B2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A1 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__B2 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__B2 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__A (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A1 (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__B2 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__A1 (.DIODE(_03893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11862__B (.DIODE(_04792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A2 (.DIODE(_04792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__11870__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__C1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__A2_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__B2 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__A1_N (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__A1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11891__C1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__D (.DIODE(_04792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11903__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__A (.DIODE(_00274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__A2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__B1 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11911__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__A_N (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11917__B2 (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11918__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__A (.DIODE(_04728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__A (.DIODE(_04728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__A (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__B1 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11954__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__11954__C (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__11960__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__11962__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__11968__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__11974__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__A2_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A2_N (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__A3 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__A1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__A1 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__B1 (.DIODE(_04924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__A1 (.DIODE(_05874_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__B (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11992__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11992__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__B2 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__12003__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A1 (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__B2 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__A1 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__B1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__B2 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__B1 (.DIODE(_04986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__A3 (.DIODE(_04986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__S (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__A1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12056__B (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__B1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A1 (.DIODE(_05731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__A2 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__C1 (.DIODE(_05013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12066__A1 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__B2 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A2 (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A3 (.DIODE(_04986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__A1 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__B2 (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__A2 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__B1 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__A (.DIODE(_00274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__B (.DIODE(_05082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__B (.DIODE(_05082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__C1 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__S (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__B1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__C1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__A2 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12154__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12154__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12158__A1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__A (.DIODE(_04590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__B (.DIODE(_04693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__C (.DIODE(_04792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12164__A (.DIODE(_04891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12164__B (.DIODE(_04986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12164__C (.DIODE(_05082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__B2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12168__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__A1 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__B2 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12170__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__A2 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__B1 (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__A (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12178__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__A1 (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12184__B2 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__B1 (.DIODE(_05172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__A3 (.DIODE(_05172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__S (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__C (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__B1 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__B2 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A2 (.DIODE(_05172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__A2 (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__12249__A (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__A2 (.DIODE(_00517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__B1 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__A1 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12264__B2 (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__A1 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__B2 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__B (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__A2 (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__C1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__B1 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A1 (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__A2 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__A1 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__B2 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__A (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__A1 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__B2 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12338__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__A1 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__B2 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12340__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A2 (.DIODE(_00811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__12342__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__C (.DIODE(_05172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__D (.DIODE(_05264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__B1 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12381__S (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__12389__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12391__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12395__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__A2 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__A3 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__12403__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__B1 (.DIODE(_05356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__A1 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__B2 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__A (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12417__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__A1 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__B1 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__B1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__B1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__S (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__B1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__C1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12469__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__B1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__12473__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__C (.DIODE(_05440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__B1 (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12479__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__A2 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__B1 (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12483__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__A1 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12495__B2 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__A (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__B (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__S (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__C1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__B1 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12526__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12526__C1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__C (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A2_N (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__B2 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__B1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__12538__A2 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A1 (.DIODE(_05507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12540__A2 (.DIODE(_05508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A1 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12544__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__A1 (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A1 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__B2 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__A (.DIODE(_00302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A (.DIODE(_00302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A2 (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12554__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__B1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__B (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__C (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__B1 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12597__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__C (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12599__B1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__C1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__A1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12605__A1 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A1 (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__B2 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12610__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__A (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12614__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__A1 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12618__B2 (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12636__B1 (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__B1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12643__C1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__C1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__C1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12655__C1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__C (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__12657__C1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__A2 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__A2 (.DIODE(_02927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A1 (.DIODE(_02434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__B1 (.DIODE(_05662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__A2 (.DIODE(_06677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__B1 (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__B2 (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__A (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__B1 (.DIODE(_02348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__B1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__12700__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__C1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__A2 (.DIODE(_02440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__C1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A1 (.DIODE(_05123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12715__C1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__A1 (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12717__B (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__A1_N (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__12735__B1 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__B1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__C (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__A2 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12755__B1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12757__A2 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12759__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__A1 (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A1 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__C1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__B (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12775__C1 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A2 (.DIODE(_05069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__B1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12777__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12781__A (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__B (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__B1 (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__A2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__A2 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12791__B1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A2 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12793__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12797__A1 (.DIODE(_06667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__A1 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__A1 (.DIODE(_04917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12799__C1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__A0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12801__A (.DIODE(_04829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A (.DIODE(_04829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__S (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__12805__A (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A (.DIODE(_06085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__S (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__A (.DIODE(_06004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A (.DIODE(_06004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__S (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A (.DIODE(_05921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__A (.DIODE(_05921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__S (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__A (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__A (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__A (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__A (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A0 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__A (.DIODE(_05634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A (.DIODE(_05634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__A (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__A (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12862__A (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__S (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__A (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__A (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__12875__A (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12876__A (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12883__A (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12889__A (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12890__A (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12897__A (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12903__A (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12904__A (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12971__S (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__B (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__C (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__B (.DIODE(_04829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__B (.DIODE(_06004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__B (.DIODE(_06004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A (.DIODE(_05988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__A1 (.DIODE(_05988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__B (.DIODE(_05921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__B (.DIODE(_05921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__B (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__B (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__B (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__B (.DIODE(_05710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__B (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__B (.DIODE(_05774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__B (.DIODE(_05634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__B (.DIODE(_05634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__B (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__B (.DIODE(_05569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__B (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13025__B (.DIODE(_05461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__B (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__B (.DIODE(_05287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__B (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__B (.DIODE(_05363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__B (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13042__B (.DIODE(_04960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__B (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__B (.DIODE(_05189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__B (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13054__B (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__B (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13064__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13066__A2 (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13070__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13072__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__B2 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13080__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__A (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__B (.DIODE(_00251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13086__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13092__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__B2 (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__A2 (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__B2 (.DIODE(_00294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__13129__B (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__A (.DIODE(_04598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13139__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13143__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__13144__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__A (.DIODE(_00320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13148__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__13149__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__A (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13151__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13152__C1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13153__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__A1 (.DIODE(_00266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13154__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13155__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__A1 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13156__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__13157__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A1 (.DIODE(_00476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13158__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__13159__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13160__A1 (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13160__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A1 (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13163__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__13164__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__C1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13167__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13168__C1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13169__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__A1 (.DIODE(_00397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13172__C1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13173__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13174__C1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__C1 (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13177__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__13178__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13179__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__13182__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13183__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__A1 (.DIODE(_00203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13184__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A1 (.DIODE(_00208_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13187__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__A1 (.DIODE(_06725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13188__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__13189__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A1 (.DIODE(_00150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13192__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13193__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__A1 (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13194__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A1 (.DIODE(_00144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__13197__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__A1 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13198__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A1 (.DIODE(_00177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13201__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__A1 (.DIODE(_00516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13202__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13203__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A1 (.DIODE(_00812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13205__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__A1 (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13206__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13207__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__B1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13318__B2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13319__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13320__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13321__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13322__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13322__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13323__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13324__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13325__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13326__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13327__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13328__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13330__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13332__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13334__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13334__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13336__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13338__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13340__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13340__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13342__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13342__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13344__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13345__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13346__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13348__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13350__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13352__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13354__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13354__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__A2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13356__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13358__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13358__B1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13360__A2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13360__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13361__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13362__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13363__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13364__B1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13365__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13366__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13370__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13372__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13372__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13374__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13376__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13378__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13380__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__A2 (.DIODE(_06661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13382__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__13384__B1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__13385__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13386__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13389__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__13393__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__13395__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13396__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__13405__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__13409__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__13413__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__13417__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13418__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13420__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13421__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__13421__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__13422__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13422__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13423__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13424__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__13425__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__13426__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13426__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13427__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__13428__A2 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13428__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13429__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__13429__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__A2 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13430__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13431__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13432__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13433__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__13433__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13434__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13435__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13436__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__13437__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13438__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13439__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13440__C1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A1 (.DIODE(_00787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13441__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13442__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13443__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__A2 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__13444__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__13445__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__13446__C (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13447__A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13448__B1 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13450__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13452__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13453__A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13453__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13454__B1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13457__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13458__B2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13459__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13462__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__13463__B2 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__13466__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13467__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13470__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13475__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13480__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13486__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13490__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13491__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13492__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13496__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13497__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13500__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13501__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13502__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13505__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__13506__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__13507__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13510__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13511__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13512__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13515__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13516__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13517__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13520__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13521__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13524__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13525__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13528__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13529__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13532__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13533__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13533__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13537__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13538__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13538__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13541__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13542__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__13543__A (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA__13545__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13546__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13554__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13555__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__13558__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13559__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13562__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13563__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13566__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13567__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13568__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13571__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13572__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13576__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13577__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13581__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13582__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13584__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13586__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13587__A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13588__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13590__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13592__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13598__C (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__13601__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__13603__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13606__B1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__13683__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13685__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13686__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13687__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13688__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13690__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13691__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13692__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13701__CLK (.DIODE(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__13744__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__13748__A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(_00230_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(_00196_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(_00477_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_A (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(_00415_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(_00414_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(_00411_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(_00376_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(_00371_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(_00267_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(_00205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(_00205_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(_00157_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(_06681_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout14_A (.DIODE(_00337_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(_00327_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(_00326_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(_00320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(_00337_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout16_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(_06661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(_06661_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(_00413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(_06694_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(_06652_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(_04873_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(_04764_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(_04764_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(_00373_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_A (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_A (.DIODE(_00367_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_A (.DIODE(_00341_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(_00341_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(_00288_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(_00202_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(_02176_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(_00468_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(_00467_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(_00466_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(_00463_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout79_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(_00442_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(_00398_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(_00273_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(_00262_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout9_A (.DIODE(_02080_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap102_A (.DIODE(_00220_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap107_A (.DIODE(_00476_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap112_A (.DIODE(_00412_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap114_A (.DIODE(_00392_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap11_A (.DIODE(_02065_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap121_A (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap148_A (.DIODE(_00340_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap153_A (.DIODE(_00319_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap55_A (.DIODE(_06730_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap73_A (.DIODE(_00464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap78_A (.DIODE(_00446_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap81_A (.DIODE(_00443_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire101_A (.DIODE(_00229_));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire122_A (.DIODE(_00372_));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06743_ (.A(net459),
    .Y(_04401_));
 sky130_fd_sc_hd__inv_2 _06744_ (.A(net255),
    .Y(_04412_));
 sky130_fd_sc_hd__inv_2 _06745_ (.A(instruction[3]),
    .Y(_04423_));
 sky130_fd_sc_hd__inv_2 _06746_ (.A(instruction[5]),
    .Y(_04434_));
 sky130_fd_sc_hd__inv_2 _06747_ (.A(instruction[41]),
    .Y(_04445_));
 sky130_fd_sc_hd__inv_2 _06748_ (.A(net292),
    .Y(_04456_));
 sky130_fd_sc_hd__inv_2 _06749_ (.A(net289),
    .Y(_04467_));
 sky130_fd_sc_hd__inv_2 _06750_ (.A(net290),
    .Y(_04478_));
 sky130_fd_sc_hd__inv_2 _06751_ (.A(reg1_val[12]),
    .Y(_04489_));
 sky130_fd_sc_hd__inv_2 _06752_ (.A(reg1_val[14]),
    .Y(_04500_));
 sky130_fd_sc_hd__inv_2 _06753_ (.A(reg1_val[18]),
    .Y(_04511_));
 sky130_fd_sc_hd__inv_2 _06754_ (.A(reg1_val[20]),
    .Y(_04521_));
 sky130_fd_sc_hd__inv_2 _06755_ (.A(reg1_val[21]),
    .Y(_04532_));
 sky130_fd_sc_hd__inv_2 _06756_ (.A(reg1_val[22]),
    .Y(_04543_));
 sky130_fd_sc_hd__inv_2 _06757_ (.A(reg1_val[23]),
    .Y(_04554_));
 sky130_fd_sc_hd__inv_2 _06758_ (.A(reg1_val[24]),
    .Y(_04565_));
 sky130_fd_sc_hd__inv_2 _06759_ (.A(reg1_val[26]),
    .Y(_04576_));
 sky130_fd_sc_hd__inv_2 _06760_ (.A(reg1_val[28]),
    .Y(_04587_));
 sky130_fd_sc_hd__inv_6 _06761_ (.A(reg1_val[31]),
    .Y(_04598_));
 sky130_fd_sc_hd__inv_2 _06762_ (.A(net295),
    .Y(_04609_));
 sky130_fd_sc_hd__inv_2 _06763_ (.A(curr_PC[3]),
    .Y(_04620_));
 sky130_fd_sc_hd__inv_2 _06764_ (.A(rst),
    .Y(_04630_));
 sky130_fd_sc_hd__nand2_1 _06765_ (.A(pred_val),
    .B(instruction[1]),
    .Y(_04641_));
 sky130_fd_sc_hd__and4_4 _06766_ (.A(instruction[0]),
    .B(pred_val),
    .C(instruction[2]),
    .D(_04641_),
    .X(_04652_));
 sky130_fd_sc_hd__mux2_8 _06767_ (.A0(instruction[23]),
    .A1(instruction[16]),
    .S(_04652_),
    .X(reg1_idx[5]));
 sky130_fd_sc_hd__mux2_8 _06768_ (.A0(instruction[20]),
    .A1(instruction[13]),
    .S(_04652_),
    .X(reg1_idx[2]));
 sky130_fd_sc_hd__mux2_8 _06769_ (.A0(instruction[21]),
    .A1(instruction[14]),
    .S(_04652_),
    .X(reg1_idx[3]));
 sky130_fd_sc_hd__mux2_8 _06770_ (.A0(instruction[18]),
    .A1(instruction[11]),
    .S(_04652_),
    .X(reg1_idx[0]));
 sky130_fd_sc_hd__mux2_8 _06771_ (.A0(instruction[19]),
    .A1(instruction[12]),
    .S(_04652_),
    .X(reg1_idx[1]));
 sky130_fd_sc_hd__mux2_8 _06772_ (.A0(instruction[22]),
    .A1(instruction[15]),
    .S(_04652_),
    .X(reg1_idx[4]));
 sky130_fd_sc_hd__and3b_1 _06773_ (.A_N(instruction[0]),
    .B(pred_val),
    .C(instruction[2]),
    .X(_04723_));
 sky130_fd_sc_hd__and3_4 _06774_ (.A(_04423_),
    .B(_04641_),
    .C(_04723_),
    .X(is_load));
 sky130_fd_sc_hd__and3_4 _06775_ (.A(instruction[3]),
    .B(_04641_),
    .C(_04723_),
    .X(is_store));
 sky130_fd_sc_hd__and4bb_1 _06776_ (.A_N(instruction[0]),
    .B_N(instruction[2]),
    .C(instruction[1]),
    .D(pred_val),
    .X(_04753_));
 sky130_fd_sc_hd__or4bb_4 _06777_ (.A(instruction[0]),
    .B(instruction[2]),
    .C_N(instruction[1]),
    .D_N(pred_val),
    .X(_04764_));
 sky130_fd_sc_hd__and2_1 _06778_ (.A(reg2_val[31]),
    .B(net269),
    .X(_04775_));
 sky130_fd_sc_hd__o31a_1 _06779_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(pred_val),
    .X(_04786_));
 sky130_fd_sc_hd__o311a_4 _06780_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[41]),
    .C1(pred_val),
    .X(_04797_));
 sky130_fd_sc_hd__and4bb_2 _06781_ (.A_N(instruction[1]),
    .B_N(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04808_));
 sky130_fd_sc_hd__or4bb_1 _06782_ (.A(instruction[1]),
    .B(instruction[2]),
    .C_N(instruction[0]),
    .D_N(pred_val),
    .X(_04819_));
 sky130_fd_sc_hd__and2_2 _06783_ (.A(instruction[25]),
    .B(net266),
    .X(_04829_));
 sky130_fd_sc_hd__o211a_2 _06784_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .X(_04840_));
 sky130_fd_sc_hd__o211ai_1 _06785_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .Y(_04851_));
 sky130_fd_sc_hd__a21o_1 _06786_ (.A1(instruction[41]),
    .A2(_04808_),
    .B1(_04840_),
    .X(_04862_));
 sky130_fd_sc_hd__a21oi_4 _06787_ (.A1(instruction[41]),
    .A2(_04808_),
    .B1(_04840_),
    .Y(_04873_));
 sky130_fd_sc_hd__a221o_1 _06788_ (.A1(instruction[24]),
    .A2(_04797_),
    .B1(_04808_),
    .B2(instruction[41]),
    .C1(_04840_),
    .X(_04884_));
 sky130_fd_sc_hd__nand2_1 _06789_ (.A(net271),
    .B(_04884_),
    .Y(_04895_));
 sky130_fd_sc_hd__o21ba_1 _06790_ (.A1(_04445_),
    .A2(net226),
    .B1_N(_04775_),
    .X(_04906_));
 sky130_fd_sc_hd__a31o_4 _06791_ (.A1(instruction[41]),
    .A2(net271),
    .A3(_04884_),
    .B1(_04775_),
    .X(_04917_));
 sky130_fd_sc_hd__or2_2 _06792_ (.A(_04598_),
    .B(_04917_),
    .X(_04928_));
 sky130_fd_sc_hd__nand2_1 _06793_ (.A(_04598_),
    .B(_04917_),
    .Y(_04938_));
 sky130_fd_sc_hd__nand2_4 _06794_ (.A(_04928_),
    .B(_04938_),
    .Y(_04949_));
 sky130_fd_sc_hd__and2_4 _06795_ (.A(instruction[37]),
    .B(net266),
    .X(_04960_));
 sky130_fd_sc_hd__nor2_1 _06796_ (.A(net247),
    .B(_04960_),
    .Y(_04971_));
 sky130_fd_sc_hd__o2bb2a_2 _06797_ (.A1_N(reg2_val[27]),
    .A2_N(net268),
    .B1(net225),
    .B2(_04971_),
    .X(_04982_));
 sky130_fd_sc_hd__a2bb2o_1 _06798_ (.A1_N(_04971_),
    .A2_N(net225),
    .B1(net268),
    .B2(reg2_val[27]),
    .X(_04993_));
 sky130_fd_sc_hd__nor2_1 _06799_ (.A(reg1_val[27]),
    .B(_04993_),
    .Y(_05004_));
 sky130_fd_sc_hd__and2_1 _06800_ (.A(reg1_val[27]),
    .B(_04993_),
    .X(_05015_));
 sky130_fd_sc_hd__nand2_1 _06801_ (.A(reg1_val[27]),
    .B(_04993_),
    .Y(_05025_));
 sky130_fd_sc_hd__nor2_2 _06802_ (.A(_05004_),
    .B(_05015_),
    .Y(_05036_));
 sky130_fd_sc_hd__and2_4 _06803_ (.A(instruction[40]),
    .B(net266),
    .X(_05047_));
 sky130_fd_sc_hd__nor2_1 _06804_ (.A(_04873_),
    .B(_05047_),
    .Y(_05058_));
 sky130_fd_sc_hd__a2bb2o_4 _06805_ (.A1_N(_05058_),
    .A2_N(net225),
    .B1(net268),
    .B2(reg2_val[30]),
    .X(_05069_));
 sky130_fd_sc_hd__inv_2 _06806_ (.A(_05069_),
    .Y(_05080_));
 sky130_fd_sc_hd__xor2_4 _06807_ (.A(net288),
    .B(_05069_),
    .X(_05091_));
 sky130_fd_sc_hd__and2_4 _06808_ (.A(instruction[39]),
    .B(net266),
    .X(_05102_));
 sky130_fd_sc_hd__nor2_1 _06809_ (.A(net247),
    .B(_05102_),
    .Y(_05113_));
 sky130_fd_sc_hd__a2bb2o_4 _06810_ (.A1_N(_05113_),
    .A2_N(net225),
    .B1(net268),
    .B2(reg2_val[29]),
    .X(_05123_));
 sky130_fd_sc_hd__inv_2 _06811_ (.A(_05123_),
    .Y(_05134_));
 sky130_fd_sc_hd__nor2_1 _06812_ (.A(reg1_val[29]),
    .B(_05123_),
    .Y(_05145_));
 sky130_fd_sc_hd__inv_2 _06813_ (.A(_05145_),
    .Y(_05156_));
 sky130_fd_sc_hd__and2_1 _06814_ (.A(reg1_val[29]),
    .B(_05123_),
    .X(_05167_));
 sky130_fd_sc_hd__nor2_2 _06815_ (.A(_05145_),
    .B(_05167_),
    .Y(_05178_));
 sky130_fd_sc_hd__and2_4 _06816_ (.A(instruction[38]),
    .B(net266),
    .X(_05189_));
 sky130_fd_sc_hd__nor2_1 _06817_ (.A(_04873_),
    .B(_05189_),
    .Y(_05200_));
 sky130_fd_sc_hd__o2bb2a_2 _06818_ (.A1_N(reg2_val[28]),
    .A2_N(net268),
    .B1(net225),
    .B2(_05200_),
    .X(_05211_));
 sky130_fd_sc_hd__a2bb2o_2 _06819_ (.A1_N(_05200_),
    .A2_N(net225),
    .B1(net268),
    .B2(reg2_val[28]),
    .X(_05221_));
 sky130_fd_sc_hd__nand2_1 _06820_ (.A(_04587_),
    .B(_05211_),
    .Y(_05232_));
 sky130_fd_sc_hd__inv_2 _06821_ (.A(_05232_),
    .Y(_05243_));
 sky130_fd_sc_hd__nand2_1 _06822_ (.A(reg1_val[28]),
    .B(_05221_),
    .Y(_05254_));
 sky130_fd_sc_hd__and2_1 _06823_ (.A(_05232_),
    .B(_05254_),
    .X(_05265_));
 sky130_fd_sc_hd__nand2_1 _06824_ (.A(_05232_),
    .B(_05254_),
    .Y(_05276_));
 sky130_fd_sc_hd__and2_4 _06825_ (.A(instruction[35]),
    .B(net266),
    .X(_05287_));
 sky130_fd_sc_hd__nor2_1 _06826_ (.A(net247),
    .B(_05287_),
    .Y(_05298_));
 sky130_fd_sc_hd__a2bb2o_4 _06827_ (.A1_N(_05298_),
    .A2_N(net225),
    .B1(net269),
    .B2(reg2_val[25]),
    .X(_05308_));
 sky130_fd_sc_hd__inv_2 _06828_ (.A(_05308_),
    .Y(_05319_));
 sky130_fd_sc_hd__nor2_1 _06829_ (.A(reg1_val[25]),
    .B(_05308_),
    .Y(_05330_));
 sky130_fd_sc_hd__and2_1 _06830_ (.A(reg1_val[25]),
    .B(_05308_),
    .X(_05341_));
 sky130_fd_sc_hd__nor2_2 _06831_ (.A(_05330_),
    .B(_05341_),
    .Y(_05352_));
 sky130_fd_sc_hd__and2_4 _06832_ (.A(instruction[36]),
    .B(net266),
    .X(_05363_));
 sky130_fd_sc_hd__nor2_1 _06833_ (.A(net247),
    .B(_05363_),
    .Y(_05374_));
 sky130_fd_sc_hd__o2bb2a_2 _06834_ (.A1_N(reg2_val[26]),
    .A2_N(net268),
    .B1(net225),
    .B2(_05374_),
    .X(_05385_));
 sky130_fd_sc_hd__a2bb2o_4 _06835_ (.A1_N(_05374_),
    .A2_N(net225),
    .B1(net268),
    .B2(reg2_val[26]),
    .X(_05395_));
 sky130_fd_sc_hd__nand2_2 _06836_ (.A(reg1_val[26]),
    .B(_05395_),
    .Y(_05406_));
 sky130_fd_sc_hd__inv_2 _06837_ (.A(_05406_),
    .Y(_05417_));
 sky130_fd_sc_hd__nand2_1 _06838_ (.A(_04576_),
    .B(_05385_),
    .Y(_05428_));
 sky130_fd_sc_hd__and2_1 _06839_ (.A(_05406_),
    .B(_05428_),
    .X(_05439_));
 sky130_fd_sc_hd__nand2_1 _06840_ (.A(_05406_),
    .B(_05428_),
    .Y(_05450_));
 sky130_fd_sc_hd__and2_4 _06841_ (.A(instruction[34]),
    .B(net266),
    .X(_05461_));
 sky130_fd_sc_hd__nor2_1 _06842_ (.A(net247),
    .B(_05461_),
    .Y(_05471_));
 sky130_fd_sc_hd__o2bb2a_2 _06843_ (.A1_N(reg2_val[24]),
    .A2_N(net268),
    .B1(net225),
    .B2(_05471_),
    .X(_05482_));
 sky130_fd_sc_hd__a2bb2o_2 _06844_ (.A1_N(_05471_),
    .A2_N(net225),
    .B1(net268),
    .B2(reg2_val[24]),
    .X(_05493_));
 sky130_fd_sc_hd__nor2_1 _06845_ (.A(reg1_val[24]),
    .B(_05493_),
    .Y(_05504_));
 sky130_fd_sc_hd__nor2_1 _06846_ (.A(_04565_),
    .B(_05482_),
    .Y(_05515_));
 sky130_fd_sc_hd__nor2_2 _06847_ (.A(_05504_),
    .B(_05515_),
    .Y(_05526_));
 sky130_fd_sc_hd__or4_1 _06848_ (.A(_05036_),
    .B(_05091_),
    .C(_05178_),
    .D(_05265_),
    .X(_05536_));
 sky130_fd_sc_hd__or4_1 _06849_ (.A(_04949_),
    .B(_05352_),
    .C(_05439_),
    .D(_05526_),
    .X(_05547_));
 sky130_fd_sc_hd__or2_1 _06850_ (.A(_05536_),
    .B(_05547_),
    .X(_05558_));
 sky130_fd_sc_hd__and2_4 _06851_ (.A(instruction[33]),
    .B(net266),
    .X(_05569_));
 sky130_fd_sc_hd__nor2_1 _06852_ (.A(net247),
    .B(_05569_),
    .Y(_05580_));
 sky130_fd_sc_hd__o2bb2a_4 _06853_ (.A1_N(reg2_val[23]),
    .A2_N(net269),
    .B1(net225),
    .B2(_05580_),
    .X(_05591_));
 sky130_fd_sc_hd__nor2_1 _06854_ (.A(_04554_),
    .B(_05591_),
    .Y(_05602_));
 sky130_fd_sc_hd__and2_1 _06855_ (.A(_04554_),
    .B(_05591_),
    .X(_05612_));
 sky130_fd_sc_hd__nor2_2 _06856_ (.A(_05602_),
    .B(_05612_),
    .Y(_05623_));
 sky130_fd_sc_hd__and2_4 _06857_ (.A(instruction[32]),
    .B(net266),
    .X(_05634_));
 sky130_fd_sc_hd__nor2_1 _06858_ (.A(net247),
    .B(_05634_),
    .Y(_05645_));
 sky130_fd_sc_hd__o2bb2a_4 _06859_ (.A1_N(reg2_val[22]),
    .A2_N(net268),
    .B1(net225),
    .B2(_05645_),
    .X(_05656_));
 sky130_fd_sc_hd__a2bb2o_2 _06860_ (.A1_N(_05645_),
    .A2_N(net225),
    .B1(net268),
    .B2(reg2_val[22]),
    .X(_05666_));
 sky130_fd_sc_hd__nand2_1 _06861_ (.A(reg1_val[22]),
    .B(_05666_),
    .Y(_05677_));
 sky130_fd_sc_hd__nand2_1 _06862_ (.A(_04543_),
    .B(_05656_),
    .Y(_05688_));
 sky130_fd_sc_hd__and2_2 _06863_ (.A(_05677_),
    .B(_05688_),
    .X(_05699_));
 sky130_fd_sc_hd__and2_4 _06864_ (.A(instruction[30]),
    .B(net266),
    .X(_05710_));
 sky130_fd_sc_hd__nor2_1 _06865_ (.A(_04873_),
    .B(_05710_),
    .Y(_05720_));
 sky130_fd_sc_hd__o2bb2a_2 _06866_ (.A1_N(reg2_val[20]),
    .A2_N(net268),
    .B1(net225),
    .B2(_05720_),
    .X(_05731_));
 sky130_fd_sc_hd__and2_1 _06867_ (.A(_04521_),
    .B(_05731_),
    .X(_05742_));
 sky130_fd_sc_hd__nor2_1 _06868_ (.A(_04521_),
    .B(_05731_),
    .Y(_05753_));
 sky130_fd_sc_hd__nor2_2 _06869_ (.A(_05742_),
    .B(_05753_),
    .Y(_05764_));
 sky130_fd_sc_hd__o311a_4 _06870_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[31]),
    .C1(pred_val),
    .X(_05774_));
 sky130_fd_sc_hd__nor2_1 _06871_ (.A(_04873_),
    .B(_05774_),
    .Y(_05785_));
 sky130_fd_sc_hd__o2bb2a_2 _06872_ (.A1_N(reg2_val[21]),
    .A2_N(net268),
    .B1(net225),
    .B2(_05785_),
    .X(_05796_));
 sky130_fd_sc_hd__a2bb2o_1 _06873_ (.A1_N(_05785_),
    .A2_N(net226),
    .B1(net268),
    .B2(reg2_val[21]),
    .X(_05807_));
 sky130_fd_sc_hd__nor2_1 _06874_ (.A(_04532_),
    .B(_05796_),
    .Y(_05816_));
 sky130_fd_sc_hd__nor2_1 _06875_ (.A(reg1_val[21]),
    .B(_05807_),
    .Y(_05826_));
 sky130_fd_sc_hd__nor2_2 _06876_ (.A(_05816_),
    .B(_05826_),
    .Y(_05835_));
 sky130_fd_sc_hd__or4_1 _06877_ (.A(_05623_),
    .B(_05699_),
    .C(_05764_),
    .D(_05835_),
    .X(_05845_));
 sky130_fd_sc_hd__and2_4 _06878_ (.A(instruction[29]),
    .B(net266),
    .X(_05854_));
 sky130_fd_sc_hd__nor2_1 _06879_ (.A(_04873_),
    .B(_05854_),
    .Y(_05864_));
 sky130_fd_sc_hd__o2bb2a_4 _06880_ (.A1_N(reg2_val[19]),
    .A2_N(net268),
    .B1(net226),
    .B2(_05864_),
    .X(_05874_));
 sky130_fd_sc_hd__and2_1 _06881_ (.A(reg1_val[19]),
    .B(_05874_),
    .X(_05883_));
 sky130_fd_sc_hd__and2b_1 _06882_ (.A_N(reg1_val[19]),
    .B(_05874_),
    .X(_05893_));
 sky130_fd_sc_hd__and2b_1 _06883_ (.A_N(_05874_),
    .B(reg1_val[19]),
    .X(_05902_));
 sky130_fd_sc_hd__nor2_2 _06884_ (.A(_05893_),
    .B(_05902_),
    .Y(_05912_));
 sky130_fd_sc_hd__and2_4 _06885_ (.A(instruction[28]),
    .B(net266),
    .X(_05921_));
 sky130_fd_sc_hd__nor2_1 _06886_ (.A(_04873_),
    .B(_05921_),
    .Y(_05931_));
 sky130_fd_sc_hd__o2bb2a_4 _06887_ (.A1_N(reg2_val[18]),
    .A2_N(net267),
    .B1(net226),
    .B2(_05931_),
    .X(_05940_));
 sky130_fd_sc_hd__a2bb2o_2 _06888_ (.A1_N(_05931_),
    .A2_N(net226),
    .B1(net267),
    .B2(reg2_val[18]),
    .X(_05949_));
 sky130_fd_sc_hd__nand2_1 _06889_ (.A(reg1_val[18]),
    .B(_05940_),
    .Y(_05959_));
 sky130_fd_sc_hd__nor2_1 _06890_ (.A(reg1_val[18]),
    .B(_05949_),
    .Y(_05968_));
 sky130_fd_sc_hd__nand2_1 _06891_ (.A(_04511_),
    .B(_05940_),
    .Y(_05978_));
 sky130_fd_sc_hd__nor2_1 _06892_ (.A(_04511_),
    .B(_05940_),
    .Y(_05986_));
 sky130_fd_sc_hd__nor2_2 _06893_ (.A(_05968_),
    .B(_05986_),
    .Y(_05995_));
 sky130_fd_sc_hd__and2_4 _06894_ (.A(instruction[27]),
    .B(_04786_),
    .X(_06004_));
 sky130_fd_sc_hd__o311ai_2 _06895_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[27]),
    .C1(pred_val),
    .Y(_06013_));
 sky130_fd_sc_hd__nor2_1 _06896_ (.A(net246),
    .B(_06004_),
    .Y(_06022_));
 sky130_fd_sc_hd__o2bb2a_4 _06897_ (.A1_N(reg2_val[17]),
    .A2_N(net267),
    .B1(net226),
    .B2(_06022_),
    .X(_06031_));
 sky130_fd_sc_hd__a2bb2o_2 _06898_ (.A1_N(_06022_),
    .A2_N(net226),
    .B1(net267),
    .B2(reg2_val[17]),
    .X(_06041_));
 sky130_fd_sc_hd__nand2_1 _06899_ (.A(reg1_val[17]),
    .B(_06031_),
    .Y(_06050_));
 sky130_fd_sc_hd__or2_1 _06900_ (.A(reg1_val[17]),
    .B(_06041_),
    .X(_06059_));
 sky130_fd_sc_hd__nand2_1 _06901_ (.A(reg1_val[17]),
    .B(_06041_),
    .Y(_06068_));
 sky130_fd_sc_hd__and2_2 _06902_ (.A(_06059_),
    .B(_06068_),
    .X(_06076_));
 sky130_fd_sc_hd__and2_2 _06903_ (.A(instruction[26]),
    .B(net266),
    .X(_06085_));
 sky130_fd_sc_hd__nand2_1 _06904_ (.A(instruction[26]),
    .B(net266),
    .Y(_06094_));
 sky130_fd_sc_hd__nor2_1 _06905_ (.A(net247),
    .B(_06085_),
    .Y(_06103_));
 sky130_fd_sc_hd__o2bb2a_2 _06906_ (.A1_N(reg2_val[16]),
    .A2_N(net267),
    .B1(net226),
    .B2(_06103_),
    .X(_06112_));
 sky130_fd_sc_hd__a2bb2o_1 _06907_ (.A1_N(_06103_),
    .A2_N(net226),
    .B1(net267),
    .B2(reg2_val[16]),
    .X(_06121_));
 sky130_fd_sc_hd__nand2_1 _06908_ (.A(reg1_val[16]),
    .B(_06112_),
    .Y(_06129_));
 sky130_fd_sc_hd__or2_1 _06909_ (.A(reg1_val[16]),
    .B(_06121_),
    .X(_06135_));
 sky130_fd_sc_hd__inv_2 _06910_ (.A(_06135_),
    .Y(_06141_));
 sky130_fd_sc_hd__and2_1 _06911_ (.A(reg1_val[16]),
    .B(_06121_),
    .X(_06147_));
 sky130_fd_sc_hd__nor2_1 _06912_ (.A(_06141_),
    .B(_06147_),
    .Y(_06153_));
 sky130_fd_sc_hd__and2_1 _06913_ (.A(reg2_val[15]),
    .B(net269),
    .X(_06159_));
 sky130_fd_sc_hd__a31o_4 _06914_ (.A1(net271),
    .A2(_04797_),
    .A3(net247),
    .B1(_06159_),
    .X(_06165_));
 sky130_fd_sc_hd__nand2b_1 _06915_ (.A_N(_06165_),
    .B(reg1_val[15]),
    .Y(_06174_));
 sky130_fd_sc_hd__or2_1 _06916_ (.A(reg1_val[15]),
    .B(_06165_),
    .X(_06185_));
 sky130_fd_sc_hd__nand2_1 _06917_ (.A(reg1_val[15]),
    .B(_06165_),
    .Y(_06196_));
 sky130_fd_sc_hd__and2_1 _06918_ (.A(_06185_),
    .B(_06196_),
    .X(_06207_));
 sky130_fd_sc_hd__nand2_1 _06919_ (.A(_06185_),
    .B(_06196_),
    .Y(_06218_));
 sky130_fd_sc_hd__and2_1 _06920_ (.A(reg2_val[14]),
    .B(_04764_),
    .X(_06229_));
 sky130_fd_sc_hd__a31o_4 _06921_ (.A1(net271),
    .A2(net246),
    .A3(_05047_),
    .B1(_06229_),
    .X(_06240_));
 sky130_fd_sc_hd__inv_2 _06922_ (.A(_06240_),
    .Y(_06251_));
 sky130_fd_sc_hd__or2_1 _06923_ (.A(_04500_),
    .B(_06240_),
    .X(_06262_));
 sky130_fd_sc_hd__or2_1 _06924_ (.A(reg1_val[14]),
    .B(_06240_),
    .X(_06273_));
 sky130_fd_sc_hd__nand2_2 _06925_ (.A(reg1_val[14]),
    .B(_06240_),
    .Y(_06284_));
 sky130_fd_sc_hd__and2_1 _06926_ (.A(_06273_),
    .B(_06284_),
    .X(_06291_));
 sky130_fd_sc_hd__nand2_1 _06927_ (.A(_06273_),
    .B(_06284_),
    .Y(_06297_));
 sky130_fd_sc_hd__and3_1 _06928_ (.A(net270),
    .B(net247),
    .C(_05102_),
    .X(_06303_));
 sky130_fd_sc_hd__a21o_2 _06929_ (.A1(reg2_val[13]),
    .A2(net267),
    .B1(_06303_),
    .X(_06309_));
 sky130_fd_sc_hd__a21oi_4 _06930_ (.A1(reg2_val[13]),
    .A2(net267),
    .B1(_06303_),
    .Y(_06315_));
 sky130_fd_sc_hd__nand2_1 _06931_ (.A(reg1_val[13]),
    .B(_06315_),
    .Y(_06321_));
 sky130_fd_sc_hd__or2_1 _06932_ (.A(reg1_val[13]),
    .B(_06309_),
    .X(_06327_));
 sky130_fd_sc_hd__nand2_1 _06933_ (.A(reg1_val[13]),
    .B(_06309_),
    .Y(_06333_));
 sky130_fd_sc_hd__nand2_1 _06934_ (.A(_06327_),
    .B(_06333_),
    .Y(_06339_));
 sky130_fd_sc_hd__inv_2 _06935_ (.A(_06339_),
    .Y(_06345_));
 sky130_fd_sc_hd__and3_1 _06936_ (.A(net271),
    .B(net246),
    .C(_05189_),
    .X(_06351_));
 sky130_fd_sc_hd__a21o_1 _06937_ (.A1(reg2_val[12]),
    .A2(net267),
    .B1(_06351_),
    .X(_06357_));
 sky130_fd_sc_hd__a21oi_4 _06938_ (.A1(reg2_val[12]),
    .A2(net267),
    .B1(_06351_),
    .Y(_06363_));
 sky130_fd_sc_hd__nand2_1 _06939_ (.A(reg1_val[12]),
    .B(_06363_),
    .Y(_06372_));
 sky130_fd_sc_hd__nand2_1 _06940_ (.A(_04489_),
    .B(_06363_),
    .Y(_06381_));
 sky130_fd_sc_hd__nand2_1 _06941_ (.A(reg1_val[12]),
    .B(_06357_),
    .Y(_06390_));
 sky130_fd_sc_hd__and2_1 _06942_ (.A(_06381_),
    .B(_06390_),
    .X(_06399_));
 sky130_fd_sc_hd__nand2_1 _06943_ (.A(_06381_),
    .B(_06390_),
    .Y(_06408_));
 sky130_fd_sc_hd__and2_1 _06944_ (.A(reg2_val[11]),
    .B(net267),
    .X(_06417_));
 sky130_fd_sc_hd__a31o_2 _06945_ (.A1(net270),
    .A2(net246),
    .A3(_04960_),
    .B1(_06417_),
    .X(_06426_));
 sky130_fd_sc_hd__a31oi_4 _06946_ (.A1(net270),
    .A2(net246),
    .A3(_04960_),
    .B1(_06417_),
    .Y(_06435_));
 sky130_fd_sc_hd__nand2_1 _06947_ (.A(net290),
    .B(_06435_),
    .Y(_06443_));
 sky130_fd_sc_hd__nand2_1 _06948_ (.A(_04478_),
    .B(_06435_),
    .Y(_06452_));
 sky130_fd_sc_hd__nand2_1 _06949_ (.A(net290),
    .B(_06426_),
    .Y(_06461_));
 sky130_fd_sc_hd__nand2_2 _06950_ (.A(_06452_),
    .B(_06461_),
    .Y(_06469_));
 sky130_fd_sc_hd__inv_2 _06951_ (.A(_06469_),
    .Y(_06478_));
 sky130_fd_sc_hd__and2_2 _06952_ (.A(reg2_val[10]),
    .B(net267),
    .X(_06487_));
 sky130_fd_sc_hd__a31o_2 _06953_ (.A1(net270),
    .A2(net246),
    .A3(_05363_),
    .B1(_06487_),
    .X(_06495_));
 sky130_fd_sc_hd__a31oi_4 _06954_ (.A1(net270),
    .A2(net246),
    .A3(_05363_),
    .B1(_06487_),
    .Y(_06502_));
 sky130_fd_sc_hd__nand2_1 _06955_ (.A(reg1_val[10]),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__nor2_1 _06956_ (.A(reg1_val[10]),
    .B(_06495_),
    .Y(_06504_));
 sky130_fd_sc_hd__nand2_1 _06957_ (.A(reg1_val[10]),
    .B(_06495_),
    .Y(_06505_));
 sky130_fd_sc_hd__nand2b_2 _06958_ (.A_N(_06504_),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__inv_2 _06959_ (.A(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__and2_1 _06960_ (.A(reg2_val[9]),
    .B(net267),
    .X(_06508_));
 sky130_fd_sc_hd__a31o_4 _06961_ (.A1(net271),
    .A2(net246),
    .A3(_05287_),
    .B1(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__nand2b_1 _06962_ (.A_N(_06509_),
    .B(reg1_val[9]),
    .Y(_06510_));
 sky130_fd_sc_hd__nor2_1 _06963_ (.A(reg1_val[9]),
    .B(_06509_),
    .Y(_06511_));
 sky130_fd_sc_hd__nand2_1 _06964_ (.A(reg1_val[9]),
    .B(_06509_),
    .Y(_06512_));
 sky130_fd_sc_hd__and2b_1 _06965_ (.A_N(_06511_),
    .B(_06512_),
    .X(_06513_));
 sky130_fd_sc_hd__nand2b_1 _06966_ (.A_N(_06511_),
    .B(_06512_),
    .Y(_06514_));
 sky130_fd_sc_hd__and2_1 _06967_ (.A(reg2_val[8]),
    .B(net267),
    .X(_06515_));
 sky130_fd_sc_hd__a31o_2 _06968_ (.A1(net270),
    .A2(net246),
    .A3(_05461_),
    .B1(_06515_),
    .X(_06516_));
 sky130_fd_sc_hd__a31oi_4 _06969_ (.A1(net270),
    .A2(net246),
    .A3(_05461_),
    .B1(_06515_),
    .Y(_06517_));
 sky130_fd_sc_hd__and2_1 _06970_ (.A(reg1_val[8]),
    .B(_06517_),
    .X(_06518_));
 sky130_fd_sc_hd__nor2_1 _06971_ (.A(reg1_val[8]),
    .B(_06516_),
    .Y(_06519_));
 sky130_fd_sc_hd__nand2_1 _06972_ (.A(reg1_val[8]),
    .B(_06516_),
    .Y(_06520_));
 sky130_fd_sc_hd__and2b_1 _06973_ (.A_N(_06519_),
    .B(_06520_),
    .X(_06521_));
 sky130_fd_sc_hd__and2_1 _06974_ (.A(reg2_val[7]),
    .B(net267),
    .X(_06522_));
 sky130_fd_sc_hd__a31o_4 _06975_ (.A1(net270),
    .A2(net247),
    .A3(_05569_),
    .B1(_06522_),
    .X(_06523_));
 sky130_fd_sc_hd__nand2b_1 _06976_ (.A_N(_06523_),
    .B(net287),
    .Y(_06524_));
 sky130_fd_sc_hd__nor2_1 _06977_ (.A(net287),
    .B(_06523_),
    .Y(_06525_));
 sky130_fd_sc_hd__nand2_1 _06978_ (.A(net287),
    .B(_06523_),
    .Y(_06526_));
 sky130_fd_sc_hd__and2b_1 _06979_ (.A_N(_06525_),
    .B(_06526_),
    .X(_06527_));
 sky130_fd_sc_hd__and2_1 _06980_ (.A(reg2_val[6]),
    .B(net267),
    .X(_06528_));
 sky130_fd_sc_hd__a31o_4 _06981_ (.A1(net271),
    .A2(net247),
    .A3(_05634_),
    .B1(_06528_),
    .X(_06529_));
 sky130_fd_sc_hd__inv_2 _06982_ (.A(_06529_),
    .Y(_06530_));
 sky130_fd_sc_hd__nand2_1 _06983_ (.A(reg1_val[6]),
    .B(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__nor2_1 _06984_ (.A(reg1_val[6]),
    .B(_06529_),
    .Y(_06532_));
 sky130_fd_sc_hd__and2_1 _06985_ (.A(reg1_val[6]),
    .B(_06529_),
    .X(_06533_));
 sky130_fd_sc_hd__nand2_1 _06986_ (.A(reg1_val[6]),
    .B(_06529_),
    .Y(_06534_));
 sky130_fd_sc_hd__nor2_1 _06987_ (.A(_06532_),
    .B(_06533_),
    .Y(_06535_));
 sky130_fd_sc_hd__o2111a_1 _06988_ (.A1(_04445_),
    .A2(_04819_),
    .B1(_04851_),
    .C1(_05774_),
    .D1(net271),
    .X(_06536_));
 sky130_fd_sc_hd__or3b_2 _06989_ (.A(net269),
    .B(_04862_),
    .C_N(_05774_),
    .X(_06537_));
 sky130_fd_sc_hd__a21oi_4 _06990_ (.A1(reg2_val[5]),
    .A2(net269),
    .B1(net245),
    .Y(_06538_));
 sky130_fd_sc_hd__a21o_2 _06991_ (.A1(reg2_val[5]),
    .A2(net269),
    .B1(net245),
    .X(_06539_));
 sky130_fd_sc_hd__nand2_1 _06992_ (.A(reg1_val[5]),
    .B(_06538_),
    .Y(_06540_));
 sky130_fd_sc_hd__nand2_2 _06993_ (.A(reg1_val[5]),
    .B(_06539_),
    .Y(_06541_));
 sky130_fd_sc_hd__inv_2 _06994_ (.A(_06541_),
    .Y(_06542_));
 sky130_fd_sc_hd__nor2_1 _06995_ (.A(reg1_val[5]),
    .B(_06539_),
    .Y(_06543_));
 sky130_fd_sc_hd__nor2_1 _06996_ (.A(_06542_),
    .B(_06543_),
    .Y(_06544_));
 sky130_fd_sc_hd__and2_1 _06997_ (.A(reg2_val[4]),
    .B(net269),
    .X(_06545_));
 sky130_fd_sc_hd__a31o_1 _06998_ (.A1(net270),
    .A2(net246),
    .A3(_05710_),
    .B1(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__a31oi_4 _06999_ (.A1(net270),
    .A2(net246),
    .A3(_05710_),
    .B1(_06545_),
    .Y(_06547_));
 sky130_fd_sc_hd__nand2_1 _07000_ (.A(reg1_val[4]),
    .B(net220),
    .Y(_06548_));
 sky130_fd_sc_hd__nor2_1 _07001_ (.A(reg1_val[4]),
    .B(net222),
    .Y(_06549_));
 sky130_fd_sc_hd__nand2_2 _07002_ (.A(reg1_val[4]),
    .B(net222),
    .Y(_06550_));
 sky130_fd_sc_hd__and2b_1 _07003_ (.A_N(_06549_),
    .B(_06550_),
    .X(_06551_));
 sky130_fd_sc_hd__and2_1 _07004_ (.A(reg2_val[3]),
    .B(net269),
    .X(_06552_));
 sky130_fd_sc_hd__a31oi_4 _07005_ (.A1(net270),
    .A2(net246),
    .A3(_05854_),
    .B1(_06552_),
    .Y(_06553_));
 sky130_fd_sc_hd__a31o_4 _07006_ (.A1(net270),
    .A2(net246),
    .A3(_05854_),
    .B1(_06552_),
    .X(_06554_));
 sky130_fd_sc_hd__nand2_1 _07007_ (.A(reg1_val[3]),
    .B(_06553_),
    .Y(_06555_));
 sky130_fd_sc_hd__nor2_1 _07008_ (.A(reg1_val[3]),
    .B(_06554_),
    .Y(_06556_));
 sky130_fd_sc_hd__nand2_2 _07009_ (.A(reg1_val[3]),
    .B(_06554_),
    .Y(_06557_));
 sky130_fd_sc_hd__and2b_1 _07010_ (.A_N(_06556_),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__and2_1 _07011_ (.A(reg2_val[2]),
    .B(net269),
    .X(_06559_));
 sky130_fd_sc_hd__a31oi_4 _07012_ (.A1(net270),
    .A2(net246),
    .A3(_05921_),
    .B1(_06559_),
    .Y(_06560_));
 sky130_fd_sc_hd__a31o_1 _07013_ (.A1(net270),
    .A2(net246),
    .A3(_05921_),
    .B1(_06559_),
    .X(_06561_));
 sky130_fd_sc_hd__nand2_1 _07014_ (.A(reg1_val[2]),
    .B(net217),
    .Y(_06562_));
 sky130_fd_sc_hd__nand2_1 _07015_ (.A(reg1_val[2]),
    .B(net216),
    .Y(_06563_));
 sky130_fd_sc_hd__nor2_1 _07016_ (.A(reg1_val[2]),
    .B(net216),
    .Y(_06564_));
 sky130_fd_sc_hd__xnor2_2 _07017_ (.A(reg1_val[2]),
    .B(_06560_),
    .Y(_06565_));
 sky130_fd_sc_hd__nand2_2 _07018_ (.A(reg2_val[1]),
    .B(net269),
    .Y(_06566_));
 sky130_fd_sc_hd__a2111o_4 _07019_ (.A1(instruction[41]),
    .A2(_04808_),
    .B1(_04840_),
    .C1(_06013_),
    .D1(net269),
    .X(_06567_));
 sky130_fd_sc_hd__and2_1 _07020_ (.A(_06566_),
    .B(_06567_),
    .X(_06568_));
 sky130_fd_sc_hd__nand2_8 _07021_ (.A(_06566_),
    .B(_06567_),
    .Y(_06569_));
 sky130_fd_sc_hd__nand2_1 _07022_ (.A(net289),
    .B(net214),
    .Y(_06570_));
 sky130_fd_sc_hd__a21oi_1 _07023_ (.A1(_06566_),
    .A2(_06567_),
    .B1(_04467_),
    .Y(_06571_));
 sky130_fd_sc_hd__nand2_1 _07024_ (.A(net289),
    .B(_06569_),
    .Y(_06572_));
 sky130_fd_sc_hd__and3_1 _07025_ (.A(_04467_),
    .B(_06566_),
    .C(_06567_),
    .X(_06573_));
 sky130_fd_sc_hd__nor2_1 _07026_ (.A(_06571_),
    .B(_06573_),
    .Y(_06574_));
 sky130_fd_sc_hd__and2_1 _07027_ (.A(reg2_val[0]),
    .B(net269),
    .X(_06575_));
 sky130_fd_sc_hd__a31oi_2 _07028_ (.A1(net270),
    .A2(net247),
    .A3(_06085_),
    .B1(_06575_),
    .Y(_06576_));
 sky130_fd_sc_hd__a31o_1 _07029_ (.A1(net270),
    .A2(net247),
    .A3(_06085_),
    .B1(_06575_),
    .X(_06577_));
 sky130_fd_sc_hd__nor2_1 _07030_ (.A(net291),
    .B(net211),
    .Y(_06578_));
 sky130_fd_sc_hd__a2bb2o_1 _07031_ (.A1_N(_06571_),
    .A2_N(_06573_),
    .B1(net206),
    .B2(net285),
    .X(_06579_));
 sky130_fd_sc_hd__a21o_1 _07032_ (.A1(_06570_),
    .A2(_06579_),
    .B1(_06565_),
    .X(_06580_));
 sky130_fd_sc_hd__a21o_1 _07033_ (.A1(_06562_),
    .A2(_06580_),
    .B1(_06558_),
    .X(_06581_));
 sky130_fd_sc_hd__a21o_1 _07034_ (.A1(_06555_),
    .A2(_06581_),
    .B1(_06551_),
    .X(_06582_));
 sky130_fd_sc_hd__a21o_1 _07035_ (.A1(_06548_),
    .A2(_06582_),
    .B1(_06544_),
    .X(_06583_));
 sky130_fd_sc_hd__a21o_1 _07036_ (.A1(_06540_),
    .A2(_06583_),
    .B1(_06535_),
    .X(_06584_));
 sky130_fd_sc_hd__a21o_1 _07037_ (.A1(_06531_),
    .A2(_06584_),
    .B1(_06527_),
    .X(_06585_));
 sky130_fd_sc_hd__a21oi_1 _07038_ (.A1(_06524_),
    .A2(_06585_),
    .B1(_06521_),
    .Y(_06586_));
 sky130_fd_sc_hd__o21ai_1 _07039_ (.A1(_06518_),
    .A2(_06586_),
    .B1(_06514_),
    .Y(_06587_));
 sky130_fd_sc_hd__a21o_1 _07040_ (.A1(_06510_),
    .A2(_06587_),
    .B1(_06507_),
    .X(_06588_));
 sky130_fd_sc_hd__a21o_1 _07041_ (.A1(_06503_),
    .A2(_06588_),
    .B1(_06478_),
    .X(_06589_));
 sky130_fd_sc_hd__a21o_1 _07042_ (.A1(_06443_),
    .A2(_06589_),
    .B1(_06399_),
    .X(_06590_));
 sky130_fd_sc_hd__a21o_1 _07043_ (.A1(_06372_),
    .A2(_06590_),
    .B1(_06345_),
    .X(_06591_));
 sky130_fd_sc_hd__a21o_1 _07044_ (.A1(_06321_),
    .A2(_06591_),
    .B1(_06291_),
    .X(_06592_));
 sky130_fd_sc_hd__a21o_1 _07045_ (.A1(_06262_),
    .A2(_06592_),
    .B1(_06207_),
    .X(_06593_));
 sky130_fd_sc_hd__a21o_1 _07046_ (.A1(_06174_),
    .A2(_06593_),
    .B1(_06153_),
    .X(_06594_));
 sky130_fd_sc_hd__a21o_1 _07047_ (.A1(_06129_),
    .A2(_06594_),
    .B1(_06076_),
    .X(_06595_));
 sky130_fd_sc_hd__a21o_1 _07048_ (.A1(_06050_),
    .A2(_06595_),
    .B1(_05995_),
    .X(_06596_));
 sky130_fd_sc_hd__a21oi_1 _07049_ (.A1(_05959_),
    .A2(_06596_),
    .B1(_05912_),
    .Y(_06597_));
 sky130_fd_sc_hd__nor2_1 _07050_ (.A(_05883_),
    .B(_06597_),
    .Y(_06598_));
 sky130_fd_sc_hd__o21bai_1 _07051_ (.A1(_05883_),
    .A2(_06597_),
    .B1_N(_05845_),
    .Y(_06599_));
 sky130_fd_sc_hd__nand2_1 _07052_ (.A(reg1_val[23]),
    .B(_05591_),
    .Y(_06600_));
 sky130_fd_sc_hd__nand2_1 _07053_ (.A(reg1_val[22]),
    .B(_05656_),
    .Y(_06601_));
 sky130_fd_sc_hd__nand2_1 _07054_ (.A(reg1_val[21]),
    .B(_05796_),
    .Y(_06602_));
 sky130_fd_sc_hd__nand2_1 _07055_ (.A(reg1_val[20]),
    .B(_05731_),
    .Y(_06603_));
 sky130_fd_sc_hd__o21a_1 _07056_ (.A1(_05835_),
    .A2(_06603_),
    .B1(_06602_),
    .X(_06604_));
 sky130_fd_sc_hd__o21a_1 _07057_ (.A1(_05699_),
    .A2(_06604_),
    .B1(_06601_),
    .X(_06605_));
 sky130_fd_sc_hd__o21a_1 _07058_ (.A1(_05623_),
    .A2(_06605_),
    .B1(_06600_),
    .X(_06606_));
 sky130_fd_sc_hd__and2_1 _07059_ (.A(_06599_),
    .B(_06606_),
    .X(_06607_));
 sky130_fd_sc_hd__nand2_1 _07060_ (.A(net288),
    .B(_05080_),
    .Y(_06608_));
 sky130_fd_sc_hd__nand2_1 _07061_ (.A(reg1_val[29]),
    .B(_05134_),
    .Y(_06609_));
 sky130_fd_sc_hd__nand2_1 _07062_ (.A(reg1_val[28]),
    .B(_05211_),
    .Y(_06610_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(reg1_val[27]),
    .B(_04982_),
    .Y(_06611_));
 sky130_fd_sc_hd__nand2_1 _07064_ (.A(reg1_val[26]),
    .B(_05385_),
    .Y(_06612_));
 sky130_fd_sc_hd__nand2_1 _07065_ (.A(reg1_val[25]),
    .B(_05319_),
    .Y(_06613_));
 sky130_fd_sc_hd__nand2_1 _07066_ (.A(reg1_val[24]),
    .B(_05482_),
    .Y(_06614_));
 sky130_fd_sc_hd__o21a_1 _07067_ (.A1(_05352_),
    .A2(_06614_),
    .B1(_06613_),
    .X(_06615_));
 sky130_fd_sc_hd__o21a_1 _07068_ (.A1(_05439_),
    .A2(_06615_),
    .B1(_06612_),
    .X(_06616_));
 sky130_fd_sc_hd__o21a_1 _07069_ (.A1(_05036_),
    .A2(_06616_),
    .B1(_06611_),
    .X(_06617_));
 sky130_fd_sc_hd__o21a_1 _07070_ (.A1(_05265_),
    .A2(_06617_),
    .B1(_06610_),
    .X(_06618_));
 sky130_fd_sc_hd__o21a_1 _07071_ (.A1(_05178_),
    .A2(_06618_),
    .B1(_06609_),
    .X(_06619_));
 sky130_fd_sc_hd__o21a_1 _07072_ (.A1(_05091_),
    .A2(_06619_),
    .B1(_06608_),
    .X(_06620_));
 sky130_fd_sc_hd__o21ba_1 _07073_ (.A1(_05558_),
    .A2(_06607_),
    .B1_N(instruction[6]),
    .X(_06621_));
 sky130_fd_sc_hd__o211a_1 _07074_ (.A1(_04949_),
    .A2(_06620_),
    .B1(_06621_),
    .C1(_04928_),
    .X(_06622_));
 sky130_fd_sc_hd__inv_2 _07075_ (.A(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__a21o_1 _07076_ (.A1(_06599_),
    .A2(_06606_),
    .B1(_05526_),
    .X(_06624_));
 sky130_fd_sc_hd__and2_1 _07077_ (.A(_06614_),
    .B(_06624_),
    .X(_06625_));
 sky130_fd_sc_hd__a21o_1 _07078_ (.A1(_06614_),
    .A2(_06624_),
    .B1(_05352_),
    .X(_06626_));
 sky130_fd_sc_hd__nand2_1 _07079_ (.A(_06613_),
    .B(_06626_),
    .Y(_06627_));
 sky130_fd_sc_hd__a21o_1 _07080_ (.A1(_06613_),
    .A2(_06626_),
    .B1(_05439_),
    .X(_06628_));
 sky130_fd_sc_hd__a21o_1 _07081_ (.A1(_06612_),
    .A2(_06628_),
    .B1(_05036_),
    .X(_06629_));
 sky130_fd_sc_hd__nand2_1 _07082_ (.A(_06611_),
    .B(_06629_),
    .Y(_06630_));
 sky130_fd_sc_hd__a21boi_1 _07083_ (.A1(_05276_),
    .A2(_06630_),
    .B1_N(_06610_),
    .Y(_06631_));
 sky130_fd_sc_hd__o21a_1 _07084_ (.A1(_05178_),
    .A2(_06631_),
    .B1(_06609_),
    .X(_06632_));
 sky130_fd_sc_hd__o21ai_1 _07085_ (.A1(_05091_),
    .A2(_06632_),
    .B1(_06608_),
    .Y(_06633_));
 sky130_fd_sc_hd__o21ai_1 _07086_ (.A1(_04949_),
    .A2(_06633_),
    .B1(_04928_),
    .Y(_06634_));
 sky130_fd_sc_hd__a21oi_1 _07087_ (.A1(instruction[6]),
    .A2(_06634_),
    .B1(_06622_),
    .Y(_06635_));
 sky130_fd_sc_hd__nor2_2 _07088_ (.A(instruction[3]),
    .B(net298),
    .Y(_06636_));
 sky130_fd_sc_hd__nand2_2 _07089_ (.A(net291),
    .B(net206),
    .Y(_06637_));
 sky130_fd_sc_hd__nand2_1 _07090_ (.A(net285),
    .B(net211),
    .Y(_06638_));
 sky130_fd_sc_hd__nand2_1 _07091_ (.A(_06637_),
    .B(_06638_),
    .Y(_06639_));
 sky130_fd_sc_hd__or4_1 _07092_ (.A(_05912_),
    .B(_05995_),
    .C(_06076_),
    .D(_06153_),
    .X(_06640_));
 sky130_fd_sc_hd__nand2_1 _07093_ (.A(_06469_),
    .B(_06506_),
    .Y(_06641_));
 sky130_fd_sc_hd__and4_1 _07094_ (.A(_06218_),
    .B(_06297_),
    .C(_06339_),
    .D(_06408_),
    .X(_06642_));
 sky130_fd_sc_hd__or4b_1 _07095_ (.A(_06513_),
    .B(_06527_),
    .C(_06641_),
    .D_N(_06642_),
    .X(_06643_));
 sky130_fd_sc_hd__or4_1 _07096_ (.A(_06535_),
    .B(_06544_),
    .C(_06551_),
    .D(_06558_),
    .X(_06644_));
 sky130_fd_sc_hd__or4b_1 _07097_ (.A(_06521_),
    .B(_06565_),
    .C(_06574_),
    .D_N(_06639_),
    .X(_06645_));
 sky130_fd_sc_hd__or4_1 _07098_ (.A(_06640_),
    .B(_06643_),
    .C(_06644_),
    .D(_06645_),
    .X(_06646_));
 sky130_fd_sc_hd__or3_1 _07099_ (.A(_05558_),
    .B(_05845_),
    .C(_06646_),
    .X(_06647_));
 sky130_fd_sc_hd__mux2_1 _07100_ (.A0(_06647_),
    .A1(_04949_),
    .S(net297),
    .X(_06648_));
 sky130_fd_sc_hd__or3_1 _07101_ (.A(instruction[3]),
    .B(net298),
    .C(_06648_),
    .X(_06649_));
 sky130_fd_sc_hd__nand2_1 _07102_ (.A(instruction[3]),
    .B(net298),
    .Y(_06650_));
 sky130_fd_sc_hd__o221a_2 _07103_ (.A1(_04423_),
    .A2(_06635_),
    .B1(_06647_),
    .B2(_06650_),
    .C1(_06649_),
    .X(_06651_));
 sky130_fd_sc_hd__xnor2_4 _07104_ (.A(instruction[5]),
    .B(_06651_),
    .Y(dest_pred_val));
 sky130_fd_sc_hd__and2_4 _07105_ (.A(instruction[1]),
    .B(_04723_),
    .X(_06652_));
 sky130_fd_sc_hd__nand2_1 _07106_ (.A(instruction[1]),
    .B(_04723_),
    .Y(_06653_));
 sky130_fd_sc_hd__a21o_4 _07107_ (.A1(_04652_),
    .A2(dest_pred_val),
    .B1(net243),
    .X(take_branch));
 sky130_fd_sc_hd__and4_1 _07108_ (.A(reg1_idx[5]),
    .B(reg1_idx[2]),
    .C(reg1_idx[3]),
    .D(_06652_),
    .X(_06654_));
 sky130_fd_sc_hd__and4_4 _07109_ (.A(reg1_idx[0]),
    .B(reg1_idx[1]),
    .C(reg1_idx[4]),
    .D(_06654_),
    .X(int_return));
 sky130_fd_sc_hd__nand2_1 _07110_ (.A(net269),
    .B(_04819_),
    .Y(_06655_));
 sky130_fd_sc_hd__and2_2 _07111_ (.A(net297),
    .B(_04434_),
    .X(_06656_));
 sky130_fd_sc_hd__and3_1 _07112_ (.A(net298),
    .B(net297),
    .C(_04434_),
    .X(_06657_));
 sky130_fd_sc_hd__nand2_2 _07113_ (.A(net298),
    .B(_06656_),
    .Y(_06658_));
 sky130_fd_sc_hd__and3_1 _07114_ (.A(net298),
    .B(_06655_),
    .C(_06656_),
    .X(_06659_));
 sky130_fd_sc_hd__nand2_1 _07115_ (.A(_06655_),
    .B(_06657_),
    .Y(_06660_));
 sky130_fd_sc_hd__nor2_4 _07116_ (.A(net255),
    .B(_06659_),
    .Y(_06661_));
 sky130_fd_sc_hd__nand2_1 _07117_ (.A(net249),
    .B(_06660_),
    .Y(_06662_));
 sky130_fd_sc_hd__nor2_8 _07118_ (.A(div_complete),
    .B(_06661_),
    .Y(busy));
 sky130_fd_sc_hd__and4b_1 _07119_ (.A_N(instruction[2]),
    .B(instruction[1]),
    .C(pred_val),
    .D(instruction[0]),
    .X(_06663_));
 sky130_fd_sc_hd__and2_4 _07120_ (.A(instruction[11]),
    .B(_06663_),
    .X(dest_pred[0]));
 sky130_fd_sc_hd__and2_4 _07121_ (.A(instruction[12]),
    .B(_06663_),
    .X(dest_pred[1]));
 sky130_fd_sc_hd__and2_4 _07122_ (.A(instruction[13]),
    .B(_06663_),
    .X(dest_pred[2]));
 sky130_fd_sc_hd__or2_2 _07123_ (.A(_04723_),
    .B(_06655_),
    .X(_06664_));
 sky130_fd_sc_hd__and2_4 _07124_ (.A(instruction[11]),
    .B(_06664_),
    .X(dest_idx[0]));
 sky130_fd_sc_hd__and2_4 _07125_ (.A(instruction[12]),
    .B(_06664_),
    .X(dest_idx[1]));
 sky130_fd_sc_hd__and2_4 _07126_ (.A(instruction[13]),
    .B(_06664_),
    .X(dest_idx[2]));
 sky130_fd_sc_hd__and2_4 _07127_ (.A(instruction[14]),
    .B(_06664_),
    .X(dest_idx[3]));
 sky130_fd_sc_hd__and2_4 _07128_ (.A(instruction[15]),
    .B(_06664_),
    .X(dest_idx[4]));
 sky130_fd_sc_hd__and2_4 _07129_ (.A(instruction[16]),
    .B(_06664_),
    .X(dest_idx[5]));
 sky130_fd_sc_hd__mux2_8 _07130_ (.A0(instruction[25]),
    .A1(instruction[18]),
    .S(_04652_),
    .X(reg2_idx[0]));
 sky130_fd_sc_hd__mux2_8 _07131_ (.A0(instruction[26]),
    .A1(instruction[19]),
    .S(_04652_),
    .X(reg2_idx[1]));
 sky130_fd_sc_hd__mux2_8 _07132_ (.A0(instruction[27]),
    .A1(instruction[20]),
    .S(_04652_),
    .X(reg2_idx[2]));
 sky130_fd_sc_hd__mux2_8 _07133_ (.A0(instruction[28]),
    .A1(instruction[21]),
    .S(_04652_),
    .X(reg2_idx[3]));
 sky130_fd_sc_hd__mux2_8 _07134_ (.A0(instruction[29]),
    .A1(instruction[22]),
    .S(_04652_),
    .X(reg2_idx[4]));
 sky130_fd_sc_hd__mux2_8 _07135_ (.A0(instruction[30]),
    .A1(instruction[23]),
    .S(_04652_),
    .X(reg2_idx[5]));
 sky130_fd_sc_hd__or3_2 _07136_ (.A(_04423_),
    .B(net298),
    .C(net297),
    .X(_06665_));
 sky130_fd_sc_hd__nor2_2 _07137_ (.A(instruction[5]),
    .B(_06665_),
    .Y(_06666_));
 sky130_fd_sc_hd__or2_4 _07138_ (.A(instruction[5]),
    .B(_06665_),
    .X(_06667_));
 sky130_fd_sc_hd__or2_1 _07139_ (.A(net297),
    .B(instruction[5]),
    .X(_06668_));
 sky130_fd_sc_hd__nand2_1 _07140_ (.A(_04423_),
    .B(net298),
    .Y(_06669_));
 sky130_fd_sc_hd__or2_2 _07141_ (.A(_06668_),
    .B(_06669_),
    .X(_06670_));
 sky130_fd_sc_hd__a31o_1 _07142_ (.A1(instruction[17]),
    .A2(_06667_),
    .A3(_06670_),
    .B1(net269),
    .X(_06671_));
 sky130_fd_sc_hd__nor2_1 _07143_ (.A(is_load),
    .B(_06656_),
    .Y(_06672_));
 sky130_fd_sc_hd__o211a_1 _07144_ (.A1(instruction[40]),
    .A2(_04819_),
    .B1(_06671_),
    .C1(_06672_),
    .X(_06673_));
 sky130_fd_sc_hd__a32o_2 _07145_ (.A1(instruction[24]),
    .A2(net296),
    .A3(is_load),
    .B1(_04862_),
    .B2(_06673_),
    .X(_06674_));
 sky130_fd_sc_hd__nand2_8 _07146_ (.A(net240),
    .B(_06674_),
    .Y(dest_mask[0]));
 sky130_fd_sc_hd__a22o_2 _07147_ (.A1(net296),
    .A2(is_load),
    .B1(net247),
    .B2(_06673_),
    .X(_06675_));
 sky130_fd_sc_hd__nand2_8 _07148_ (.A(net240),
    .B(_06675_),
    .Y(dest_mask[1]));
 sky130_fd_sc_hd__or2_2 _07149_ (.A(net297),
    .B(_04434_),
    .X(_06676_));
 sky130_fd_sc_hd__and4b_4 _07150_ (.A_N(net297),
    .B(instruction[5]),
    .C(net296),
    .D(_06636_),
    .X(_06677_));
 sky130_fd_sc_hd__or4_1 _07151_ (.A(instruction[3]),
    .B(net298),
    .C(net284),
    .D(_06676_),
    .X(_06678_));
 sky130_fd_sc_hd__a31o_2 _07152_ (.A1(net298),
    .A2(net297),
    .A3(instruction[5]),
    .B1(_06677_),
    .X(_06679_));
 sky130_fd_sc_hd__and2_1 _07153_ (.A(net296),
    .B(_04949_),
    .X(_06680_));
 sky130_fd_sc_hd__nand2_4 _07154_ (.A(net296),
    .B(_04949_),
    .Y(_06681_));
 sky130_fd_sc_hd__and2_1 _07155_ (.A(reg1_val[31]),
    .B(net293),
    .X(_06682_));
 sky130_fd_sc_hd__nand2_2 _07156_ (.A(reg1_val[31]),
    .B(net293),
    .Y(_06683_));
 sky130_fd_sc_hd__or3_2 _07157_ (.A(net292),
    .B(net289),
    .C(reg1_val[2]),
    .X(_06684_));
 sky130_fd_sc_hd__or4_2 _07158_ (.A(net292),
    .B(net289),
    .C(reg1_val[2]),
    .D(reg1_val[3]),
    .X(_06685_));
 sky130_fd_sc_hd__nor2_1 _07159_ (.A(reg1_val[4]),
    .B(_06685_),
    .Y(_06686_));
 sky130_fd_sc_hd__xnor2_2 _07160_ (.A(reg1_val[5]),
    .B(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__or2_1 _07161_ (.A(reg1_val[5]),
    .B(net260),
    .X(_06688_));
 sky130_fd_sc_hd__o21ai_2 _07162_ (.A1(net259),
    .A2(_06687_),
    .B1(_06688_),
    .Y(_06689_));
 sky130_fd_sc_hd__o21a_1 _07163_ (.A1(net259),
    .A2(_06687_),
    .B1(_06688_),
    .X(_06690_));
 sky130_fd_sc_hd__xor2_2 _07164_ (.A(reg1_val[3]),
    .B(_06684_),
    .X(_06691_));
 sky130_fd_sc_hd__or2_2 _07165_ (.A(reg1_val[3]),
    .B(net260),
    .X(_06692_));
 sky130_fd_sc_hd__o21ai_4 _07166_ (.A1(net259),
    .A2(_06691_),
    .B1(_06692_),
    .Y(_06693_));
 sky130_fd_sc_hd__o21a_4 _07167_ (.A1(net259),
    .A2(_06691_),
    .B1(_06692_),
    .X(_06694_));
 sky130_fd_sc_hd__xor2_1 _07168_ (.A(reg1_val[4]),
    .B(_06685_),
    .X(_06695_));
 sky130_fd_sc_hd__mux2_1 _07169_ (.A0(reg1_val[4]),
    .A1(_06695_),
    .S(net260),
    .X(_06696_));
 sky130_fd_sc_hd__nor2_2 _07170_ (.A(_06694_),
    .B(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__or2_1 _07171_ (.A(_06694_),
    .B(_06696_),
    .X(_06698_));
 sky130_fd_sc_hd__nand2_1 _07172_ (.A(_06694_),
    .B(_06696_),
    .Y(_06699_));
 sky130_fd_sc_hd__nor2_2 _07173_ (.A(net179),
    .B(_06699_),
    .Y(_06700_));
 sky130_fd_sc_hd__a21oi_4 _07174_ (.A1(net179),
    .A2(_06697_),
    .B1(_06700_),
    .Y(_06701_));
 sky130_fd_sc_hd__a21o_4 _07175_ (.A1(net179),
    .A2(_06697_),
    .B1(_06700_),
    .X(_06702_));
 sky130_fd_sc_hd__and2_4 _07176_ (.A(net293),
    .B(_04917_),
    .X(_06703_));
 sky130_fd_sc_hd__nand2_1 _07177_ (.A(net293),
    .B(_04917_),
    .Y(_06704_));
 sky130_fd_sc_hd__or2_1 _07178_ (.A(_06165_),
    .B(_06240_),
    .X(_06705_));
 sky130_fd_sc_hd__and4_4 _07179_ (.A(_06553_),
    .B(_06560_),
    .C(net214),
    .D(net211),
    .X(_06706_));
 sky130_fd_sc_hd__and4bb_4 _07180_ (.A_N(_06523_),
    .B_N(_06529_),
    .C(_06538_),
    .D(_06547_),
    .X(_06707_));
 sky130_fd_sc_hd__and2_1 _07181_ (.A(_06706_),
    .B(_06707_),
    .X(_06708_));
 sky130_fd_sc_hd__nand2_2 _07182_ (.A(_06706_),
    .B(_06707_),
    .Y(_06709_));
 sky130_fd_sc_hd__nor2_1 _07183_ (.A(_06509_),
    .B(_06516_),
    .Y(_06710_));
 sky130_fd_sc_hd__nor4_1 _07184_ (.A(_06426_),
    .B(_06495_),
    .C(_06509_),
    .D(_06516_),
    .Y(_06711_));
 sky130_fd_sc_hd__and3_1 _07185_ (.A(_06706_),
    .B(_06707_),
    .C(_06711_),
    .X(_06712_));
 sky130_fd_sc_hd__and4_2 _07186_ (.A(_06363_),
    .B(_06706_),
    .C(_06707_),
    .D(net176),
    .X(_06713_));
 sky130_fd_sc_hd__and4b_2 _07187_ (.A_N(_06705_),
    .B(net176),
    .C(_06315_),
    .D(_06363_),
    .X(_06714_));
 sky130_fd_sc_hd__or4b_1 _07188_ (.A(_06309_),
    .B(_06357_),
    .C(_06705_),
    .D_N(net176),
    .X(_06715_));
 sky130_fd_sc_hd__nand2_1 _07189_ (.A(_06708_),
    .B(_06714_),
    .Y(_06716_));
 sky130_fd_sc_hd__nand2_1 _07190_ (.A(_06031_),
    .B(_06112_),
    .Y(_06717_));
 sky130_fd_sc_hd__and4_1 _07191_ (.A(_05874_),
    .B(_05940_),
    .C(_06031_),
    .D(_06112_),
    .X(_06718_));
 sky130_fd_sc_hd__and3_4 _07192_ (.A(_06708_),
    .B(_06714_),
    .C(_06718_),
    .X(_06719_));
 sky130_fd_sc_hd__or3b_4 _07193_ (.A(_06709_),
    .B(_06715_),
    .C_N(_06718_),
    .X(_06720_));
 sky130_fd_sc_hd__nor2_1 _07194_ (.A(_05731_),
    .B(net177),
    .Y(_06721_));
 sky130_fd_sc_hd__a211o_2 _07195_ (.A1(_05731_),
    .A2(_06719_),
    .B1(net177),
    .C1(_05807_),
    .X(_06722_));
 sky130_fd_sc_hd__a211o_2 _07196_ (.A1(_06703_),
    .A2(_06720_),
    .B1(_06721_),
    .C1(_05796_),
    .X(_06723_));
 sky130_fd_sc_hd__and2_1 _07197_ (.A(_06722_),
    .B(_06723_),
    .X(_06724_));
 sky130_fd_sc_hd__nand2_8 _07198_ (.A(_06722_),
    .B(_06723_),
    .Y(_06725_));
 sky130_fd_sc_hd__and2_4 _07199_ (.A(_06698_),
    .B(_06699_),
    .X(_06726_));
 sky130_fd_sc_hd__nand2_2 _07200_ (.A(_06698_),
    .B(_06699_),
    .Y(_06727_));
 sky130_fd_sc_hd__and2_2 _07201_ (.A(_05731_),
    .B(_05796_),
    .X(_06728_));
 sky130_fd_sc_hd__a21o_2 _07202_ (.A1(_06719_),
    .A2(_06728_),
    .B1(net177),
    .X(_06729_));
 sky130_fd_sc_hd__xnor2_4 _07203_ (.A(_05666_),
    .B(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__xnor2_2 _07204_ (.A(_05656_),
    .B(_06729_),
    .Y(_06731_));
 sky130_fd_sc_hd__o22a_1 _07205_ (.A1(net133),
    .A2(net56),
    .B1(net158),
    .B2(net53),
    .X(_06732_));
 sky130_fd_sc_hd__xnor2_2 _07206_ (.A(net179),
    .B(_06732_),
    .Y(_06733_));
 sky130_fd_sc_hd__xor2_1 _07207_ (.A(net292),
    .B(net289),
    .X(_06734_));
 sky130_fd_sc_hd__or2_1 _07208_ (.A(net259),
    .B(_06734_),
    .X(_06735_));
 sky130_fd_sc_hd__o21a_2 _07209_ (.A1(net289),
    .A2(net260),
    .B1(_06735_),
    .X(_06736_));
 sky130_fd_sc_hd__o21ai_4 _07210_ (.A1(net289),
    .A2(net260),
    .B1(_06735_),
    .Y(_06737_));
 sky130_fd_sc_hd__and3_1 _07211_ (.A(_05591_),
    .B(_05656_),
    .C(_06728_),
    .X(_06738_));
 sky130_fd_sc_hd__nand3_2 _07212_ (.A(_05591_),
    .B(_05656_),
    .C(_06728_),
    .Y(_06739_));
 sky130_fd_sc_hd__nand2_1 _07213_ (.A(_06719_),
    .B(_06738_),
    .Y(_06740_));
 sky130_fd_sc_hd__nor2_1 _07214_ (.A(_05308_),
    .B(_05493_),
    .Y(_06741_));
 sky130_fd_sc_hd__a31o_2 _07215_ (.A1(_06719_),
    .A2(_06738_),
    .A3(_06741_),
    .B1(net177),
    .X(_06742_));
 sky130_fd_sc_hd__xnor2_4 _07216_ (.A(_05395_),
    .B(_06742_),
    .Y(_00136_));
 sky130_fd_sc_hd__xnor2_2 _07217_ (.A(_05385_),
    .B(_06742_),
    .Y(_00137_));
 sky130_fd_sc_hd__nor2_8 _07218_ (.A(net292),
    .B(_04467_),
    .Y(_00138_));
 sky130_fd_sc_hd__nand2_1 _07219_ (.A(net285),
    .B(net289),
    .Y(_00139_));
 sky130_fd_sc_hd__a21oi_1 _07220_ (.A1(_06719_),
    .A2(_06738_),
    .B1(net177),
    .Y(_00140_));
 sky130_fd_sc_hd__nor2_1 _07221_ (.A(_05482_),
    .B(net177),
    .Y(_00141_));
 sky130_fd_sc_hd__a31o_2 _07222_ (.A1(_05482_),
    .A2(_06719_),
    .A3(_06738_),
    .B1(net177),
    .X(_00142_));
 sky130_fd_sc_hd__xnor2_2 _07223_ (.A(_05319_),
    .B(_00142_),
    .Y(_00143_));
 sky130_fd_sc_hd__xnor2_4 _07224_ (.A(_05308_),
    .B(_00142_),
    .Y(_00144_));
 sky130_fd_sc_hd__o22a_1 _07225_ (.A1(net285),
    .A2(net51),
    .B1(net236),
    .B2(net49),
    .X(_00145_));
 sky130_fd_sc_hd__xnor2_2 _07226_ (.A(net199),
    .B(_00145_),
    .Y(_00146_));
 sky130_fd_sc_hd__nand2_1 _07227_ (.A(_06733_),
    .B(_00146_),
    .Y(_00147_));
 sky130_fd_sc_hd__a31oi_4 _07228_ (.A1(_05656_),
    .A2(_06719_),
    .A3(_06728_),
    .B1(net177),
    .Y(_00148_));
 sky130_fd_sc_hd__xor2_2 _07229_ (.A(_05591_),
    .B(_00148_),
    .X(_00149_));
 sky130_fd_sc_hd__xnor2_4 _07230_ (.A(_05591_),
    .B(_00148_),
    .Y(_00150_));
 sky130_fd_sc_hd__o21ai_1 _07231_ (.A1(net292),
    .A2(net289),
    .B1(reg1_val[2]),
    .Y(_00151_));
 sky130_fd_sc_hd__and3_1 _07232_ (.A(net260),
    .B(_06684_),
    .C(_00151_),
    .X(_00152_));
 sky130_fd_sc_hd__a21o_1 _07233_ (.A1(reg1_val[2]),
    .A2(net259),
    .B1(_00152_),
    .X(_00153_));
 sky130_fd_sc_hd__nor2_4 _07234_ (.A(net199),
    .B(_00153_),
    .Y(_00154_));
 sky130_fd_sc_hd__and2_2 _07235_ (.A(net199),
    .B(_00153_),
    .X(_00155_));
 sky130_fd_sc_hd__and2_1 _07236_ (.A(net201),
    .B(_00155_),
    .X(_00156_));
 sky130_fd_sc_hd__a21oi_2 _07237_ (.A1(net200),
    .A2(_00154_),
    .B1(_00156_),
    .Y(_00157_));
 sky130_fd_sc_hd__mux2_8 _07238_ (.A0(_00154_),
    .A1(_00155_),
    .S(net201),
    .X(_00158_));
 sky130_fd_sc_hd__nor2_8 _07239_ (.A(_00154_),
    .B(_00155_),
    .Y(_00159_));
 sky130_fd_sc_hd__or2_2 _07240_ (.A(_00154_),
    .B(_00155_),
    .X(_00160_));
 sky130_fd_sc_hd__o2bb2a_4 _07241_ (.A1_N(_06740_),
    .A2_N(_00141_),
    .B1(_00140_),
    .B2(_05493_),
    .X(_00161_));
 sky130_fd_sc_hd__a2bb2o_1 _07242_ (.A1_N(_05493_),
    .A2_N(_00140_),
    .B1(_00141_),
    .B2(_06740_),
    .X(_00162_));
 sky130_fd_sc_hd__o22a_1 _07243_ (.A1(net47),
    .A2(net132),
    .B1(net157),
    .B2(net45),
    .X(_00163_));
 sky130_fd_sc_hd__xnor2_2 _07244_ (.A(net201),
    .B(_00163_),
    .Y(_00164_));
 sky130_fd_sc_hd__xnor2_2 _07245_ (.A(_06733_),
    .B(_00146_),
    .Y(_00165_));
 sky130_fd_sc_hd__o21ai_1 _07246_ (.A1(_00164_),
    .A2(_00165_),
    .B1(_00147_),
    .Y(_00166_));
 sky130_fd_sc_hd__o22a_1 _07247_ (.A1(net49),
    .A2(net157),
    .B1(net45),
    .B2(net132),
    .X(_00167_));
 sky130_fd_sc_hd__xnor2_1 _07248_ (.A(net201),
    .B(_00167_),
    .Y(_00168_));
 sky130_fd_sc_hd__o22a_1 _07249_ (.A1(net133),
    .A2(net53),
    .B1(net47),
    .B2(net158),
    .X(_00169_));
 sky130_fd_sc_hd__xnor2_2 _07250_ (.A(net179),
    .B(_00169_),
    .Y(_00170_));
 sky130_fd_sc_hd__nor2_1 _07251_ (.A(_04982_),
    .B(_06703_),
    .Y(_00171_));
 sky130_fd_sc_hd__or4_2 _07252_ (.A(_04993_),
    .B(_05308_),
    .C(_05395_),
    .D(_05493_),
    .X(_00172_));
 sky130_fd_sc_hd__nor3_4 _07253_ (.A(_06720_),
    .B(_06739_),
    .C(_00172_),
    .Y(_00173_));
 sky130_fd_sc_hd__or3_4 _07254_ (.A(_06720_),
    .B(_06739_),
    .C(_00172_),
    .X(_00174_));
 sky130_fd_sc_hd__a41o_1 _07255_ (.A1(_05385_),
    .A2(_06719_),
    .A3(_06738_),
    .A4(_06741_),
    .B1(_04982_),
    .X(_00175_));
 sky130_fd_sc_hd__a31oi_1 _07256_ (.A1(_06703_),
    .A2(_00174_),
    .A3(_00175_),
    .B1(_00171_),
    .Y(_00176_));
 sky130_fd_sc_hd__a31o_4 _07257_ (.A1(_06703_),
    .A2(_00174_),
    .A3(_00175_),
    .B1(_00171_),
    .X(_00177_));
 sky130_fd_sc_hd__o22a_1 _07258_ (.A1(net51),
    .A2(net236),
    .B1(net44),
    .B2(net286),
    .X(_00178_));
 sky130_fd_sc_hd__xnor2_2 _07259_ (.A(net199),
    .B(_00178_),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_1 _07260_ (.A(_00170_),
    .B(_00179_),
    .Y(_00180_));
 sky130_fd_sc_hd__xnor2_2 _07261_ (.A(_00170_),
    .B(_00179_),
    .Y(_00181_));
 sky130_fd_sc_hd__or2_1 _07262_ (.A(_00168_),
    .B(_00181_),
    .X(_00182_));
 sky130_fd_sc_hd__nand2_1 _07263_ (.A(_00168_),
    .B(_00181_),
    .Y(_00183_));
 sky130_fd_sc_hd__xnor2_1 _07264_ (.A(_00168_),
    .B(_00181_),
    .Y(_00184_));
 sky130_fd_sc_hd__or4_4 _07265_ (.A(reg1_val[4]),
    .B(reg1_val[5]),
    .C(reg1_val[6]),
    .D(_06685_),
    .X(_00185_));
 sky130_fd_sc_hd__xor2_2 _07266_ (.A(net287),
    .B(_00185_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_2 _07267_ (.A0(net287),
    .A1(_00186_),
    .S(net260),
    .X(_00187_));
 sky130_fd_sc_hd__inv_6 _07268_ (.A(net174),
    .Y(_00188_));
 sky130_fd_sc_hd__o31ai_1 _07269_ (.A1(reg1_val[4]),
    .A2(reg1_val[5]),
    .A3(_06685_),
    .B1(reg1_val[6]),
    .Y(_00189_));
 sky130_fd_sc_hd__and2_1 _07270_ (.A(_00185_),
    .B(_00189_),
    .X(_00190_));
 sky130_fd_sc_hd__or2_1 _07271_ (.A(reg1_val[6]),
    .B(net260),
    .X(_00191_));
 sky130_fd_sc_hd__o21ai_2 _07272_ (.A1(net259),
    .A2(_00190_),
    .B1(_00191_),
    .Y(_00192_));
 sky130_fd_sc_hd__nand2_1 _07273_ (.A(net181),
    .B(_00192_),
    .Y(_00193_));
 sky130_fd_sc_hd__or2_1 _07274_ (.A(net181),
    .B(_00192_),
    .X(_00194_));
 sky130_fd_sc_hd__nor2_1 _07275_ (.A(net174),
    .B(_00194_),
    .Y(_00195_));
 sky130_fd_sc_hd__o21ba_2 _07276_ (.A1(_00188_),
    .A2(_00193_),
    .B1_N(_00195_),
    .X(_00196_));
 sky130_fd_sc_hd__o21bai_1 _07277_ (.A1(_00188_),
    .A2(_00193_),
    .B1_N(_00195_),
    .Y(_00197_));
 sky130_fd_sc_hd__o31a_4 _07278_ (.A1(_06709_),
    .A2(_06715_),
    .A3(_06717_),
    .B1(_06703_),
    .X(_00198_));
 sky130_fd_sc_hd__nor2_1 _07279_ (.A(_05940_),
    .B(net178),
    .Y(_00199_));
 sky130_fd_sc_hd__o21ai_4 _07280_ (.A1(_00198_),
    .A2(_00199_),
    .B1(_05874_),
    .Y(_00200_));
 sky130_fd_sc_hd__or3_4 _07281_ (.A(_05874_),
    .B(_00198_),
    .C(_00199_),
    .X(_00201_));
 sky130_fd_sc_hd__and2_4 _07282_ (.A(_00200_),
    .B(_00201_),
    .X(_00202_));
 sky130_fd_sc_hd__nand2_8 _07283_ (.A(_00200_),
    .B(_00201_),
    .Y(_00203_));
 sky130_fd_sc_hd__and2_1 _07284_ (.A(_00193_),
    .B(_00194_),
    .X(_00204_));
 sky130_fd_sc_hd__nand2_2 _07285_ (.A(_00193_),
    .B(_00194_),
    .Y(_00205_));
 sky130_fd_sc_hd__o21a_2 _07286_ (.A1(net177),
    .A2(_06719_),
    .B1(_05731_),
    .X(_00206_));
 sky130_fd_sc_hd__and2_2 _07287_ (.A(_06720_),
    .B(_06721_),
    .X(_00207_));
 sky130_fd_sc_hd__nor2_8 _07288_ (.A(_00206_),
    .B(_00207_),
    .Y(_00208_));
 sky130_fd_sc_hd__or2_1 _07289_ (.A(_00206_),
    .B(_00207_),
    .X(_00209_));
 sky130_fd_sc_hd__o22a_1 _07290_ (.A1(net105),
    .A2(net42),
    .B1(net131),
    .B2(net40),
    .X(_00210_));
 sky130_fd_sc_hd__xnor2_1 _07291_ (.A(_00188_),
    .B(_00210_),
    .Y(_00211_));
 sky130_fd_sc_hd__or3_2 _07292_ (.A(net287),
    .B(reg1_val[8]),
    .C(_00185_),
    .X(_00212_));
 sky130_fd_sc_hd__or2_2 _07293_ (.A(reg1_val[8]),
    .B(reg1_val[9]),
    .X(_00213_));
 sky130_fd_sc_hd__xor2_2 _07294_ (.A(reg1_val[9]),
    .B(_00212_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _07295_ (.A0(reg1_val[9]),
    .A1(_00214_),
    .S(net260),
    .X(_00215_));
 sky130_fd_sc_hd__a21oi_1 _07296_ (.A1(_06708_),
    .A2(_06714_),
    .B1(net177),
    .Y(_00216_));
 sky130_fd_sc_hd__nor2_1 _07297_ (.A(_06112_),
    .B(net177),
    .Y(_00217_));
 sky130_fd_sc_hd__a31o_4 _07298_ (.A1(_06112_),
    .A2(_06708_),
    .A3(_06714_),
    .B1(net177),
    .X(_00218_));
 sky130_fd_sc_hd__xnor2_4 _07299_ (.A(_06031_),
    .B(_00218_),
    .Y(_00219_));
 sky130_fd_sc_hd__xnor2_4 _07300_ (.A(_06041_),
    .B(_00218_),
    .Y(_00220_));
 sky130_fd_sc_hd__and2_1 _07301_ (.A(reg1_val[8]),
    .B(net259),
    .X(_00221_));
 sky130_fd_sc_hd__o21ai_1 _07302_ (.A1(net287),
    .A2(_00185_),
    .B1(reg1_val[8]),
    .Y(_00222_));
 sky130_fd_sc_hd__a31o_1 _07303_ (.A1(net260),
    .A2(_00212_),
    .A3(_00222_),
    .B1(_00221_),
    .X(_00223_));
 sky130_fd_sc_hd__nor2_2 _07304_ (.A(net174),
    .B(_00223_),
    .Y(_00224_));
 sky130_fd_sc_hd__and2_1 _07305_ (.A(net174),
    .B(_00223_),
    .X(_00225_));
 sky130_fd_sc_hd__and2b_1 _07306_ (.A_N(net155),
    .B(_00225_),
    .X(_00226_));
 sky130_fd_sc_hd__a21oi_4 _07307_ (.A1(net155),
    .A2(_00224_),
    .B1(_00226_),
    .Y(_00227_));
 sky130_fd_sc_hd__mux2_2 _07308_ (.A0(_00225_),
    .A1(_00224_),
    .S(net155),
    .X(_00228_));
 sky130_fd_sc_hd__xnor2_4 _07309_ (.A(_05940_),
    .B(_00198_),
    .Y(_00229_));
 sky130_fd_sc_hd__xnor2_4 _07310_ (.A(_05949_),
    .B(_00198_),
    .Y(_00230_));
 sky130_fd_sc_hd__nor2_2 _07311_ (.A(_00224_),
    .B(_00225_),
    .Y(_00231_));
 sky130_fd_sc_hd__or2_2 _07312_ (.A(_00224_),
    .B(_00225_),
    .X(_00232_));
 sky130_fd_sc_hd__a22o_1 _07313_ (.A1(_00220_),
    .A2(net129),
    .B1(_00229_),
    .B2(net127),
    .X(_00233_));
 sky130_fd_sc_hd__xnor2_1 _07314_ (.A(net154),
    .B(_00233_),
    .Y(_00234_));
 sky130_fd_sc_hd__nor2_1 _07315_ (.A(_00211_),
    .B(_00234_),
    .Y(_00235_));
 sky130_fd_sc_hd__xnor2_1 _07316_ (.A(_00166_),
    .B(_00184_),
    .Y(_00236_));
 sky130_fd_sc_hd__a32o_2 _07317_ (.A1(_00166_),
    .A2(_00182_),
    .A3(_00183_),
    .B1(_00235_),
    .B2(_00236_),
    .X(_00237_));
 sky130_fd_sc_hd__nand2_2 _07318_ (.A(_04554_),
    .B(net259),
    .Y(_00238_));
 sky130_fd_sc_hd__nor4_4 _07319_ (.A(net287),
    .B(reg1_val[10]),
    .C(_00185_),
    .D(_00213_),
    .Y(_00239_));
 sky130_fd_sc_hd__or4_2 _07320_ (.A(net287),
    .B(reg1_val[10]),
    .C(_00185_),
    .D(_00213_),
    .X(_00240_));
 sky130_fd_sc_hd__or3_1 _07321_ (.A(net290),
    .B(reg1_val[12]),
    .C(_00240_),
    .X(_00241_));
 sky130_fd_sc_hd__nor2_1 _07322_ (.A(reg1_val[12]),
    .B(reg1_val[13]),
    .Y(_00242_));
 sky130_fd_sc_hd__or2_1 _07323_ (.A(reg1_val[12]),
    .B(reg1_val[13]),
    .X(_00243_));
 sky130_fd_sc_hd__and3_1 _07324_ (.A(_04478_),
    .B(_00239_),
    .C(_00242_),
    .X(_00244_));
 sky130_fd_sc_hd__or4_2 _07325_ (.A(net290),
    .B(reg1_val[14]),
    .C(_00240_),
    .D(_00243_),
    .X(_00245_));
 sky130_fd_sc_hd__or2_1 _07326_ (.A(reg1_val[14]),
    .B(reg1_val[15]),
    .X(_00246_));
 sky130_fd_sc_hd__nor4_2 _07327_ (.A(net290),
    .B(_00240_),
    .C(_00243_),
    .D(_00246_),
    .Y(_00247_));
 sky130_fd_sc_hd__or4_4 _07328_ (.A(net290),
    .B(_00240_),
    .C(_00243_),
    .D(_00246_),
    .X(_00248_));
 sky130_fd_sc_hd__or2_4 _07329_ (.A(reg1_val[16]),
    .B(reg1_val[17]),
    .X(_00249_));
 sky130_fd_sc_hd__nor3_2 _07330_ (.A(reg1_val[18]),
    .B(reg1_val[19]),
    .C(_00249_),
    .Y(_00250_));
 sky130_fd_sc_hd__or3_4 _07331_ (.A(reg1_val[18]),
    .B(reg1_val[19]),
    .C(_00249_),
    .X(_00251_));
 sky130_fd_sc_hd__nor2_1 _07332_ (.A(reg1_val[20]),
    .B(reg1_val[21]),
    .Y(_00252_));
 sky130_fd_sc_hd__or2_1 _07333_ (.A(reg1_val[20]),
    .B(reg1_val[21]),
    .X(_00253_));
 sky130_fd_sc_hd__and4_2 _07334_ (.A(_04543_),
    .B(_04554_),
    .C(_00250_),
    .D(_00252_),
    .X(_00254_));
 sky130_fd_sc_hd__or4_4 _07335_ (.A(reg1_val[22]),
    .B(reg1_val[23]),
    .C(_00251_),
    .D(_00253_),
    .X(_00255_));
 sky130_fd_sc_hd__nand2_1 _07336_ (.A(net173),
    .B(_00254_),
    .Y(_00256_));
 sky130_fd_sc_hd__nand2_1 _07337_ (.A(net173),
    .B(_00250_),
    .Y(_00257_));
 sky130_fd_sc_hd__or3_1 _07338_ (.A(_00248_),
    .B(_00251_),
    .C(_00253_),
    .X(_00258_));
 sky130_fd_sc_hd__or4_1 _07339_ (.A(reg1_val[22]),
    .B(_00248_),
    .C(_00251_),
    .D(_00253_),
    .X(_00259_));
 sky130_fd_sc_hd__a41o_1 _07340_ (.A1(_04543_),
    .A2(net173),
    .A3(_00250_),
    .A4(_00252_),
    .B1(_04554_),
    .X(_00260_));
 sky130_fd_sc_hd__a21o_2 _07341_ (.A1(_00256_),
    .A2(_00260_),
    .B1(net258),
    .X(_00261_));
 sky130_fd_sc_hd__and2_4 _07342_ (.A(_00238_),
    .B(_00261_),
    .X(_00262_));
 sky130_fd_sc_hd__nand2_2 _07343_ (.A(_00238_),
    .B(_00261_),
    .Y(_00263_));
 sky130_fd_sc_hd__o21a_2 _07344_ (.A1(net178),
    .A2(_06706_),
    .B1(_06547_),
    .X(_00264_));
 sky130_fd_sc_hd__and3b_2 _07345_ (.A_N(_06706_),
    .B(_06703_),
    .C(net222),
    .X(_00265_));
 sky130_fd_sc_hd__nor2_8 _07346_ (.A(_00264_),
    .B(_00265_),
    .Y(_00266_));
 sky130_fd_sc_hd__or2_4 _07347_ (.A(_00264_),
    .B(_00265_),
    .X(_00267_));
 sky130_fd_sc_hd__nand2_4 _07348_ (.A(_04532_),
    .B(net258),
    .Y(_00268_));
 sky130_fd_sc_hd__or3_1 _07349_ (.A(reg1_val[20]),
    .B(_00248_),
    .C(_00251_),
    .X(_00269_));
 sky130_fd_sc_hd__a31o_1 _07350_ (.A1(_04521_),
    .A2(net173),
    .A3(_00250_),
    .B1(_04532_),
    .X(_00270_));
 sky130_fd_sc_hd__and2_1 _07351_ (.A(_00258_),
    .B(_00270_),
    .X(_00271_));
 sky130_fd_sc_hd__a21o_2 _07352_ (.A1(_00258_),
    .A2(_00270_),
    .B1(net258),
    .X(_00272_));
 sky130_fd_sc_hd__and2_4 _07353_ (.A(_00268_),
    .B(_00272_),
    .X(_00273_));
 sky130_fd_sc_hd__nand2_8 _07354_ (.A(_00268_),
    .B(_00272_),
    .Y(_00274_));
 sky130_fd_sc_hd__a31o_1 _07355_ (.A1(net173),
    .A2(_00250_),
    .A3(_00252_),
    .B1(_04543_),
    .X(_00275_));
 sky130_fd_sc_hd__a21o_1 _07356_ (.A1(_00259_),
    .A2(_00275_),
    .B1(net258),
    .X(_00276_));
 sky130_fd_sc_hd__nand2_1 _07357_ (.A(_04543_),
    .B(net259),
    .Y(_00277_));
 sky130_fd_sc_hd__and2_1 _07358_ (.A(_00276_),
    .B(_00277_),
    .X(_00278_));
 sky130_fd_sc_hd__a22o_1 _07359_ (.A1(_00268_),
    .A2(_00272_),
    .B1(_00276_),
    .B2(_00277_),
    .X(_00279_));
 sky130_fd_sc_hd__nand4_2 _07360_ (.A(_00268_),
    .B(_00272_),
    .C(_00276_),
    .D(_00277_),
    .Y(_00280_));
 sky130_fd_sc_hd__nor2_1 _07361_ (.A(net98),
    .B(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__mux2_1 _07362_ (.A0(_00279_),
    .A1(_00280_),
    .S(_00263_),
    .X(_00282_));
 sky130_fd_sc_hd__or3b_1 _07363_ (.A(net283),
    .B(_06547_),
    .C_N(_04917_),
    .X(_00283_));
 sky130_fd_sc_hd__a211o_2 _07364_ (.A1(_06547_),
    .A2(_06706_),
    .B1(net178),
    .C1(_06539_),
    .X(_00284_));
 sky130_fd_sc_hd__o211ai_4 _07365_ (.A1(net178),
    .A2(_06706_),
    .B1(_00283_),
    .C1(_06539_),
    .Y(_00285_));
 sky130_fd_sc_hd__and2_4 _07366_ (.A(_00284_),
    .B(_00285_),
    .X(_00286_));
 sky130_fd_sc_hd__nand2_8 _07367_ (.A(_00284_),
    .B(_00285_),
    .Y(_00287_));
 sky130_fd_sc_hd__nand2_2 _07368_ (.A(_00279_),
    .B(_00280_),
    .Y(_00288_));
 sky130_fd_sc_hd__o22a_1 _07369_ (.A1(net125),
    .A2(net39),
    .B1(_00286_),
    .B2(net37),
    .X(_00289_));
 sky130_fd_sc_hd__xnor2_1 _07370_ (.A(net99),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__or2_2 _07371_ (.A(reg1_val[27]),
    .B(net261),
    .X(_00291_));
 sky130_fd_sc_hd__nor2_1 _07372_ (.A(reg1_val[24]),
    .B(reg1_val[25]),
    .Y(_00292_));
 sky130_fd_sc_hd__or2_2 _07373_ (.A(reg1_val[24]),
    .B(reg1_val[25]),
    .X(_00293_));
 sky130_fd_sc_hd__or3_4 _07374_ (.A(reg1_val[26]),
    .B(reg1_val[27]),
    .C(_00293_),
    .X(_00294_));
 sky130_fd_sc_hd__inv_2 _07375_ (.A(_00294_),
    .Y(_00295_));
 sky130_fd_sc_hd__and3_1 _07376_ (.A(net173),
    .B(_00254_),
    .C(_00295_),
    .X(_00296_));
 sky130_fd_sc_hd__and3_1 _07377_ (.A(net173),
    .B(_00254_),
    .C(_00292_),
    .X(_00297_));
 sky130_fd_sc_hd__or4_1 _07378_ (.A(reg1_val[26]),
    .B(_00248_),
    .C(_00255_),
    .D(_00293_),
    .X(_00298_));
 sky130_fd_sc_hd__o41a_1 _07379_ (.A1(reg1_val[26]),
    .A2(_00248_),
    .A3(_00255_),
    .A4(_00293_),
    .B1(reg1_val[27]),
    .X(_00299_));
 sky130_fd_sc_hd__o21ai_4 _07380_ (.A1(_00296_),
    .A2(_00299_),
    .B1(net261),
    .Y(_00300_));
 sky130_fd_sc_hd__and2_1 _07381_ (.A(_00291_),
    .B(_00300_),
    .X(_00301_));
 sky130_fd_sc_hd__nand2_4 _07382_ (.A(_00291_),
    .B(_00300_),
    .Y(_00302_));
 sky130_fd_sc_hd__or2_2 _07383_ (.A(reg1_val[25]),
    .B(net261),
    .X(_00303_));
 sky130_fd_sc_hd__or3_1 _07384_ (.A(reg1_val[24]),
    .B(_00248_),
    .C(_00255_),
    .X(_00304_));
 sky130_fd_sc_hd__o31a_1 _07385_ (.A1(reg1_val[24]),
    .A2(_00248_),
    .A3(_00255_),
    .B1(reg1_val[25]),
    .X(_00305_));
 sky130_fd_sc_hd__nor2_1 _07386_ (.A(_00297_),
    .B(_00305_),
    .Y(_00306_));
 sky130_fd_sc_hd__o21ai_4 _07387_ (.A1(_00297_),
    .A2(_00305_),
    .B1(net261),
    .Y(_00307_));
 sky130_fd_sc_hd__and2_2 _07388_ (.A(_00303_),
    .B(_00307_),
    .X(_00308_));
 sky130_fd_sc_hd__nand2_4 _07389_ (.A(_00303_),
    .B(_00307_),
    .Y(_00309_));
 sky130_fd_sc_hd__a31o_1 _07390_ (.A1(net173),
    .A2(_00254_),
    .A3(_00292_),
    .B1(_04576_),
    .X(_00310_));
 sky130_fd_sc_hd__a21o_1 _07391_ (.A1(_00298_),
    .A2(_00310_),
    .B1(_06683_),
    .X(_00311_));
 sky130_fd_sc_hd__nand2_1 _07392_ (.A(_04576_),
    .B(net259),
    .Y(_00312_));
 sky130_fd_sc_hd__and2_1 _07393_ (.A(_00311_),
    .B(_00312_),
    .X(_00313_));
 sky130_fd_sc_hd__a22o_1 _07394_ (.A1(_00303_),
    .A2(_00307_),
    .B1(_00311_),
    .B2(_00312_),
    .X(_00314_));
 sky130_fd_sc_hd__nand4_2 _07395_ (.A(_00303_),
    .B(_00307_),
    .C(_00311_),
    .D(_00312_),
    .Y(_00315_));
 sky130_fd_sc_hd__nor2_1 _07396_ (.A(net93),
    .B(_00315_),
    .Y(_00316_));
 sky130_fd_sc_hd__mux2_1 _07397_ (.A0(_00314_),
    .A1(_00315_),
    .S(_00302_),
    .X(_00317_));
 sky130_fd_sc_hd__and3_4 _07398_ (.A(net293),
    .B(_04917_),
    .C(net206),
    .X(_00318_));
 sky130_fd_sc_hd__xnor2_4 _07399_ (.A(net214),
    .B(_00318_),
    .Y(_00319_));
 sky130_fd_sc_hd__xnor2_4 _07400_ (.A(_06569_),
    .B(_00318_),
    .Y(_00320_));
 sky130_fd_sc_hd__nand2_1 _07401_ (.A(_00314_),
    .B(_00315_),
    .Y(_00321_));
 sky130_fd_sc_hd__o22a_1 _07402_ (.A1(net212),
    .A2(net35),
    .B1(net152),
    .B2(net33),
    .X(_00322_));
 sky130_fd_sc_hd__xnor2_1 _07403_ (.A(net95),
    .B(_00322_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _07404_ (.A(_00290_),
    .B(_00323_),
    .Y(_00324_));
 sky130_fd_sc_hd__o211a_4 _07405_ (.A1(_06569_),
    .A2(net206),
    .B1(net293),
    .C1(_04917_),
    .X(_00325_));
 sky130_fd_sc_hd__xnor2_4 _07406_ (.A(net216),
    .B(_00325_),
    .Y(_00326_));
 sky130_fd_sc_hd__xnor2_4 _07407_ (.A(_06560_),
    .B(_00325_),
    .Y(_00327_));
 sky130_fd_sc_hd__a21o_1 _07408_ (.A1(net173),
    .A2(_00254_),
    .B1(_04565_),
    .X(_00328_));
 sky130_fd_sc_hd__a21o_1 _07409_ (.A1(_00304_),
    .A2(_00328_),
    .B1(net258),
    .X(_00329_));
 sky130_fd_sc_hd__nand2_1 _07410_ (.A(_04565_),
    .B(net259),
    .Y(_00330_));
 sky130_fd_sc_hd__and2_1 _07411_ (.A(_00329_),
    .B(_00330_),
    .X(_00331_));
 sky130_fd_sc_hd__nor2_1 _07412_ (.A(net98),
    .B(_00331_),
    .Y(_00332_));
 sky130_fd_sc_hd__a22o_1 _07413_ (.A1(_00238_),
    .A2(_00261_),
    .B1(_00329_),
    .B2(_00330_),
    .X(_00333_));
 sky130_fd_sc_hd__nand4_4 _07414_ (.A(_00238_),
    .B(_00261_),
    .C(_00329_),
    .D(_00330_),
    .Y(_00334_));
 sky130_fd_sc_hd__nor2_1 _07415_ (.A(net92),
    .B(_00334_),
    .Y(_00335_));
 sky130_fd_sc_hd__mux2_2 _07416_ (.A0(_00333_),
    .A1(_00334_),
    .S(_00309_),
    .X(_00336_));
 sky130_fd_sc_hd__a21o_1 _07417_ (.A1(net92),
    .A2(_00332_),
    .B1(_00335_),
    .X(_00337_));
 sky130_fd_sc_hd__o311a_4 _07418_ (.A1(net216),
    .A2(_06569_),
    .A3(net206),
    .B1(_04917_),
    .C1(net293),
    .X(_00338_));
 sky130_fd_sc_hd__xnor2_4 _07419_ (.A(_06554_),
    .B(_00338_),
    .Y(_00339_));
 sky130_fd_sc_hd__xnor2_4 _07420_ (.A(_06553_),
    .B(_00338_),
    .Y(_00340_));
 sky130_fd_sc_hd__and2_2 _07421_ (.A(_00333_),
    .B(_00334_),
    .X(_00341_));
 sky130_fd_sc_hd__nand2_2 _07422_ (.A(_00333_),
    .B(_00334_),
    .Y(_00342_));
 sky130_fd_sc_hd__a22o_1 _07423_ (.A1(net150),
    .A2(net14),
    .B1(net148),
    .B2(net30),
    .X(_00343_));
 sky130_fd_sc_hd__xnor2_1 _07424_ (.A(net92),
    .B(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__or2_1 _07425_ (.A(_00290_),
    .B(_00323_),
    .X(_00345_));
 sky130_fd_sc_hd__nand2_1 _07426_ (.A(_00324_),
    .B(_00345_),
    .Y(_00346_));
 sky130_fd_sc_hd__or2_1 _07427_ (.A(_00344_),
    .B(_00346_),
    .X(_00347_));
 sky130_fd_sc_hd__nor2_1 _07428_ (.A(reg1_val[19]),
    .B(net261),
    .Y(_00348_));
 sky130_fd_sc_hd__inv_2 _07429_ (.A(_00348_),
    .Y(_00349_));
 sky130_fd_sc_hd__or3_1 _07430_ (.A(reg1_val[18]),
    .B(_00248_),
    .C(_00249_),
    .X(_00350_));
 sky130_fd_sc_hd__o31ai_4 _07431_ (.A1(reg1_val[18]),
    .A2(_00248_),
    .A3(_00249_),
    .B1(reg1_val[19]),
    .Y(_00351_));
 sky130_fd_sc_hd__a21o_1 _07432_ (.A1(_00257_),
    .A2(_00351_),
    .B1(net258),
    .X(_00352_));
 sky130_fd_sc_hd__and2_1 _07433_ (.A(_00349_),
    .B(_00352_),
    .X(_00353_));
 sky130_fd_sc_hd__or2_2 _07434_ (.A(reg1_val[17]),
    .B(net261),
    .X(_00354_));
 sky130_fd_sc_hd__or2_1 _07435_ (.A(_00248_),
    .B(_00249_),
    .X(_00355_));
 sky130_fd_sc_hd__o21ai_1 _07436_ (.A1(reg1_val[16]),
    .A2(_00248_),
    .B1(reg1_val[17]),
    .Y(_00356_));
 sky130_fd_sc_hd__a21o_2 _07437_ (.A1(_00355_),
    .A2(_00356_),
    .B1(net258),
    .X(_00357_));
 sky130_fd_sc_hd__and2_1 _07438_ (.A(_00354_),
    .B(_00357_),
    .X(_00358_));
 sky130_fd_sc_hd__nand2_8 _07439_ (.A(_00354_),
    .B(_00357_),
    .Y(_00359_));
 sky130_fd_sc_hd__o21ai_1 _07440_ (.A1(_00248_),
    .A2(_00249_),
    .B1(reg1_val[18]),
    .Y(_00360_));
 sky130_fd_sc_hd__a21o_1 _07441_ (.A1(_00350_),
    .A2(_00360_),
    .B1(net258),
    .X(_00361_));
 sky130_fd_sc_hd__nand2_1 _07442_ (.A(_04511_),
    .B(net258),
    .Y(_00362_));
 sky130_fd_sc_hd__and2_1 _07443_ (.A(_00361_),
    .B(_00362_),
    .X(_00363_));
 sky130_fd_sc_hd__a22o_1 _07444_ (.A1(_00354_),
    .A2(_00357_),
    .B1(_00361_),
    .B2(_00362_),
    .X(_00364_));
 sky130_fd_sc_hd__nand4_2 _07445_ (.A(_00354_),
    .B(_00357_),
    .C(_00361_),
    .D(_00362_),
    .Y(_00365_));
 sky130_fd_sc_hd__nor2_1 _07446_ (.A(net89),
    .B(_00365_),
    .Y(_00366_));
 sky130_fd_sc_hd__mux2_4 _07447_ (.A0(_00365_),
    .A1(_00364_),
    .S(net89),
    .X(_00367_));
 sky130_fd_sc_hd__a21oi_1 _07448_ (.A1(_06706_),
    .A2(_06707_),
    .B1(net178),
    .Y(_00368_));
 sky130_fd_sc_hd__nor2_1 _07449_ (.A(_06517_),
    .B(net178),
    .Y(_00369_));
 sky130_fd_sc_hd__a31o_4 _07450_ (.A1(_06517_),
    .A2(_06706_),
    .A3(_06707_),
    .B1(net178),
    .X(_00370_));
 sky130_fd_sc_hd__xor2_4 _07451_ (.A(_06509_),
    .B(_00370_),
    .X(_00371_));
 sky130_fd_sc_hd__xnor2_4 _07452_ (.A(_06509_),
    .B(_00370_),
    .Y(_00372_));
 sky130_fd_sc_hd__nand2_2 _07453_ (.A(_00364_),
    .B(_00365_),
    .Y(_00373_));
 sky130_fd_sc_hd__a31o_4 _07454_ (.A1(_06706_),
    .A2(_06707_),
    .A3(_06710_),
    .B1(net178),
    .X(_00374_));
 sky130_fd_sc_hd__xnor2_4 _07455_ (.A(_06495_),
    .B(_00374_),
    .Y(_00375_));
 sky130_fd_sc_hd__xnor2_4 _07456_ (.A(_06502_),
    .B(_00374_),
    .Y(_00376_));
 sky130_fd_sc_hd__o22a_1 _07457_ (.A1(net28),
    .A2(net123),
    .B1(net26),
    .B2(net120),
    .X(_00377_));
 sky130_fd_sc_hd__xnor2_1 _07458_ (.A(net88),
    .B(_00377_),
    .Y(_00378_));
 sky130_fd_sc_hd__xor2_1 _07459_ (.A(reg1_val[15]),
    .B(_00245_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _07460_ (.A0(reg1_val[15]),
    .A1(_00379_),
    .S(net260),
    .X(_00380_));
 sky130_fd_sc_hd__inv_6 _07461_ (.A(net117),
    .Y(_00381_));
 sky130_fd_sc_hd__xnor2_1 _07462_ (.A(reg1_val[16]),
    .B(_00247_),
    .Y(_00382_));
 sky130_fd_sc_hd__mux2_2 _07463_ (.A0(reg1_val[16]),
    .A1(_00382_),
    .S(net261),
    .X(_00383_));
 sky130_fd_sc_hd__and2_1 _07464_ (.A(net117),
    .B(_00383_),
    .X(_00384_));
 sky130_fd_sc_hd__nand2_1 _07465_ (.A(net118),
    .B(_00383_),
    .Y(_00385_));
 sky130_fd_sc_hd__nor2_1 _07466_ (.A(net118),
    .B(_00383_),
    .Y(_00386_));
 sky130_fd_sc_hd__or2_1 _07467_ (.A(net118),
    .B(_00383_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _07468_ (.A0(_00385_),
    .A1(_00387_),
    .S(net87),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _07469_ (.A0(_00384_),
    .A1(_00386_),
    .S(net87),
    .X(_00389_));
 sky130_fd_sc_hd__a41o_4 _07470_ (.A1(_06502_),
    .A2(_06706_),
    .A3(_06707_),
    .A4(_06710_),
    .B1(net178),
    .X(_00390_));
 sky130_fd_sc_hd__xnor2_4 _07471_ (.A(_06435_),
    .B(_00390_),
    .Y(_00391_));
 sky130_fd_sc_hd__xnor2_4 _07472_ (.A(_06426_),
    .B(_00390_),
    .Y(_00392_));
 sky130_fd_sc_hd__nor2_1 _07473_ (.A(_00384_),
    .B(_00386_),
    .Y(_00393_));
 sky130_fd_sc_hd__nand2_1 _07474_ (.A(_00385_),
    .B(_00387_),
    .Y(_00394_));
 sky130_fd_sc_hd__o21ai_4 _07475_ (.A1(net178),
    .A2(_06712_),
    .B1(_06363_),
    .Y(_00395_));
 sky130_fd_sc_hd__or3_4 _07476_ (.A(_06363_),
    .B(net178),
    .C(_06712_),
    .X(_00396_));
 sky130_fd_sc_hd__and2_4 _07477_ (.A(_00395_),
    .B(_00396_),
    .X(_00397_));
 sky130_fd_sc_hd__nand2_4 _07478_ (.A(_00395_),
    .B(_00396_),
    .Y(_00398_));
 sky130_fd_sc_hd__o22a_1 _07479_ (.A1(net24),
    .A2(net115),
    .B1(net22),
    .B2(net85),
    .X(_00399_));
 sky130_fd_sc_hd__xnor2_1 _07480_ (.A(net86),
    .B(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__a21o_1 _07481_ (.A1(net173),
    .A2(_00250_),
    .B1(_04521_),
    .X(_00401_));
 sky130_fd_sc_hd__a21o_1 _07482_ (.A1(_00269_),
    .A2(_00401_),
    .B1(net258),
    .X(_00402_));
 sky130_fd_sc_hd__nand2_1 _07483_ (.A(_04521_),
    .B(net258),
    .Y(_00403_));
 sky130_fd_sc_hd__and2_1 _07484_ (.A(_00402_),
    .B(_00403_),
    .X(_00404_));
 sky130_fd_sc_hd__a22o_1 _07485_ (.A1(_00349_),
    .A2(_00352_),
    .B1(_00402_),
    .B2(_00403_),
    .X(_00405_));
 sky130_fd_sc_hd__nand4_2 _07486_ (.A(_00349_),
    .B(_00352_),
    .C(_00402_),
    .D(_00403_),
    .Y(_00406_));
 sky130_fd_sc_hd__nor2_1 _07487_ (.A(net97),
    .B(_00406_),
    .Y(_00407_));
 sky130_fd_sc_hd__mux2_1 _07488_ (.A0(_00405_),
    .A1(_00406_),
    .S(_00274_),
    .X(_00408_));
 sky130_fd_sc_hd__a31o_4 _07489_ (.A1(_06538_),
    .A2(_06547_),
    .A3(_06706_),
    .B1(net178),
    .X(_00409_));
 sky130_fd_sc_hd__a41o_4 _07490_ (.A1(_06530_),
    .A2(_06538_),
    .A3(_06547_),
    .A4(_06706_),
    .B1(net178),
    .X(_00410_));
 sky130_fd_sc_hd__xor2_4 _07491_ (.A(_06523_),
    .B(_00410_),
    .X(_00411_));
 sky130_fd_sc_hd__xnor2_4 _07492_ (.A(_06523_),
    .B(_00410_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_2 _07493_ (.A(_00405_),
    .B(_00406_),
    .Y(_00413_));
 sky130_fd_sc_hd__o2bb2a_4 _07494_ (.A1_N(_06709_),
    .A2_N(_00369_),
    .B1(_00368_),
    .B2(_06516_),
    .X(_00414_));
 sky130_fd_sc_hd__a2bb2o_2 _07495_ (.A1_N(_06516_),
    .A2_N(_00368_),
    .B1(_00369_),
    .B2(_06709_),
    .X(_00415_));
 sky130_fd_sc_hd__o22a_1 _07496_ (.A1(net21),
    .A2(_00411_),
    .B1(net19),
    .B2(net110),
    .X(_00416_));
 sky130_fd_sc_hd__xnor2_1 _07497_ (.A(net96),
    .B(_00416_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _07498_ (.A(_00400_),
    .B(_00417_),
    .Y(_00418_));
 sky130_fd_sc_hd__or2_1 _07499_ (.A(_00400_),
    .B(_00417_),
    .X(_00419_));
 sky130_fd_sc_hd__nand2_1 _07500_ (.A(_00418_),
    .B(_00419_),
    .Y(_00420_));
 sky130_fd_sc_hd__inv_2 _07501_ (.A(_00420_),
    .Y(_00421_));
 sky130_fd_sc_hd__xor2_1 _07502_ (.A(_00378_),
    .B(_00420_),
    .X(_00422_));
 sky130_fd_sc_hd__a21oi_1 _07503_ (.A1(_00324_),
    .A2(_00347_),
    .B1(_00422_),
    .Y(_00423_));
 sky130_fd_sc_hd__and3_1 _07504_ (.A(_00324_),
    .B(_00347_),
    .C(_00422_),
    .X(_00424_));
 sky130_fd_sc_hd__nor2_2 _07505_ (.A(_00423_),
    .B(_00424_),
    .Y(_00425_));
 sky130_fd_sc_hd__xor2_4 _07506_ (.A(_00237_),
    .B(_00425_),
    .X(_00426_));
 sky130_fd_sc_hd__nor2_1 _07507_ (.A(reg1_val[13]),
    .B(net260),
    .Y(_00427_));
 sky130_fd_sc_hd__o31a_1 _07508_ (.A1(net290),
    .A2(reg1_val[12]),
    .A3(_00240_),
    .B1(reg1_val[13]),
    .X(_00428_));
 sky130_fd_sc_hd__o21a_2 _07509_ (.A1(_00244_),
    .A2(_00428_),
    .B1(net260),
    .X(_00429_));
 sky130_fd_sc_hd__nor2_1 _07510_ (.A(_00427_),
    .B(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__inv_8 _07511_ (.A(net108),
    .Y(_00431_));
 sky130_fd_sc_hd__a31o_1 _07512_ (.A1(_04478_),
    .A2(_00239_),
    .A3(_00242_),
    .B1(_04500_),
    .X(_00432_));
 sky130_fd_sc_hd__and2_1 _07513_ (.A(_00245_),
    .B(_00432_),
    .X(_00433_));
 sky130_fd_sc_hd__a21oi_2 _07514_ (.A1(_00245_),
    .A2(_00432_),
    .B1(net259),
    .Y(_00434_));
 sky130_fd_sc_hd__nor2_1 _07515_ (.A(reg1_val[14]),
    .B(net261),
    .Y(_00435_));
 sky130_fd_sc_hd__nor2_1 _07516_ (.A(_00434_),
    .B(_00435_),
    .Y(_00436_));
 sky130_fd_sc_hd__or4_1 _07517_ (.A(_00427_),
    .B(_00429_),
    .C(_00434_),
    .D(_00435_),
    .X(_00437_));
 sky130_fd_sc_hd__nor2_1 _07518_ (.A(net117),
    .B(_00437_),
    .Y(_00438_));
 sky130_fd_sc_hd__o22ai_2 _07519_ (.A1(_00427_),
    .A2(_00429_),
    .B1(_00434_),
    .B2(_00435_),
    .Y(_00439_));
 sky130_fd_sc_hd__mux2_1 _07520_ (.A0(_00437_),
    .A1(_00439_),
    .S(net117),
    .X(_00440_));
 sky130_fd_sc_hd__nor2_4 _07521_ (.A(net177),
    .B(_06713_),
    .Y(_00441_));
 sky130_fd_sc_hd__xnor2_4 _07522_ (.A(_06309_),
    .B(_00441_),
    .Y(_00442_));
 sky130_fd_sc_hd__xnor2_4 _07523_ (.A(_06315_),
    .B(_00441_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_2 _07524_ (.A(_00437_),
    .B(_00439_),
    .Y(_00444_));
 sky130_fd_sc_hd__a21oi_4 _07525_ (.A1(_06315_),
    .A2(_06713_),
    .B1(net178),
    .Y(_00445_));
 sky130_fd_sc_hd__xnor2_4 _07526_ (.A(_06251_),
    .B(_00445_),
    .Y(_00446_));
 sky130_fd_sc_hd__xnor2_2 _07527_ (.A(_06240_),
    .B(_00445_),
    .Y(_00447_));
 sky130_fd_sc_hd__o22a_1 _07528_ (.A1(net83),
    .A2(_00442_),
    .B1(net79),
    .B2(net77),
    .X(_00448_));
 sky130_fd_sc_hd__xnor2_1 _07529_ (.A(net116),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__nor2_1 _07530_ (.A(net290),
    .B(net260),
    .Y(_00450_));
 sky130_fd_sc_hd__xnor2_2 _07531_ (.A(_04478_),
    .B(_00239_),
    .Y(_00451_));
 sky130_fd_sc_hd__a21oi_2 _07532_ (.A1(net260),
    .A2(_00451_),
    .B1(_00450_),
    .Y(_00452_));
 sky130_fd_sc_hd__a21o_1 _07533_ (.A1(_04478_),
    .A2(_00239_),
    .B1(_04489_),
    .X(_00453_));
 sky130_fd_sc_hd__a21o_2 _07534_ (.A1(_00241_),
    .A2(_00453_),
    .B1(net259),
    .X(_00454_));
 sky130_fd_sc_hd__nand2_2 _07535_ (.A(_04489_),
    .B(net259),
    .Y(_00455_));
 sky130_fd_sc_hd__and2_1 _07536_ (.A(_00454_),
    .B(_00455_),
    .X(_00456_));
 sky130_fd_sc_hd__and3_1 _07537_ (.A(net145),
    .B(_00454_),
    .C(_00455_),
    .X(_00457_));
 sky130_fd_sc_hd__o2111a_2 _07538_ (.A1(_00427_),
    .A2(_00429_),
    .B1(net145),
    .C1(_00454_),
    .D1(_00455_),
    .X(_00458_));
 sky130_fd_sc_hd__a21oi_4 _07539_ (.A1(_00454_),
    .A2(_00455_),
    .B1(net145),
    .Y(_00459_));
 sky130_fd_sc_hd__a21oi_4 _07540_ (.A1(net108),
    .A2(_00459_),
    .B1(_00458_),
    .Y(_00460_));
 sky130_fd_sc_hd__a21o_4 _07541_ (.A1(net108),
    .A2(_00459_),
    .B1(_00458_),
    .X(_00461_));
 sky130_fd_sc_hd__a31o_4 _07542_ (.A1(_06251_),
    .A2(_06315_),
    .A3(_06713_),
    .B1(net177),
    .X(_00462_));
 sky130_fd_sc_hd__xor2_4 _07543_ (.A(_06165_),
    .B(_00462_),
    .X(_00463_));
 sky130_fd_sc_hd__xnor2_4 _07544_ (.A(_06165_),
    .B(_00462_),
    .Y(_00464_));
 sky130_fd_sc_hd__nor2_4 _07545_ (.A(_00457_),
    .B(_00459_),
    .Y(_00465_));
 sky130_fd_sc_hd__or2_4 _07546_ (.A(_00457_),
    .B(_00459_),
    .X(_00466_));
 sky130_fd_sc_hd__o2bb2a_4 _07547_ (.A1_N(_06716_),
    .A2_N(_00217_),
    .B1(_00216_),
    .B2(_06121_),
    .X(_00467_));
 sky130_fd_sc_hd__a2bb2o_2 _07548_ (.A1_N(_06121_),
    .A2_N(_00216_),
    .B1(_00217_),
    .B2(_06716_),
    .X(_00468_));
 sky130_fd_sc_hd__a22o_1 _07549_ (.A1(_00461_),
    .A2(_00464_),
    .B1(_00465_),
    .B2(net71),
    .X(_00469_));
 sky130_fd_sc_hd__xnor2_1 _07550_ (.A(_00431_),
    .B(_00469_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_2 _07551_ (.A(_00449_),
    .B(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__or2_1 _07552_ (.A(_00449_),
    .B(_00470_),
    .X(_00472_));
 sky130_fd_sc_hd__nand2_1 _07553_ (.A(_00471_),
    .B(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__o22a_1 _07554_ (.A1(net120),
    .A2(net24),
    .B1(_00391_),
    .B2(net22),
    .X(_00474_));
 sky130_fd_sc_hd__xnor2_1 _07555_ (.A(net87),
    .B(_00474_),
    .Y(_00475_));
 sky130_fd_sc_hd__xnor2_4 _07556_ (.A(_06529_),
    .B(_00409_),
    .Y(_00476_));
 sky130_fd_sc_hd__xnor2_4 _07557_ (.A(_06530_),
    .B(_00409_),
    .Y(_00477_));
 sky130_fd_sc_hd__o22a_1 _07558_ (.A1(_00411_),
    .A2(net19),
    .B1(net106),
    .B2(net21),
    .X(_00478_));
 sky130_fd_sc_hd__xnor2_1 _07559_ (.A(net97),
    .B(_00478_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _07560_ (.A(_00475_),
    .B(_00479_),
    .Y(_00480_));
 sky130_fd_sc_hd__o22a_1 _07561_ (.A1(net123),
    .A2(net26),
    .B1(net110),
    .B2(net28),
    .X(_00481_));
 sky130_fd_sc_hd__xor2_1 _07562_ (.A(net88),
    .B(_00481_),
    .X(_00482_));
 sky130_fd_sc_hd__xnor2_1 _07563_ (.A(_00475_),
    .B(_00479_),
    .Y(_00483_));
 sky130_fd_sc_hd__or2_1 _07564_ (.A(_00482_),
    .B(_00483_),
    .X(_00484_));
 sky130_fd_sc_hd__a21oi_1 _07565_ (.A1(_00480_),
    .A2(_00484_),
    .B1(_00473_),
    .Y(_00485_));
 sky130_fd_sc_hd__and3_1 _07566_ (.A(_00473_),
    .B(_00480_),
    .C(_00484_),
    .X(_00486_));
 sky130_fd_sc_hd__or2_1 _07567_ (.A(_00485_),
    .B(_00486_),
    .X(_00487_));
 sky130_fd_sc_hd__o22a_1 _07568_ (.A1(net85),
    .A2(net83),
    .B1(net82),
    .B2(net79),
    .X(_00488_));
 sky130_fd_sc_hd__xnor2_1 _07569_ (.A(net118),
    .B(_00488_),
    .Y(_00489_));
 sky130_fd_sc_hd__o31a_1 _07570_ (.A1(net287),
    .A2(_00185_),
    .A3(_00213_),
    .B1(reg1_val[10]),
    .X(_00490_));
 sky130_fd_sc_hd__nor2_1 _07571_ (.A(_00239_),
    .B(_00490_),
    .Y(_00491_));
 sky130_fd_sc_hd__mux2_1 _07572_ (.A0(reg1_val[10]),
    .A1(_00491_),
    .S(net260),
    .X(_00492_));
 sky130_fd_sc_hd__nor2_1 _07573_ (.A(net155),
    .B(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__and2_1 _07574_ (.A(net155),
    .B(_00492_),
    .X(_00494_));
 sky130_fd_sc_hd__and3b_1 _07575_ (.A_N(net145),
    .B(_00492_),
    .C(net154),
    .X(_00495_));
 sky130_fd_sc_hd__a21oi_1 _07576_ (.A1(net145),
    .A2(_00493_),
    .B1(_00495_),
    .Y(_00496_));
 sky130_fd_sc_hd__or2_2 _07577_ (.A(_00493_),
    .B(_00494_),
    .X(_00497_));
 sky130_fd_sc_hd__o22a_1 _07578_ (.A1(net70),
    .A2(net68),
    .B1(net66),
    .B2(net103),
    .X(_00498_));
 sky130_fd_sc_hd__xnor2_1 _07579_ (.A(net146),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__and2_1 _07580_ (.A(_00489_),
    .B(_00499_),
    .X(_00500_));
 sky130_fd_sc_hd__a22o_1 _07581_ (.A1(net78),
    .A2(_00461_),
    .B1(_00464_),
    .B2(_00465_),
    .X(_00501_));
 sky130_fd_sc_hd__xnor2_1 _07582_ (.A(_00431_),
    .B(_00501_),
    .Y(_00502_));
 sky130_fd_sc_hd__nor2_1 _07583_ (.A(_00489_),
    .B(_00499_),
    .Y(_00503_));
 sky130_fd_sc_hd__or2_1 _07584_ (.A(_00500_),
    .B(_00503_),
    .X(_00504_));
 sky130_fd_sc_hd__inv_2 _07585_ (.A(_00504_),
    .Y(_00505_));
 sky130_fd_sc_hd__a21o_1 _07586_ (.A1(_00502_),
    .A2(_00505_),
    .B1(_00500_),
    .X(_00506_));
 sky130_fd_sc_hd__and2b_1 _07587_ (.A_N(_00487_),
    .B(_00506_),
    .X(_00507_));
 sky130_fd_sc_hd__xor2_1 _07588_ (.A(_00487_),
    .B(_00506_),
    .X(_00508_));
 sky130_fd_sc_hd__o22a_1 _07589_ (.A1(net49),
    .A2(net132),
    .B1(net157),
    .B2(net51),
    .X(_00509_));
 sky130_fd_sc_hd__xnor2_2 _07590_ (.A(net202),
    .B(_00509_),
    .Y(_00510_));
 sky130_fd_sc_hd__o22a_1 _07591_ (.A1(net133),
    .A2(net47),
    .B1(net45),
    .B2(net158),
    .X(_00511_));
 sky130_fd_sc_hd__xnor2_2 _07592_ (.A(net179),
    .B(_00511_),
    .Y(_00512_));
 sky130_fd_sc_hd__a21oi_4 _07593_ (.A1(_06703_),
    .A2(_00174_),
    .B1(_05221_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_2 _07594_ (.A(_05221_),
    .B(_06703_),
    .Y(_00514_));
 sky130_fd_sc_hd__nor2_8 _07595_ (.A(_00173_),
    .B(_00514_),
    .Y(_00515_));
 sky130_fd_sc_hd__nor2_8 _07596_ (.A(_00513_),
    .B(_00515_),
    .Y(_00516_));
 sky130_fd_sc_hd__or2_4 _07597_ (.A(_00513_),
    .B(_00515_),
    .X(_00517_));
 sky130_fd_sc_hd__o22a_1 _07598_ (.A1(net236),
    .A2(net44),
    .B1(_00517_),
    .B2(net286),
    .X(_00518_));
 sky130_fd_sc_hd__xnor2_2 _07599_ (.A(net199),
    .B(_00518_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _07600_ (.A(_00512_),
    .B(_00519_),
    .Y(_00520_));
 sky130_fd_sc_hd__xnor2_2 _07601_ (.A(_00512_),
    .B(_00519_),
    .Y(_00521_));
 sky130_fd_sc_hd__or2_1 _07602_ (.A(_00510_),
    .B(_00521_),
    .X(_00522_));
 sky130_fd_sc_hd__xnor2_2 _07603_ (.A(_00510_),
    .B(_00521_),
    .Y(_00523_));
 sky130_fd_sc_hd__o22a_1 _07604_ (.A1(net56),
    .A2(net131),
    .B1(net40),
    .B2(net105),
    .X(_00524_));
 sky130_fd_sc_hd__xnor2_1 _07605_ (.A(net174),
    .B(_00524_),
    .Y(_00525_));
 sky130_fd_sc_hd__a22o_1 _07606_ (.A1(net129),
    .A2(_00229_),
    .B1(net126),
    .B2(_00203_),
    .X(_00526_));
 sky130_fd_sc_hd__xor2_1 _07607_ (.A(net154),
    .B(_00526_),
    .X(_00527_));
 sky130_fd_sc_hd__nand2_1 _07608_ (.A(_00525_),
    .B(_00527_),
    .Y(_00528_));
 sky130_fd_sc_hd__a22o_1 _07609_ (.A1(_00203_),
    .A2(net129),
    .B1(net127),
    .B2(_00208_),
    .X(_00529_));
 sky130_fd_sc_hd__xnor2_2 _07610_ (.A(net154),
    .B(_00529_),
    .Y(_00530_));
 sky130_fd_sc_hd__o22a_1 _07611_ (.A1(net103),
    .A2(net68),
    .B1(net66),
    .B2(net100),
    .X(_00531_));
 sky130_fd_sc_hd__xnor2_2 _07612_ (.A(net146),
    .B(_00531_),
    .Y(_00532_));
 sky130_fd_sc_hd__o22a_1 _07613_ (.A1(net56),
    .A2(net105),
    .B1(net131),
    .B2(net53),
    .X(_00533_));
 sky130_fd_sc_hd__xnor2_2 _07614_ (.A(net174),
    .B(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__nand2_1 _07615_ (.A(_00532_),
    .B(_00534_),
    .Y(_00535_));
 sky130_fd_sc_hd__xnor2_2 _07616_ (.A(_00532_),
    .B(_00534_),
    .Y(_00536_));
 sky130_fd_sc_hd__xnor2_2 _07617_ (.A(_00530_),
    .B(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__or2_1 _07618_ (.A(_00528_),
    .B(_00537_),
    .X(_00538_));
 sky130_fd_sc_hd__xnor2_2 _07619_ (.A(_00528_),
    .B(_00537_),
    .Y(_00539_));
 sky130_fd_sc_hd__xnor2_2 _07620_ (.A(_00523_),
    .B(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__a22o_1 _07621_ (.A1(net14),
    .A2(net148),
    .B1(net30),
    .B2(_00266_),
    .X(_00541_));
 sky130_fd_sc_hd__xnor2_1 _07622_ (.A(net92),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__o22a_1 _07623_ (.A1(net35),
    .A2(net152),
    .B1(net33),
    .B2(net151),
    .X(_00543_));
 sky130_fd_sc_hd__xnor2_1 _07624_ (.A(net95),
    .B(_00543_),
    .Y(_00544_));
 sky130_fd_sc_hd__o22a_1 _07625_ (.A1(net39),
    .A2(_00286_),
    .B1(net37),
    .B2(_00477_),
    .X(_00545_));
 sky130_fd_sc_hd__xnor2_1 _07626_ (.A(net99),
    .B(_00545_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _07627_ (.A(_00544_),
    .B(_00546_),
    .Y(_00547_));
 sky130_fd_sc_hd__xnor2_1 _07628_ (.A(_00544_),
    .B(_00546_),
    .Y(_00548_));
 sky130_fd_sc_hd__or2_1 _07629_ (.A(_00542_),
    .B(_00548_),
    .X(_00549_));
 sky130_fd_sc_hd__nand2_1 _07630_ (.A(_00542_),
    .B(_00548_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _07631_ (.A(_00549_),
    .B(_00550_),
    .Y(_00551_));
 sky130_fd_sc_hd__nor2_1 _07632_ (.A(_00540_),
    .B(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__xor2_2 _07633_ (.A(_00540_),
    .B(_00551_),
    .X(_00553_));
 sky130_fd_sc_hd__or4_4 _07634_ (.A(reg1_val[28]),
    .B(_00248_),
    .C(_00255_),
    .D(_00294_),
    .X(_00554_));
 sky130_fd_sc_hd__a31o_1 _07635_ (.A1(_00247_),
    .A2(_00254_),
    .A3(_00295_),
    .B1(_04587_),
    .X(_00555_));
 sky130_fd_sc_hd__a21o_1 _07636_ (.A1(_00554_),
    .A2(_00555_),
    .B1(net258),
    .X(_00556_));
 sky130_fd_sc_hd__nand2_1 _07637_ (.A(_04587_),
    .B(net258),
    .Y(_00557_));
 sky130_fd_sc_hd__and2_1 _07638_ (.A(_00556_),
    .B(_00557_),
    .X(_00558_));
 sky130_fd_sc_hd__nor2_1 _07639_ (.A(net93),
    .B(_00558_),
    .Y(_00559_));
 sky130_fd_sc_hd__a22o_1 _07640_ (.A1(_00291_),
    .A2(_00300_),
    .B1(_00556_),
    .B2(_00557_),
    .X(_00560_));
 sky130_fd_sc_hd__nand4_2 _07641_ (.A(_00291_),
    .B(_00300_),
    .C(_00556_),
    .D(_00557_),
    .Y(_00561_));
 sky130_fd_sc_hd__and2_1 _07642_ (.A(_00560_),
    .B(_00561_),
    .X(_00562_));
 sky130_fd_sc_hd__nand2_1 _07643_ (.A(net207),
    .B(net17),
    .Y(_00563_));
 sky130_fd_sc_hd__nand3b_1 _07644_ (.A_N(_00563_),
    .B(_00182_),
    .C(_00180_),
    .Y(_00564_));
 sky130_fd_sc_hd__a21bo_1 _07645_ (.A1(_00180_),
    .A2(_00182_),
    .B1_N(_00563_),
    .X(_00565_));
 sky130_fd_sc_hd__nand2_1 _07646_ (.A(_00564_),
    .B(_00565_),
    .Y(_00566_));
 sky130_fd_sc_hd__xnor2_1 _07647_ (.A(_00553_),
    .B(_00566_),
    .Y(_00567_));
 sky130_fd_sc_hd__nor2_1 _07648_ (.A(_00508_),
    .B(_00567_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _07649_ (.A(_00508_),
    .B(_00567_),
    .Y(_00569_));
 sky130_fd_sc_hd__and2b_1 _07650_ (.A_N(_00568_),
    .B(_00569_),
    .X(_00570_));
 sky130_fd_sc_hd__xor2_4 _07651_ (.A(_00426_),
    .B(_00570_),
    .X(_00571_));
 sky130_fd_sc_hd__nand2_1 _07652_ (.A(_00344_),
    .B(_00346_),
    .Y(_00572_));
 sky130_fd_sc_hd__nand2_1 _07653_ (.A(_00347_),
    .B(_00572_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _07654_ (.A(_00482_),
    .B(_00483_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _07655_ (.A(_00484_),
    .B(_00574_),
    .Y(_00575_));
 sky130_fd_sc_hd__xnor2_1 _07656_ (.A(_00235_),
    .B(_00236_),
    .Y(_00576_));
 sky130_fd_sc_hd__nor2_1 _07657_ (.A(_00575_),
    .B(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__xor2_1 _07658_ (.A(_00575_),
    .B(_00576_),
    .X(_00578_));
 sky130_fd_sc_hd__xnor2_1 _07659_ (.A(_00573_),
    .B(_00578_),
    .Y(_00579_));
 sky130_fd_sc_hd__o22a_1 _07660_ (.A1(net74),
    .A2(net68),
    .B1(net66),
    .B2(net70),
    .X(_00580_));
 sky130_fd_sc_hd__xnor2_1 _07661_ (.A(net146),
    .B(_00580_),
    .Y(_00581_));
 sky130_fd_sc_hd__o22a_1 _07662_ (.A1(net115),
    .A2(net83),
    .B1(net79),
    .B2(net85),
    .X(_00582_));
 sky130_fd_sc_hd__xnor2_1 _07663_ (.A(net116),
    .B(_00582_),
    .Y(_00583_));
 sky130_fd_sc_hd__and2_1 _07664_ (.A(_00581_),
    .B(_00583_),
    .X(_00584_));
 sky130_fd_sc_hd__o22a_1 _07665_ (.A1(net82),
    .A2(net75),
    .B1(net72),
    .B2(net76),
    .X(_00585_));
 sky130_fd_sc_hd__xnor2_1 _07666_ (.A(net108),
    .B(_00585_),
    .Y(_00586_));
 sky130_fd_sc_hd__nor2_1 _07667_ (.A(_00581_),
    .B(_00583_),
    .Y(_00587_));
 sky130_fd_sc_hd__or2_1 _07668_ (.A(_00584_),
    .B(_00587_),
    .X(_00588_));
 sky130_fd_sc_hd__inv_2 _07669_ (.A(_00588_),
    .Y(_00589_));
 sky130_fd_sc_hd__a21o_1 _07670_ (.A1(_00586_),
    .A2(_00589_),
    .B1(_00584_),
    .X(_00590_));
 sky130_fd_sc_hd__or2_1 _07671_ (.A(_00525_),
    .B(_00527_),
    .X(_00591_));
 sky130_fd_sc_hd__nand2_1 _07672_ (.A(_00528_),
    .B(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__o22a_1 _07673_ (.A1(_00371_),
    .A2(net24),
    .B1(net22),
    .B2(net119),
    .X(_00593_));
 sky130_fd_sc_hd__xnor2_1 _07674_ (.A(net86),
    .B(_00593_),
    .Y(_00594_));
 sky130_fd_sc_hd__o22a_1 _07675_ (.A1(_00286_),
    .A2(net21),
    .B1(net19),
    .B2(_00477_),
    .X(_00595_));
 sky130_fd_sc_hd__xnor2_1 _07676_ (.A(net96),
    .B(_00595_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_1 _07677_ (.A(_00594_),
    .B(_00596_),
    .Y(_00597_));
 sky130_fd_sc_hd__o22a_1 _07678_ (.A1(net28),
    .A2(_00411_),
    .B1(net110),
    .B2(net26),
    .X(_00598_));
 sky130_fd_sc_hd__xor2_1 _07679_ (.A(net88),
    .B(_00598_),
    .X(_00599_));
 sky130_fd_sc_hd__xnor2_1 _07680_ (.A(_00594_),
    .B(_00596_),
    .Y(_00600_));
 sky130_fd_sc_hd__or2_1 _07681_ (.A(_00599_),
    .B(_00600_),
    .X(_00601_));
 sky130_fd_sc_hd__a21oi_1 _07682_ (.A1(_00597_),
    .A2(_00601_),
    .B1(_00592_),
    .Y(_00602_));
 sky130_fd_sc_hd__and3_1 _07683_ (.A(_00592_),
    .B(_00597_),
    .C(_00601_),
    .X(_00603_));
 sky130_fd_sc_hd__or2_1 _07684_ (.A(_00602_),
    .B(_00603_),
    .X(_00604_));
 sky130_fd_sc_hd__and2b_1 _07685_ (.A_N(_00604_),
    .B(_00590_),
    .X(_00605_));
 sky130_fd_sc_hd__xnor2_1 _07686_ (.A(_00590_),
    .B(_00604_),
    .Y(_00606_));
 sky130_fd_sc_hd__xor2_2 _07687_ (.A(_00164_),
    .B(_00165_),
    .X(_00607_));
 sky130_fd_sc_hd__nand2_1 _07688_ (.A(net95),
    .B(_00607_),
    .Y(_00608_));
 sky130_fd_sc_hd__o22a_1 _07689_ (.A1(net53),
    .A2(net132),
    .B1(net157),
    .B2(net47),
    .X(_00609_));
 sky130_fd_sc_hd__xnor2_1 _07690_ (.A(net201),
    .B(_00609_),
    .Y(_00610_));
 sky130_fd_sc_hd__o22a_1 _07691_ (.A1(net286),
    .A2(net49),
    .B1(net45),
    .B2(net236),
    .X(_00611_));
 sky130_fd_sc_hd__xnor2_1 _07692_ (.A(net199),
    .B(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2b_1 _07693_ (.A_N(_00610_),
    .B(_00612_),
    .Y(_00613_));
 sky130_fd_sc_hd__xnor2_2 _07694_ (.A(net95),
    .B(_00607_),
    .Y(_00614_));
 sky130_fd_sc_hd__o21a_1 _07695_ (.A1(_00613_),
    .A2(_00614_),
    .B1(_00608_),
    .X(_00615_));
 sky130_fd_sc_hd__xor2_1 _07696_ (.A(_00502_),
    .B(_00504_),
    .X(_00616_));
 sky130_fd_sc_hd__o22a_1 _07697_ (.A1(_00267_),
    .A2(net37),
    .B1(_00339_),
    .B2(net39),
    .X(_00617_));
 sky130_fd_sc_hd__xnor2_1 _07698_ (.A(net99),
    .B(_00617_),
    .Y(_00618_));
 sky130_fd_sc_hd__nor2_1 _07699_ (.A(net212),
    .B(net33),
    .Y(_00619_));
 sky130_fd_sc_hd__xnor2_1 _07700_ (.A(net95),
    .B(_00619_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2b_1 _07701_ (.A_N(_00620_),
    .B(_00618_),
    .Y(_00621_));
 sky130_fd_sc_hd__a22o_1 _07702_ (.A1(net153),
    .A2(net14),
    .B1(net30),
    .B2(_00327_),
    .X(_00622_));
 sky130_fd_sc_hd__xnor2_1 _07703_ (.A(net91),
    .B(_00622_),
    .Y(_00623_));
 sky130_fd_sc_hd__xnor2_1 _07704_ (.A(_00618_),
    .B(_00620_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _07705_ (.A(_00623_),
    .B(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__a21o_1 _07706_ (.A1(_00621_),
    .A2(_00625_),
    .B1(_00616_),
    .X(_00626_));
 sky130_fd_sc_hd__nand3_1 _07707_ (.A(_00616_),
    .B(_00621_),
    .C(_00625_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _07708_ (.A(_00626_),
    .B(_00627_),
    .Y(_00628_));
 sky130_fd_sc_hd__xnor2_1 _07709_ (.A(_00615_),
    .B(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__xnor2_1 _07710_ (.A(_00579_),
    .B(_00606_),
    .Y(_00630_));
 sky130_fd_sc_hd__or2_1 _07711_ (.A(_00629_),
    .B(_00630_),
    .X(_00631_));
 sky130_fd_sc_hd__a21bo_1 _07712_ (.A1(_00579_),
    .A2(_00606_),
    .B1_N(_00631_),
    .X(_00632_));
 sky130_fd_sc_hd__xnor2_2 _07713_ (.A(_00613_),
    .B(_00614_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_1 _07714_ (.A(_00599_),
    .B(_00600_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _07715_ (.A(_00601_),
    .B(_00634_),
    .Y(_00635_));
 sky130_fd_sc_hd__or2_1 _07716_ (.A(_00633_),
    .B(_00635_),
    .X(_00636_));
 sky130_fd_sc_hd__or2_1 _07717_ (.A(_00623_),
    .B(_00624_),
    .X(_00637_));
 sky130_fd_sc_hd__nand2_1 _07718_ (.A(_00625_),
    .B(_00637_),
    .Y(_00638_));
 sky130_fd_sc_hd__xnor2_2 _07719_ (.A(_00633_),
    .B(_00635_),
    .Y(_00639_));
 sky130_fd_sc_hd__o21ai_2 _07720_ (.A1(_00638_),
    .A2(_00639_),
    .B1(_00636_),
    .Y(_00640_));
 sky130_fd_sc_hd__nand2_1 _07721_ (.A(_00211_),
    .B(_00234_),
    .Y(_00641_));
 sky130_fd_sc_hd__nand2b_1 _07722_ (.A_N(_00235_),
    .B(_00641_),
    .Y(_00642_));
 sky130_fd_sc_hd__o22a_1 _07723_ (.A1(net76),
    .A2(net68),
    .B1(net66),
    .B2(net74),
    .X(_00643_));
 sky130_fd_sc_hd__xnor2_1 _07724_ (.A(net146),
    .B(_00643_),
    .Y(_00644_));
 sky130_fd_sc_hd__o22a_1 _07725_ (.A1(net119),
    .A2(net83),
    .B1(net79),
    .B2(_00391_),
    .X(_00645_));
 sky130_fd_sc_hd__xnor2_1 _07726_ (.A(net116),
    .B(_00645_),
    .Y(_00646_));
 sky130_fd_sc_hd__nand2_1 _07727_ (.A(_00644_),
    .B(_00646_),
    .Y(_00647_));
 sky130_fd_sc_hd__o22a_1 _07728_ (.A1(net85),
    .A2(net75),
    .B1(net72),
    .B2(net82),
    .X(_00648_));
 sky130_fd_sc_hd__xnor2_1 _07729_ (.A(net108),
    .B(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__inv_2 _07730_ (.A(_00649_),
    .Y(_00650_));
 sky130_fd_sc_hd__or2_1 _07731_ (.A(_00644_),
    .B(_00646_),
    .X(_00651_));
 sky130_fd_sc_hd__nand2_1 _07732_ (.A(_00647_),
    .B(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hd__or2_1 _07733_ (.A(_00650_),
    .B(_00652_),
    .X(_00653_));
 sky130_fd_sc_hd__a21oi_1 _07734_ (.A1(_00647_),
    .A2(_00653_),
    .B1(_00642_),
    .Y(_00654_));
 sky130_fd_sc_hd__a22o_1 _07735_ (.A1(_00220_),
    .A2(net127),
    .B1(net71),
    .B2(net128),
    .X(_00655_));
 sky130_fd_sc_hd__xor2_1 _07736_ (.A(net154),
    .B(_00655_),
    .X(_00656_));
 sky130_fd_sc_hd__o22a_1 _07737_ (.A1(net56),
    .A2(net158),
    .B1(net40),
    .B2(net133),
    .X(_00657_));
 sky130_fd_sc_hd__xnor2_1 _07738_ (.A(net179),
    .B(_00657_),
    .Y(_00658_));
 sky130_fd_sc_hd__o22a_1 _07739_ (.A1(net42),
    .A2(net131),
    .B1(net100),
    .B2(net105),
    .X(_00659_));
 sky130_fd_sc_hd__xnor2_1 _07740_ (.A(_00188_),
    .B(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__xnor2_1 _07741_ (.A(_00656_),
    .B(_00658_),
    .Y(_00661_));
 sky130_fd_sc_hd__nor2_1 _07742_ (.A(_00660_),
    .B(_00661_),
    .Y(_00662_));
 sky130_fd_sc_hd__a21oi_1 _07743_ (.A1(_00656_),
    .A2(_00658_),
    .B1(_00662_),
    .Y(_00663_));
 sky130_fd_sc_hd__and3_1 _07744_ (.A(_00642_),
    .B(_00647_),
    .C(_00653_),
    .X(_00664_));
 sky130_fd_sc_hd__nor2_1 _07745_ (.A(_00654_),
    .B(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__and2b_1 _07746_ (.A_N(_00663_),
    .B(_00665_),
    .X(_00666_));
 sky130_fd_sc_hd__nor2_1 _07747_ (.A(_00654_),
    .B(_00666_),
    .Y(_00667_));
 sky130_fd_sc_hd__o21a_1 _07748_ (.A1(_00654_),
    .A2(_00666_),
    .B1(_00640_),
    .X(_00668_));
 sky130_fd_sc_hd__xor2_1 _07749_ (.A(_00586_),
    .B(_00588_),
    .X(_00669_));
 sky130_fd_sc_hd__o22a_1 _07750_ (.A1(net125),
    .A2(net21),
    .B1(net19),
    .B2(_00286_),
    .X(_00670_));
 sky130_fd_sc_hd__xnor2_1 _07751_ (.A(net96),
    .B(_00670_),
    .Y(_00671_));
 sky130_fd_sc_hd__o22a_1 _07752_ (.A1(net123),
    .A2(net22),
    .B1(net110),
    .B2(net24),
    .X(_00672_));
 sky130_fd_sc_hd__xnor2_1 _07753_ (.A(net86),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__nand2_1 _07754_ (.A(_00671_),
    .B(_00673_),
    .Y(_00674_));
 sky130_fd_sc_hd__o22a_1 _07755_ (.A1(net26),
    .A2(net113),
    .B1(_00477_),
    .B2(net28),
    .X(_00675_));
 sky130_fd_sc_hd__xor2_1 _07756_ (.A(net88),
    .B(_00675_),
    .X(_00676_));
 sky130_fd_sc_hd__xnor2_1 _07757_ (.A(_00671_),
    .B(_00673_),
    .Y(_00677_));
 sky130_fd_sc_hd__or2_1 _07758_ (.A(_00676_),
    .B(_00677_),
    .X(_00678_));
 sky130_fd_sc_hd__a21oi_1 _07759_ (.A1(_00674_),
    .A2(_00678_),
    .B1(_00669_),
    .Y(_00679_));
 sky130_fd_sc_hd__o22a_1 _07760_ (.A1(net56),
    .A2(net132),
    .B1(net157),
    .B2(net53),
    .X(_00680_));
 sky130_fd_sc_hd__xnor2_2 _07761_ (.A(net200),
    .B(_00680_),
    .Y(_00681_));
 sky130_fd_sc_hd__o22a_1 _07762_ (.A1(net236),
    .A2(net47),
    .B1(net45),
    .B2(net286),
    .X(_00682_));
 sky130_fd_sc_hd__xnor2_1 _07763_ (.A(_06736_),
    .B(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__o22a_1 _07764_ (.A1(net39),
    .A2(net151),
    .B1(_00339_),
    .B2(net37),
    .X(_00684_));
 sky130_fd_sc_hd__xnor2_1 _07765_ (.A(net99),
    .B(_00684_),
    .Y(_00685_));
 sky130_fd_sc_hd__and3_1 _07766_ (.A(_00681_),
    .B(_00683_),
    .C(_00685_),
    .X(_00686_));
 sky130_fd_sc_hd__a22o_1 _07767_ (.A1(net207),
    .A2(net14),
    .B1(net30),
    .B2(net153),
    .X(_00687_));
 sky130_fd_sc_hd__xnor2_1 _07768_ (.A(net92),
    .B(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__a21oi_1 _07769_ (.A1(_00681_),
    .A2(_00683_),
    .B1(_00685_),
    .Y(_00689_));
 sky130_fd_sc_hd__or3_1 _07770_ (.A(_00686_),
    .B(_00688_),
    .C(_00689_),
    .X(_00690_));
 sky130_fd_sc_hd__nand2b_1 _07771_ (.A_N(_00686_),
    .B(_00690_),
    .Y(_00691_));
 sky130_fd_sc_hd__and3_1 _07772_ (.A(_00669_),
    .B(_00674_),
    .C(_00678_),
    .X(_00692_));
 sky130_fd_sc_hd__nor2_1 _07773_ (.A(_00679_),
    .B(_00692_),
    .Y(_00693_));
 sky130_fd_sc_hd__or2_1 _07774_ (.A(_00679_),
    .B(_00692_),
    .X(_00694_));
 sky130_fd_sc_hd__a21o_1 _07775_ (.A1(_00691_),
    .A2(_00693_),
    .B1(_00679_),
    .X(_00695_));
 sky130_fd_sc_hd__xnor2_2 _07776_ (.A(_00640_),
    .B(_00667_),
    .Y(_00696_));
 sky130_fd_sc_hd__a21o_1 _07777_ (.A1(_00695_),
    .A2(_00696_),
    .B1(_00668_),
    .X(_00697_));
 sky130_fd_sc_hd__o21ai_2 _07778_ (.A1(_00615_),
    .A2(_00628_),
    .B1(_00626_),
    .Y(_00698_));
 sky130_fd_sc_hd__a31o_1 _07779_ (.A1(_00347_),
    .A2(_00572_),
    .A3(_00578_),
    .B1(_00577_),
    .X(_00699_));
 sky130_fd_sc_hd__nor2_1 _07780_ (.A(_00602_),
    .B(_00605_),
    .Y(_00700_));
 sky130_fd_sc_hd__o21a_1 _07781_ (.A1(_00602_),
    .A2(_00605_),
    .B1(_00699_),
    .X(_00701_));
 sky130_fd_sc_hd__xnor2_2 _07782_ (.A(_00699_),
    .B(_00700_),
    .Y(_00702_));
 sky130_fd_sc_hd__xor2_1 _07783_ (.A(_00698_),
    .B(_00702_),
    .X(_00703_));
 sky130_fd_sc_hd__xnor2_1 _07784_ (.A(_00697_),
    .B(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__nand2b_1 _07785_ (.A_N(_00704_),
    .B(_00632_),
    .Y(_00705_));
 sky130_fd_sc_hd__xnor2_2 _07786_ (.A(_00632_),
    .B(_00704_),
    .Y(_00706_));
 sky130_fd_sc_hd__and2_1 _07787_ (.A(_00571_),
    .B(_00706_),
    .X(_00707_));
 sky130_fd_sc_hd__xor2_1 _07788_ (.A(_00610_),
    .B(_00612_),
    .X(_00708_));
 sky130_fd_sc_hd__o22a_1 _07789_ (.A1(net123),
    .A2(net84),
    .B1(net80),
    .B2(net119),
    .X(_00709_));
 sky130_fd_sc_hd__xnor2_2 _07790_ (.A(net116),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__o22a_1 _07791_ (.A1(net82),
    .A2(net68),
    .B1(net66),
    .B2(net76),
    .X(_00711_));
 sky130_fd_sc_hd__xnor2_2 _07792_ (.A(net146),
    .B(_00711_),
    .Y(_00712_));
 sky130_fd_sc_hd__and2_1 _07793_ (.A(_00710_),
    .B(_00712_),
    .X(_00713_));
 sky130_fd_sc_hd__o22a_1 _07794_ (.A1(net115),
    .A2(net75),
    .B1(net72),
    .B2(net85),
    .X(_00714_));
 sky130_fd_sc_hd__xnor2_2 _07795_ (.A(net108),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__xor2_2 _07796_ (.A(_00710_),
    .B(_00712_),
    .X(_00716_));
 sky130_fd_sc_hd__a21oi_2 _07797_ (.A1(_00715_),
    .A2(_00716_),
    .B1(_00713_),
    .Y(_00717_));
 sky130_fd_sc_hd__xor2_1 _07798_ (.A(_00708_),
    .B(_00717_),
    .X(_00718_));
 sky130_fd_sc_hd__o22a_1 _07799_ (.A1(net133),
    .A2(net42),
    .B1(net40),
    .B2(net158),
    .X(_00719_));
 sky130_fd_sc_hd__xnor2_1 _07800_ (.A(net179),
    .B(_00719_),
    .Y(_00720_));
 sky130_fd_sc_hd__a22o_1 _07801_ (.A1(net128),
    .A2(_00464_),
    .B1(net71),
    .B2(net126),
    .X(_00721_));
 sky130_fd_sc_hd__xor2_1 _07802_ (.A(net154),
    .B(_00721_),
    .X(_00722_));
 sky130_fd_sc_hd__and2_1 _07803_ (.A(_00720_),
    .B(_00722_),
    .X(_00723_));
 sky130_fd_sc_hd__o22a_1 _07804_ (.A1(net105),
    .A2(net103),
    .B1(net100),
    .B2(net131),
    .X(_00724_));
 sky130_fd_sc_hd__xnor2_2 _07805_ (.A(net174),
    .B(_00724_),
    .Y(_00725_));
 sky130_fd_sc_hd__inv_2 _07806_ (.A(_00725_),
    .Y(_00726_));
 sky130_fd_sc_hd__xnor2_1 _07807_ (.A(_00720_),
    .B(_00722_),
    .Y(_00727_));
 sky130_fd_sc_hd__nor2_1 _07808_ (.A(_00726_),
    .B(_00727_),
    .Y(_00728_));
 sky130_fd_sc_hd__o21ai_1 _07809_ (.A1(_00723_),
    .A2(_00728_),
    .B1(_00718_),
    .Y(_00729_));
 sky130_fd_sc_hd__o21a_1 _07810_ (.A1(_00708_),
    .A2(_00717_),
    .B1(_00729_),
    .X(_00730_));
 sky130_fd_sc_hd__xnor2_1 _07811_ (.A(_00649_),
    .B(_00652_),
    .Y(_00731_));
 sky130_fd_sc_hd__o21ai_1 _07812_ (.A1(_00686_),
    .A2(_00689_),
    .B1(_00688_),
    .Y(_00732_));
 sky130_fd_sc_hd__and3_1 _07813_ (.A(_00690_),
    .B(_00731_),
    .C(_00732_),
    .X(_00733_));
 sky130_fd_sc_hd__nand2_1 _07814_ (.A(_00676_),
    .B(_00677_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand2_1 _07815_ (.A(_00678_),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__a21oi_1 _07816_ (.A1(_00690_),
    .A2(_00732_),
    .B1(_00731_),
    .Y(_00736_));
 sky130_fd_sc_hd__or3_1 _07817_ (.A(_00733_),
    .B(_00735_),
    .C(_00736_),
    .X(_00737_));
 sky130_fd_sc_hd__o21ba_1 _07818_ (.A1(_00735_),
    .A2(_00736_),
    .B1_N(_00733_),
    .X(_00738_));
 sky130_fd_sc_hd__and2_1 _07819_ (.A(_00660_),
    .B(_00661_),
    .X(_00739_));
 sky130_fd_sc_hd__or2_1 _07820_ (.A(_00662_),
    .B(_00739_),
    .X(_00740_));
 sky130_fd_sc_hd__o22a_1 _07821_ (.A1(net24),
    .A2(net113),
    .B1(net110),
    .B2(net22),
    .X(_00741_));
 sky130_fd_sc_hd__xnor2_2 _07822_ (.A(net86),
    .B(_00741_),
    .Y(_00742_));
 sky130_fd_sc_hd__o22a_1 _07823_ (.A1(net149),
    .A2(net21),
    .B1(net19),
    .B2(_00267_),
    .X(_00743_));
 sky130_fd_sc_hd__xnor2_2 _07824_ (.A(net96),
    .B(_00743_),
    .Y(_00744_));
 sky130_fd_sc_hd__and2_1 _07825_ (.A(_00742_),
    .B(_00744_),
    .X(_00745_));
 sky130_fd_sc_hd__o22a_1 _07826_ (.A1(net124),
    .A2(net28),
    .B1(net26),
    .B2(net106),
    .X(_00746_));
 sky130_fd_sc_hd__xnor2_2 _07827_ (.A(net88),
    .B(_00746_),
    .Y(_00747_));
 sky130_fd_sc_hd__xor2_2 _07828_ (.A(_00742_),
    .B(_00744_),
    .X(_00748_));
 sky130_fd_sc_hd__a21o_1 _07829_ (.A1(_00747_),
    .A2(_00748_),
    .B1(_00745_),
    .X(_00749_));
 sky130_fd_sc_hd__or3b_1 _07830_ (.A(_00662_),
    .B(_00739_),
    .C_N(_00749_),
    .X(_00750_));
 sky130_fd_sc_hd__o22a_1 _07831_ (.A1(net39),
    .A2(net152),
    .B1(net151),
    .B2(net37),
    .X(_00751_));
 sky130_fd_sc_hd__xnor2_2 _07832_ (.A(net99),
    .B(_00751_),
    .Y(_00752_));
 sky130_fd_sc_hd__nand2_1 _07833_ (.A(net207),
    .B(net30),
    .Y(_00753_));
 sky130_fd_sc_hd__mux2_1 _07834_ (.A0(_00752_),
    .A1(net92),
    .S(_00753_),
    .X(_00754_));
 sky130_fd_sc_hd__inv_2 _07835_ (.A(_00754_),
    .Y(_00755_));
 sky130_fd_sc_hd__xor2_1 _07836_ (.A(_00740_),
    .B(_00749_),
    .X(_00756_));
 sky130_fd_sc_hd__or2_1 _07837_ (.A(_00755_),
    .B(_00756_),
    .X(_00757_));
 sky130_fd_sc_hd__xnor2_1 _07838_ (.A(_00730_),
    .B(_00738_),
    .Y(_00758_));
 sky130_fd_sc_hd__a21o_1 _07839_ (.A1(_00750_),
    .A2(_00757_),
    .B1(_00758_),
    .X(_00759_));
 sky130_fd_sc_hd__o21ai_2 _07840_ (.A1(_00730_),
    .A2(_00738_),
    .B1(_00759_),
    .Y(_00760_));
 sky130_fd_sc_hd__xor2_2 _07841_ (.A(_00695_),
    .B(_00696_),
    .X(_00761_));
 sky130_fd_sc_hd__xor2_1 _07842_ (.A(_00638_),
    .B(_00639_),
    .X(_00762_));
 sky130_fd_sc_hd__xnor2_1 _07843_ (.A(_00663_),
    .B(_00665_),
    .Y(_00763_));
 sky130_fd_sc_hd__xnor2_1 _07844_ (.A(_00762_),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__xor2_1 _07845_ (.A(_00691_),
    .B(_00694_),
    .X(_00765_));
 sky130_fd_sc_hd__or2_1 _07846_ (.A(_00764_),
    .B(_00765_),
    .X(_00766_));
 sky130_fd_sc_hd__a21bo_1 _07847_ (.A1(_00762_),
    .A2(_00763_),
    .B1_N(_00766_),
    .X(_00767_));
 sky130_fd_sc_hd__xnor2_2 _07848_ (.A(_00760_),
    .B(_00761_),
    .Y(_00768_));
 sky130_fd_sc_hd__nand2b_1 _07849_ (.A_N(_00768_),
    .B(_00767_),
    .Y(_00769_));
 sky130_fd_sc_hd__a21bo_1 _07850_ (.A1(_00760_),
    .A2(_00761_),
    .B1_N(_00769_),
    .X(_00770_));
 sky130_fd_sc_hd__xor2_4 _07851_ (.A(_00571_),
    .B(_00706_),
    .X(_00771_));
 sky130_fd_sc_hd__a21oi_4 _07852_ (.A1(_00770_),
    .A2(_00771_),
    .B1(_00707_),
    .Y(_00772_));
 sky130_fd_sc_hd__a21bo_2 _07853_ (.A1(_00697_),
    .A2(_00703_),
    .B1_N(_00705_),
    .X(_00773_));
 sky130_fd_sc_hd__o21a_2 _07854_ (.A1(_00523_),
    .A2(_00539_),
    .B1(_00538_),
    .X(_00774_));
 sky130_fd_sc_hd__o22a_1 _07855_ (.A1(net28),
    .A2(net120),
    .B1(net115),
    .B2(net26),
    .X(_00775_));
 sky130_fd_sc_hd__xnor2_2 _07856_ (.A(net88),
    .B(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__o22a_1 _07857_ (.A1(net123),
    .A2(net19),
    .B1(net110),
    .B2(net21),
    .X(_00777_));
 sky130_fd_sc_hd__xnor2_1 _07858_ (.A(net96),
    .B(_00777_),
    .Y(_00778_));
 sky130_fd_sc_hd__o22a_1 _07859_ (.A1(net24),
    .A2(net85),
    .B1(_00442_),
    .B2(net22),
    .X(_00779_));
 sky130_fd_sc_hd__xnor2_1 _07860_ (.A(net86),
    .B(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__and2_1 _07861_ (.A(_00778_),
    .B(_00780_),
    .X(_00781_));
 sky130_fd_sc_hd__or2_1 _07862_ (.A(_00778_),
    .B(_00780_),
    .X(_00782_));
 sky130_fd_sc_hd__nand2b_1 _07863_ (.A_N(_00781_),
    .B(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__xnor2_2 _07864_ (.A(_00776_),
    .B(_00783_),
    .Y(_00784_));
 sky130_fd_sc_hd__or2_1 _07865_ (.A(reg1_val[29]),
    .B(net261),
    .X(_00785_));
 sky130_fd_sc_hd__xor2_2 _07866_ (.A(reg1_val[29]),
    .B(_00554_),
    .X(_00786_));
 sky130_fd_sc_hd__o21a_4 _07867_ (.A1(net258),
    .A2(_00786_),
    .B1(_00785_),
    .X(_00787_));
 sky130_fd_sc_hd__o21ai_2 _07868_ (.A1(net258),
    .A2(_00786_),
    .B1(_00785_),
    .Y(_00788_));
 sky130_fd_sc_hd__nand2_1 _07869_ (.A(_00563_),
    .B(net65),
    .Y(_00789_));
 sky130_fd_sc_hd__and3_1 _07870_ (.A(_00564_),
    .B(_00784_),
    .C(_00789_),
    .X(_00790_));
 sky130_fd_sc_hd__a21oi_2 _07871_ (.A1(_00564_),
    .A2(_00789_),
    .B1(_00784_),
    .Y(_00791_));
 sky130_fd_sc_hd__nor2_2 _07872_ (.A(_00790_),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__xnor2_4 _07873_ (.A(_00774_),
    .B(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_1 _07874_ (.A(_00520_),
    .B(_00522_),
    .Y(_00794_));
 sky130_fd_sc_hd__o21a_1 _07875_ (.A1(_00530_),
    .A2(_00536_),
    .B1(_00535_),
    .X(_00795_));
 sky130_fd_sc_hd__nor2_1 _07876_ (.A(_00561_),
    .B(_00787_),
    .Y(_00796_));
 sky130_fd_sc_hd__mux2_2 _07877_ (.A0(_00560_),
    .A1(_00561_),
    .S(net64),
    .X(_00797_));
 sky130_fd_sc_hd__a21o_1 _07878_ (.A1(_00559_),
    .A2(_00787_),
    .B1(_00796_),
    .X(_00798_));
 sky130_fd_sc_hd__a22o_1 _07879_ (.A1(net153),
    .A2(net17),
    .B1(net13),
    .B2(net207),
    .X(_00799_));
 sky130_fd_sc_hd__xnor2_1 _07880_ (.A(net65),
    .B(_00799_),
    .Y(_00800_));
 sky130_fd_sc_hd__nand2b_1 _07881_ (.A_N(_00795_),
    .B(_00800_),
    .Y(_00801_));
 sky130_fd_sc_hd__xnor2_1 _07882_ (.A(_00795_),
    .B(_00800_),
    .Y(_00802_));
 sky130_fd_sc_hd__a21bo_1 _07883_ (.A1(_00520_),
    .A2(_00522_),
    .B1_N(_00802_),
    .X(_00803_));
 sky130_fd_sc_hd__xor2_1 _07884_ (.A(_00794_),
    .B(_00802_),
    .X(_00804_));
 sky130_fd_sc_hd__o22a_1 _07885_ (.A1(net51),
    .A2(net132),
    .B1(net157),
    .B2(net44),
    .X(_00805_));
 sky130_fd_sc_hd__xnor2_2 _07886_ (.A(net202),
    .B(_00805_),
    .Y(_00806_));
 sky130_fd_sc_hd__o22a_1 _07887_ (.A1(net158),
    .A2(net49),
    .B1(net45),
    .B2(net133),
    .X(_00807_));
 sky130_fd_sc_hd__xnor2_1 _07888_ (.A(net179),
    .B(_00807_),
    .Y(_00808_));
 sky130_fd_sc_hd__a211o_4 _07889_ (.A1(_05211_),
    .A2(_00173_),
    .B1(net178),
    .C1(_05123_),
    .X(_00809_));
 sky130_fd_sc_hd__o211ai_4 _07890_ (.A1(net177),
    .A2(_00173_),
    .B1(_00514_),
    .C1(_05123_),
    .Y(_00810_));
 sky130_fd_sc_hd__and2_4 _07891_ (.A(_00809_),
    .B(_00810_),
    .X(_00811_));
 sky130_fd_sc_hd__nand2_8 _07892_ (.A(_00809_),
    .B(_00810_),
    .Y(_00812_));
 sky130_fd_sc_hd__a21o_1 _07893_ (.A1(_00809_),
    .A2(_00810_),
    .B1(net286),
    .X(_00813_));
 sky130_fd_sc_hd__or3_1 _07894_ (.A(net236),
    .B(_00513_),
    .C(_00515_),
    .X(_00814_));
 sky130_fd_sc_hd__nand3_1 _07895_ (.A(net197),
    .B(_00813_),
    .C(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__a21o_1 _07896_ (.A1(_00813_),
    .A2(_00814_),
    .B1(net198),
    .X(_00816_));
 sky130_fd_sc_hd__and3_1 _07897_ (.A(_00808_),
    .B(_00815_),
    .C(_00816_),
    .X(_00817_));
 sky130_fd_sc_hd__a21oi_1 _07898_ (.A1(_00815_),
    .A2(_00816_),
    .B1(_00808_),
    .Y(_00818_));
 sky130_fd_sc_hd__or2_1 _07899_ (.A(_00817_),
    .B(_00818_),
    .X(_00819_));
 sky130_fd_sc_hd__xor2_2 _07900_ (.A(_00806_),
    .B(_00819_),
    .X(_00820_));
 sky130_fd_sc_hd__o22a_1 _07901_ (.A1(net40),
    .A2(_00227_),
    .B1(_00232_),
    .B2(net56),
    .X(_00821_));
 sky130_fd_sc_hd__xor2_2 _07902_ (.A(net154),
    .B(_00821_),
    .X(_00822_));
 sky130_fd_sc_hd__o22a_1 _07903_ (.A1(net100),
    .A2(net68),
    .B1(net66),
    .B2(net42),
    .X(_00823_));
 sky130_fd_sc_hd__xnor2_2 _07904_ (.A(net146),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__o22a_1 _07905_ (.A1(net53),
    .A2(net105),
    .B1(net131),
    .B2(net47),
    .X(_00825_));
 sky130_fd_sc_hd__xnor2_2 _07906_ (.A(net174),
    .B(_00825_),
    .Y(_00826_));
 sky130_fd_sc_hd__nand2_1 _07907_ (.A(_00824_),
    .B(_00826_),
    .Y(_00827_));
 sky130_fd_sc_hd__xnor2_2 _07908_ (.A(_00824_),
    .B(_00826_),
    .Y(_00828_));
 sky130_fd_sc_hd__xnor2_2 _07909_ (.A(_00822_),
    .B(_00828_),
    .Y(_00829_));
 sky130_fd_sc_hd__nor2_1 _07910_ (.A(_00471_),
    .B(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__xor2_2 _07911_ (.A(_00471_),
    .B(_00829_),
    .X(_00831_));
 sky130_fd_sc_hd__xnor2_1 _07912_ (.A(_00820_),
    .B(_00831_),
    .Y(_00832_));
 sky130_fd_sc_hd__a22o_1 _07913_ (.A1(_00266_),
    .A2(net14),
    .B1(net30),
    .B2(_00287_),
    .X(_00833_));
 sky130_fd_sc_hd__xnor2_1 _07914_ (.A(net91),
    .B(_00833_),
    .Y(_00834_));
 sky130_fd_sc_hd__inv_2 _07915_ (.A(_00834_),
    .Y(_00835_));
 sky130_fd_sc_hd__o22a_1 _07916_ (.A1(net35),
    .A2(net151),
    .B1(net149),
    .B2(net33),
    .X(_00836_));
 sky130_fd_sc_hd__xnor2_1 _07917_ (.A(net95),
    .B(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__o22a_1 _07918_ (.A1(net37),
    .A2(_00411_),
    .B1(_00477_),
    .B2(net39),
    .X(_00838_));
 sky130_fd_sc_hd__xnor2_1 _07919_ (.A(net99),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__nand2_1 _07920_ (.A(_00837_),
    .B(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hd__or2_1 _07921_ (.A(_00837_),
    .B(_00839_),
    .X(_00841_));
 sky130_fd_sc_hd__nand2_1 _07922_ (.A(_00840_),
    .B(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__or2_1 _07923_ (.A(_00835_),
    .B(_00842_),
    .X(_00843_));
 sky130_fd_sc_hd__nand2_1 _07924_ (.A(_00835_),
    .B(_00842_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _07925_ (.A(_00843_),
    .B(_00844_),
    .Y(_00845_));
 sky130_fd_sc_hd__nor2_1 _07926_ (.A(_00832_),
    .B(_00845_),
    .Y(_00846_));
 sky130_fd_sc_hd__xor2_1 _07927_ (.A(_00832_),
    .B(_00845_),
    .X(_00847_));
 sky130_fd_sc_hd__nand2_1 _07928_ (.A(_00804_),
    .B(_00847_),
    .Y(_00848_));
 sky130_fd_sc_hd__or2_1 _07929_ (.A(_00804_),
    .B(_00847_),
    .X(_00849_));
 sky130_fd_sc_hd__nand2_2 _07930_ (.A(_00848_),
    .B(_00849_),
    .Y(_00850_));
 sky130_fd_sc_hd__a21bo_2 _07931_ (.A1(_00378_),
    .A2(_00421_),
    .B1_N(_00418_),
    .X(_00851_));
 sky130_fd_sc_hd__a22o_1 _07932_ (.A1(_00220_),
    .A2(_00465_),
    .B1(net71),
    .B2(_00461_),
    .X(_00852_));
 sky130_fd_sc_hd__xnor2_1 _07933_ (.A(_00431_),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__o22a_1 _07934_ (.A1(net83),
    .A2(net76),
    .B1(net74),
    .B2(net79),
    .X(_00854_));
 sky130_fd_sc_hd__xnor2_1 _07935_ (.A(net116),
    .B(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__nand2_1 _07936_ (.A(_00853_),
    .B(_00855_),
    .Y(_00856_));
 sky130_fd_sc_hd__or2_1 _07937_ (.A(_00853_),
    .B(_00855_),
    .X(_00857_));
 sky130_fd_sc_hd__nand2_1 _07938_ (.A(_00856_),
    .B(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__a21oi_1 _07939_ (.A1(_00547_),
    .A2(_00549_),
    .B1(_00858_),
    .Y(_00859_));
 sky130_fd_sc_hd__and3_1 _07940_ (.A(_00547_),
    .B(_00549_),
    .C(_00858_),
    .X(_00860_));
 sky130_fd_sc_hd__or2_2 _07941_ (.A(_00859_),
    .B(_00860_),
    .X(_00861_));
 sky130_fd_sc_hd__and2b_1 _07942_ (.A_N(_00861_),
    .B(_00851_),
    .X(_00862_));
 sky130_fd_sc_hd__xnor2_4 _07943_ (.A(_00851_),
    .B(_00861_),
    .Y(_00863_));
 sky130_fd_sc_hd__xnor2_4 _07944_ (.A(_00850_),
    .B(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__xor2_4 _07945_ (.A(_00793_),
    .B(_00864_),
    .X(_00865_));
 sky130_fd_sc_hd__a21o_2 _07946_ (.A1(_00426_),
    .A2(_00569_),
    .B1(_00568_),
    .X(_00866_));
 sky130_fd_sc_hd__a21o_2 _07947_ (.A1(_00237_),
    .A2(_00425_),
    .B1(_00423_),
    .X(_00867_));
 sky130_fd_sc_hd__or2_2 _07948_ (.A(_00485_),
    .B(_00507_),
    .X(_00868_));
 sky130_fd_sc_hd__a21oi_2 _07949_ (.A1(_00553_),
    .A2(_00566_),
    .B1(_00552_),
    .Y(_00869_));
 sky130_fd_sc_hd__o21ba_1 _07950_ (.A1(_00485_),
    .A2(_00507_),
    .B1_N(_00869_),
    .X(_00870_));
 sky130_fd_sc_hd__xnor2_4 _07951_ (.A(_00868_),
    .B(_00869_),
    .Y(_00871_));
 sky130_fd_sc_hd__xnor2_4 _07952_ (.A(_00867_),
    .B(_00871_),
    .Y(_00872_));
 sky130_fd_sc_hd__a21oi_4 _07953_ (.A1(_00698_),
    .A2(_00702_),
    .B1(_00701_),
    .Y(_00873_));
 sky130_fd_sc_hd__xnor2_4 _07954_ (.A(_00872_),
    .B(_00873_),
    .Y(_00874_));
 sky130_fd_sc_hd__nand2b_1 _07955_ (.A_N(_00874_),
    .B(_00866_),
    .Y(_00875_));
 sky130_fd_sc_hd__xnor2_4 _07956_ (.A(_00866_),
    .B(_00874_),
    .Y(_00876_));
 sky130_fd_sc_hd__and2_1 _07957_ (.A(_00865_),
    .B(_00876_),
    .X(_00877_));
 sky130_fd_sc_hd__xor2_4 _07958_ (.A(_00865_),
    .B(_00876_),
    .X(_00878_));
 sky130_fd_sc_hd__xnor2_4 _07959_ (.A(_00773_),
    .B(_00878_),
    .Y(_00879_));
 sky130_fd_sc_hd__and2_1 _07960_ (.A(_00772_),
    .B(_00879_),
    .X(_00880_));
 sky130_fd_sc_hd__or2_1 _07961_ (.A(_00772_),
    .B(_00879_),
    .X(_00881_));
 sky130_fd_sc_hd__xnor2_4 _07962_ (.A(_00772_),
    .B(_00879_),
    .Y(_00882_));
 sky130_fd_sc_hd__xnor2_2 _07963_ (.A(_00770_),
    .B(_00771_),
    .Y(_00883_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(_00629_),
    .B(_00630_),
    .Y(_00884_));
 sky130_fd_sc_hd__and2_2 _07965_ (.A(_00631_),
    .B(_00884_),
    .X(_00885_));
 sky130_fd_sc_hd__xnor2_2 _07966_ (.A(_00767_),
    .B(_00768_),
    .Y(_00886_));
 sky130_fd_sc_hd__and2_1 _07967_ (.A(_00885_),
    .B(_00886_),
    .X(_00887_));
 sky130_fd_sc_hd__nand3_1 _07968_ (.A(_00750_),
    .B(_00757_),
    .C(_00758_),
    .Y(_00888_));
 sky130_fd_sc_hd__nand2_2 _07969_ (.A(_00759_),
    .B(_00888_),
    .Y(_00889_));
 sky130_fd_sc_hd__xor2_1 _07970_ (.A(_00681_),
    .B(_00683_),
    .X(_00890_));
 sky130_fd_sc_hd__o22a_1 _07971_ (.A1(net85),
    .A2(net68),
    .B1(net66),
    .B2(net82),
    .X(_00891_));
 sky130_fd_sc_hd__xnor2_2 _07972_ (.A(net146),
    .B(_00891_),
    .Y(_00892_));
 sky130_fd_sc_hd__o22a_1 _07973_ (.A1(net131),
    .A2(net103),
    .B1(net70),
    .B2(net104),
    .X(_00893_));
 sky130_fd_sc_hd__xnor2_2 _07974_ (.A(net174),
    .B(_00893_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_1 _07975_ (.A(_00892_),
    .B(_00894_),
    .Y(_00895_));
 sky130_fd_sc_hd__a22o_1 _07976_ (.A1(net128),
    .A2(net78),
    .B1(_00464_),
    .B2(net126),
    .X(_00896_));
 sky130_fd_sc_hd__xnor2_2 _07977_ (.A(net154),
    .B(_00896_),
    .Y(_00897_));
 sky130_fd_sc_hd__xnor2_2 _07978_ (.A(_00892_),
    .B(_00894_),
    .Y(_00898_));
 sky130_fd_sc_hd__o21a_1 _07979_ (.A1(_00897_),
    .A2(_00898_),
    .B1(_00895_),
    .X(_00899_));
 sky130_fd_sc_hd__and2b_1 _07980_ (.A_N(_00899_),
    .B(_00890_),
    .X(_00900_));
 sky130_fd_sc_hd__a22o_1 _07981_ (.A1(_06726_),
    .A2(_00203_),
    .B1(_00229_),
    .B2(_06702_),
    .X(_00901_));
 sky130_fd_sc_hd__xnor2_2 _07982_ (.A(net181),
    .B(_00901_),
    .Y(_00902_));
 sky130_fd_sc_hd__o22a_1 _07983_ (.A1(net53),
    .A2(net236),
    .B1(net47),
    .B2(net286),
    .X(_00903_));
 sky130_fd_sc_hd__xnor2_2 _07984_ (.A(net199),
    .B(_00903_),
    .Y(_00904_));
 sky130_fd_sc_hd__and2_1 _07985_ (.A(_00902_),
    .B(_00904_),
    .X(_00905_));
 sky130_fd_sc_hd__o22a_2 _07986_ (.A1(net56),
    .A2(_00160_),
    .B1(net40),
    .B2(net132),
    .X(_00906_));
 sky130_fd_sc_hd__xnor2_4 _07987_ (.A(net200),
    .B(_00906_),
    .Y(_00907_));
 sky130_fd_sc_hd__or2_1 _07988_ (.A(_00902_),
    .B(_00904_),
    .X(_00908_));
 sky130_fd_sc_hd__xnor2_2 _07989_ (.A(_00902_),
    .B(_00904_),
    .Y(_00909_));
 sky130_fd_sc_hd__a21o_1 _07990_ (.A1(_00907_),
    .A2(_00908_),
    .B1(_00905_),
    .X(_00910_));
 sky130_fd_sc_hd__xnor2_1 _07991_ (.A(_00890_),
    .B(_00899_),
    .Y(_00911_));
 sky130_fd_sc_hd__a21o_1 _07992_ (.A1(_00910_),
    .A2(_00911_),
    .B1(_00900_),
    .X(_00912_));
 sky130_fd_sc_hd__xnor2_2 _07993_ (.A(_00715_),
    .B(_00716_),
    .Y(_00913_));
 sky130_fd_sc_hd__xor2_2 _07994_ (.A(_00752_),
    .B(_00753_),
    .X(_00914_));
 sky130_fd_sc_hd__or2_1 _07995_ (.A(_00913_),
    .B(_00914_),
    .X(_00915_));
 sky130_fd_sc_hd__xnor2_2 _07996_ (.A(_00747_),
    .B(_00748_),
    .Y(_00916_));
 sky130_fd_sc_hd__xnor2_2 _07997_ (.A(_00913_),
    .B(_00914_),
    .Y(_00917_));
 sky130_fd_sc_hd__o21ai_2 _07998_ (.A1(_00916_),
    .A2(_00917_),
    .B1(_00915_),
    .Y(_00918_));
 sky130_fd_sc_hd__o22a_1 _07999_ (.A1(net22),
    .A2(net113),
    .B1(net106),
    .B2(net24),
    .X(_00919_));
 sky130_fd_sc_hd__xnor2_1 _08000_ (.A(_00359_),
    .B(_00919_),
    .Y(_00920_));
 sky130_fd_sc_hd__o22a_1 _08001_ (.A1(net119),
    .A2(net75),
    .B1(net72),
    .B2(net115),
    .X(_00921_));
 sky130_fd_sc_hd__xnor2_1 _08002_ (.A(_00431_),
    .B(_00921_),
    .Y(_00922_));
 sky130_fd_sc_hd__or2_1 _08003_ (.A(_00920_),
    .B(_00922_),
    .X(_00923_));
 sky130_fd_sc_hd__o22a_1 _08004_ (.A1(net110),
    .A2(net84),
    .B1(net80),
    .B2(net123),
    .X(_00924_));
 sky130_fd_sc_hd__xnor2_1 _08005_ (.A(_00381_),
    .B(_00924_),
    .Y(_00925_));
 sky130_fd_sc_hd__xnor2_1 _08006_ (.A(_00920_),
    .B(_00922_),
    .Y(_00926_));
 sky130_fd_sc_hd__o21a_1 _08007_ (.A1(_00925_),
    .A2(_00926_),
    .B1(_00923_),
    .X(_00927_));
 sky130_fd_sc_hd__xnor2_1 _08008_ (.A(_00725_),
    .B(_00727_),
    .Y(_00928_));
 sky130_fd_sc_hd__and2b_1 _08009_ (.A_N(_00927_),
    .B(_00928_),
    .X(_00929_));
 sky130_fd_sc_hd__o22a_1 _08010_ (.A1(_00267_),
    .A2(net28),
    .B1(net26),
    .B2(net124),
    .X(_00930_));
 sky130_fd_sc_hd__xnor2_1 _08011_ (.A(net88),
    .B(_00930_),
    .Y(_00931_));
 sky130_fd_sc_hd__o22a_1 _08012_ (.A1(net151),
    .A2(net21),
    .B1(net19),
    .B2(net149),
    .X(_00932_));
 sky130_fd_sc_hd__xnor2_1 _08013_ (.A(net96),
    .B(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(_00931_),
    .B(_00933_),
    .Y(_00934_));
 sky130_fd_sc_hd__inv_2 _08015_ (.A(_00934_),
    .Y(_00935_));
 sky130_fd_sc_hd__xnor2_1 _08016_ (.A(_00927_),
    .B(_00928_),
    .Y(_00936_));
 sky130_fd_sc_hd__a21oi_1 _08017_ (.A1(_00935_),
    .A2(_00936_),
    .B1(_00929_),
    .Y(_00937_));
 sky130_fd_sc_hd__xor2_1 _08018_ (.A(_00912_),
    .B(_00918_),
    .X(_00938_));
 sky130_fd_sc_hd__and2b_1 _08019_ (.A_N(_00937_),
    .B(_00938_),
    .X(_00939_));
 sky130_fd_sc_hd__a21oi_2 _08020_ (.A1(_00912_),
    .A2(_00918_),
    .B1(_00939_),
    .Y(_00940_));
 sky130_fd_sc_hd__or3_1 _08021_ (.A(_00718_),
    .B(_00723_),
    .C(_00728_),
    .X(_00941_));
 sky130_fd_sc_hd__and2_1 _08022_ (.A(_00729_),
    .B(_00941_),
    .X(_00942_));
 sky130_fd_sc_hd__o21ai_1 _08023_ (.A1(_00733_),
    .A2(_00736_),
    .B1(_00735_),
    .Y(_00943_));
 sky130_fd_sc_hd__and3_1 _08024_ (.A(_00737_),
    .B(_00942_),
    .C(_00943_),
    .X(_00944_));
 sky130_fd_sc_hd__a21oi_1 _08025_ (.A1(_00737_),
    .A2(_00943_),
    .B1(_00942_),
    .Y(_00945_));
 sky130_fd_sc_hd__nor2_1 _08026_ (.A(_00944_),
    .B(_00945_),
    .Y(_00946_));
 sky130_fd_sc_hd__nand2_1 _08027_ (.A(_00755_),
    .B(_00756_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _08028_ (.A(_00757_),
    .B(_00947_),
    .Y(_00948_));
 sky130_fd_sc_hd__a31o_1 _08029_ (.A1(_00757_),
    .A2(_00946_),
    .A3(_00947_),
    .B1(_00944_),
    .X(_00949_));
 sky130_fd_sc_hd__xnor2_1 _08030_ (.A(_00889_),
    .B(_00940_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand2b_1 _08031_ (.A_N(_00950_),
    .B(_00949_),
    .Y(_00951_));
 sky130_fd_sc_hd__o21ai_4 _08032_ (.A1(_00889_),
    .A2(_00940_),
    .B1(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__xor2_4 _08033_ (.A(_00885_),
    .B(_00886_),
    .X(_00953_));
 sky130_fd_sc_hd__a21oi_2 _08034_ (.A1(_00952_),
    .A2(_00953_),
    .B1(_00887_),
    .Y(_00954_));
 sky130_fd_sc_hd__and2_1 _08035_ (.A(_00883_),
    .B(_00954_),
    .X(_00955_));
 sky130_fd_sc_hd__nand2_1 _08036_ (.A(_00764_),
    .B(_00765_),
    .Y(_00956_));
 sky130_fd_sc_hd__and2_1 _08037_ (.A(_00766_),
    .B(_00956_),
    .X(_00957_));
 sky130_fd_sc_hd__xnor2_1 _08038_ (.A(_00949_),
    .B(_00950_),
    .Y(_00958_));
 sky130_fd_sc_hd__xor2_1 _08039_ (.A(_00937_),
    .B(_00938_),
    .X(_00959_));
 sky130_fd_sc_hd__xnor2_1 _08040_ (.A(_00931_),
    .B(_00933_),
    .Y(_00960_));
 sky130_fd_sc_hd__xnor2_2 _08041_ (.A(_00897_),
    .B(_00898_),
    .Y(_00961_));
 sky130_fd_sc_hd__or2_1 _08042_ (.A(_00960_),
    .B(_00961_),
    .X(_00962_));
 sky130_fd_sc_hd__xnor2_1 _08043_ (.A(_00960_),
    .B(_00961_),
    .Y(_00963_));
 sky130_fd_sc_hd__xnor2_1 _08044_ (.A(_00925_),
    .B(_00926_),
    .Y(_00964_));
 sky130_fd_sc_hd__o21a_1 _08045_ (.A1(_00963_),
    .A2(_00964_),
    .B1(_00962_),
    .X(_00965_));
 sky130_fd_sc_hd__o22a_1 _08046_ (.A1(net105),
    .A2(net74),
    .B1(net70),
    .B2(net131),
    .X(_00966_));
 sky130_fd_sc_hd__xnor2_1 _08047_ (.A(net174),
    .B(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__o22a_1 _08048_ (.A1(net115),
    .A2(net68),
    .B1(net66),
    .B2(net85),
    .X(_00968_));
 sky130_fd_sc_hd__xnor2_1 _08049_ (.A(net146),
    .B(_00968_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_1 _08050_ (.A(_00967_),
    .B(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__o22a_1 _08051_ (.A1(_00227_),
    .A2(net82),
    .B1(net76),
    .B2(_00232_),
    .X(_00971_));
 sky130_fd_sc_hd__xnor2_1 _08052_ (.A(net154),
    .B(_00971_),
    .Y(_00972_));
 sky130_fd_sc_hd__inv_2 _08053_ (.A(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__xnor2_1 _08054_ (.A(_00967_),
    .B(_00969_),
    .Y(_00974_));
 sky130_fd_sc_hd__o21ai_1 _08055_ (.A1(_00973_),
    .A2(_00974_),
    .B1(_00970_),
    .Y(_00975_));
 sky130_fd_sc_hd__o22a_1 _08056_ (.A1(net212),
    .A2(net39),
    .B1(net37),
    .B2(net152),
    .X(_00976_));
 sky130_fd_sc_hd__xnor2_1 _08057_ (.A(net99),
    .B(_00976_),
    .Y(_00977_));
 sky130_fd_sc_hd__nand2_1 _08058_ (.A(_00975_),
    .B(_00977_),
    .Y(_00978_));
 sky130_fd_sc_hd__o22a_1 _08059_ (.A1(net133),
    .A2(net103),
    .B1(net100),
    .B2(net158),
    .X(_00979_));
 sky130_fd_sc_hd__xnor2_2 _08060_ (.A(net179),
    .B(_00979_),
    .Y(_00980_));
 sky130_fd_sc_hd__a22o_1 _08061_ (.A1(net292),
    .A2(_06730_),
    .B1(_00138_),
    .B2(_06725_),
    .X(_00981_));
 sky130_fd_sc_hd__xnor2_2 _08062_ (.A(net198),
    .B(_00981_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_1 _08063_ (.A(_00980_),
    .B(_00982_),
    .Y(_00983_));
 sky130_fd_sc_hd__xnor2_2 _08064_ (.A(_00980_),
    .B(_00982_),
    .Y(_00984_));
 sky130_fd_sc_hd__o22a_1 _08065_ (.A1(net132),
    .A2(net42),
    .B1(net40),
    .B2(_00160_),
    .X(_00985_));
 sky130_fd_sc_hd__xnor2_1 _08066_ (.A(net201),
    .B(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hd__o21ai_2 _08067_ (.A1(_00984_),
    .A2(_00986_),
    .B1(_00983_),
    .Y(_00987_));
 sky130_fd_sc_hd__xor2_1 _08068_ (.A(_00975_),
    .B(_00977_),
    .X(_00988_));
 sky130_fd_sc_hd__a21boi_2 _08069_ (.A1(_00987_),
    .A2(_00988_),
    .B1_N(_00978_),
    .Y(_00989_));
 sky130_fd_sc_hd__nor2_1 _08070_ (.A(_00965_),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__xnor2_4 _08071_ (.A(_00907_),
    .B(_00909_),
    .Y(_00991_));
 sky130_fd_sc_hd__o22a_1 _08072_ (.A1(net124),
    .A2(net24),
    .B1(net22),
    .B2(net106),
    .X(_00992_));
 sky130_fd_sc_hd__xnor2_1 _08073_ (.A(_00359_),
    .B(_00992_),
    .Y(_00993_));
 sky130_fd_sc_hd__o22a_1 _08074_ (.A1(net123),
    .A2(net75),
    .B1(net72),
    .B2(net119),
    .X(_00994_));
 sky130_fd_sc_hd__xnor2_1 _08075_ (.A(_00431_),
    .B(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__or2_1 _08076_ (.A(_00993_),
    .B(_00995_),
    .X(_00996_));
 sky130_fd_sc_hd__o22a_1 _08077_ (.A1(net113),
    .A2(net84),
    .B1(net80),
    .B2(net110),
    .X(_00997_));
 sky130_fd_sc_hd__xnor2_1 _08078_ (.A(net116),
    .B(_00997_),
    .Y(_00998_));
 sky130_fd_sc_hd__inv_2 _08079_ (.A(_00998_),
    .Y(_00999_));
 sky130_fd_sc_hd__xnor2_1 _08080_ (.A(_00993_),
    .B(_00995_),
    .Y(_01000_));
 sky130_fd_sc_hd__o21a_1 _08081_ (.A1(_00999_),
    .A2(_01000_),
    .B1(_00996_),
    .X(_01001_));
 sky130_fd_sc_hd__and2b_1 _08082_ (.A_N(_01001_),
    .B(_00991_),
    .X(_01002_));
 sky130_fd_sc_hd__o22a_1 _08083_ (.A1(net152),
    .A2(net21),
    .B1(net19),
    .B2(_00326_),
    .X(_01003_));
 sky130_fd_sc_hd__xnor2_2 _08084_ (.A(net96),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__o22a_1 _08085_ (.A1(_00339_),
    .A2(net28),
    .B1(net26),
    .B2(net125),
    .X(_01005_));
 sky130_fd_sc_hd__xnor2_2 _08086_ (.A(net88),
    .B(_01005_),
    .Y(_01006_));
 sky130_fd_sc_hd__nand2_1 _08087_ (.A(_01004_),
    .B(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hd__xnor2_2 _08088_ (.A(_00991_),
    .B(_01001_),
    .Y(_01008_));
 sky130_fd_sc_hd__a31o_1 _08089_ (.A1(_01004_),
    .A2(_01006_),
    .A3(_01008_),
    .B1(_01002_),
    .X(_01009_));
 sky130_fd_sc_hd__xor2_2 _08090_ (.A(_00965_),
    .B(_00989_),
    .X(_01010_));
 sky130_fd_sc_hd__a21oi_2 _08091_ (.A1(_01009_),
    .A2(_01010_),
    .B1(_00990_),
    .Y(_01011_));
 sky130_fd_sc_hd__xnor2_1 _08092_ (.A(_00910_),
    .B(_00911_),
    .Y(_01012_));
 sky130_fd_sc_hd__xor2_2 _08093_ (.A(_00916_),
    .B(_00917_),
    .X(_01013_));
 sky130_fd_sc_hd__and2b_1 _08094_ (.A_N(_01012_),
    .B(_01013_),
    .X(_01014_));
 sky130_fd_sc_hd__xnor2_1 _08095_ (.A(_00934_),
    .B(_00936_),
    .Y(_01015_));
 sky130_fd_sc_hd__xnor2_1 _08096_ (.A(_01012_),
    .B(_01013_),
    .Y(_01016_));
 sky130_fd_sc_hd__a21o_1 _08097_ (.A1(_01015_),
    .A2(_01016_),
    .B1(_01014_),
    .X(_01017_));
 sky130_fd_sc_hd__xnor2_1 _08098_ (.A(_00959_),
    .B(_01011_),
    .Y(_01018_));
 sky130_fd_sc_hd__nand2b_1 _08099_ (.A_N(_01018_),
    .B(_01017_),
    .Y(_01019_));
 sky130_fd_sc_hd__o21ai_1 _08100_ (.A1(_00959_),
    .A2(_01011_),
    .B1(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__xnor2_1 _08101_ (.A(_00957_),
    .B(_00958_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2b_1 _08102_ (.A_N(_01021_),
    .B(_01020_),
    .Y(_01022_));
 sky130_fd_sc_hd__a21bo_2 _08103_ (.A1(_00957_),
    .A2(_00958_),
    .B1_N(_01022_),
    .X(_01023_));
 sky130_fd_sc_hd__xor2_4 _08104_ (.A(_00952_),
    .B(_00953_),
    .X(_01024_));
 sky130_fd_sc_hd__nand2_1 _08105_ (.A(_01023_),
    .B(_01024_),
    .Y(_01025_));
 sky130_fd_sc_hd__or2_1 _08106_ (.A(_00883_),
    .B(_00954_),
    .X(_01026_));
 sky130_fd_sc_hd__a21o_1 _08107_ (.A1(_01025_),
    .A2(_01026_),
    .B1(_00955_),
    .X(_01027_));
 sky130_fd_sc_hd__xnor2_1 _08108_ (.A(_00946_),
    .B(_00948_),
    .Y(_01028_));
 sky130_fd_sc_hd__xnor2_1 _08109_ (.A(_01017_),
    .B(_01018_),
    .Y(_01029_));
 sky130_fd_sc_hd__nand2_1 _08110_ (.A(_01028_),
    .B(_01029_),
    .Y(_01030_));
 sky130_fd_sc_hd__xnor2_2 _08111_ (.A(_01009_),
    .B(_01010_),
    .Y(_01031_));
 sky130_fd_sc_hd__xnor2_1 _08112_ (.A(_01004_),
    .B(_01006_),
    .Y(_01032_));
 sky130_fd_sc_hd__xnor2_1 _08113_ (.A(_00973_),
    .B(_00974_),
    .Y(_01033_));
 sky130_fd_sc_hd__nor2_1 _08114_ (.A(_01032_),
    .B(_01033_),
    .Y(_01034_));
 sky130_fd_sc_hd__xnor2_1 _08115_ (.A(_00998_),
    .B(_01000_),
    .Y(_01035_));
 sky130_fd_sc_hd__xor2_1 _08116_ (.A(_01032_),
    .B(_01033_),
    .X(_01036_));
 sky130_fd_sc_hd__a21oi_2 _08117_ (.A1(_01035_),
    .A2(_01036_),
    .B1(_01034_),
    .Y(_01037_));
 sky130_fd_sc_hd__nor2_1 _08118_ (.A(net212),
    .B(net37),
    .Y(_01038_));
 sky130_fd_sc_hd__a22o_1 _08119_ (.A1(_06726_),
    .A2(_00220_),
    .B1(net71),
    .B2(_06702_),
    .X(_01039_));
 sky130_fd_sc_hd__xnor2_1 _08120_ (.A(net179),
    .B(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__a21o_1 _08121_ (.A1(_06722_),
    .A2(_06723_),
    .B1(net285),
    .X(_01041_));
 sky130_fd_sc_hd__or3_1 _08122_ (.A(net236),
    .B(_00206_),
    .C(_00207_),
    .X(_01042_));
 sky130_fd_sc_hd__and3_1 _08123_ (.A(net198),
    .B(_01041_),
    .C(_01042_),
    .X(_01043_));
 sky130_fd_sc_hd__a21oi_1 _08124_ (.A1(_01041_),
    .A2(_01042_),
    .B1(net198),
    .Y(_01044_));
 sky130_fd_sc_hd__or3_1 _08125_ (.A(_01040_),
    .B(_01043_),
    .C(_01044_),
    .X(_01045_));
 sky130_fd_sc_hd__o21ai_1 _08126_ (.A1(_01043_),
    .A2(_01044_),
    .B1(_01040_),
    .Y(_01046_));
 sky130_fd_sc_hd__a22o_1 _08127_ (.A1(_00159_),
    .A2(_00203_),
    .B1(_00229_),
    .B2(_00158_),
    .X(_01047_));
 sky130_fd_sc_hd__xnor2_1 _08128_ (.A(net202),
    .B(_01047_),
    .Y(_01048_));
 sky130_fd_sc_hd__nand3_1 _08129_ (.A(_01045_),
    .B(_01046_),
    .C(_01048_),
    .Y(_01049_));
 sky130_fd_sc_hd__nand2_1 _08130_ (.A(_01045_),
    .B(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__mux2_1 _08131_ (.A0(net99),
    .A1(_01050_),
    .S(_01038_),
    .X(_01051_));
 sky130_fd_sc_hd__and2b_1 _08132_ (.A_N(_01037_),
    .B(_01051_),
    .X(_01052_));
 sky130_fd_sc_hd__xnor2_1 _08133_ (.A(_00984_),
    .B(_00986_),
    .Y(_01053_));
 sky130_fd_sc_hd__o22a_1 _08134_ (.A1(net119),
    .A2(net69),
    .B1(net67),
    .B2(net115),
    .X(_01054_));
 sky130_fd_sc_hd__xnor2_1 _08135_ (.A(net147),
    .B(_01054_),
    .Y(_01055_));
 sky130_fd_sc_hd__o22a_1 _08136_ (.A1(net104),
    .A2(net76),
    .B1(net74),
    .B2(net130),
    .X(_01056_));
 sky130_fd_sc_hd__xnor2_1 _08137_ (.A(net175),
    .B(_01056_),
    .Y(_01057_));
 sky130_fd_sc_hd__a22o_1 _08138_ (.A1(net128),
    .A2(_00397_),
    .B1(net81),
    .B2(net126),
    .X(_01058_));
 sky130_fd_sc_hd__xnor2_1 _08139_ (.A(net154),
    .B(_01058_),
    .Y(_01059_));
 sky130_fd_sc_hd__xnor2_1 _08140_ (.A(_01055_),
    .B(_01057_),
    .Y(_01060_));
 sky130_fd_sc_hd__or2_1 _08141_ (.A(_01059_),
    .B(_01060_),
    .X(_01061_));
 sky130_fd_sc_hd__a21bo_1 _08142_ (.A1(_01055_),
    .A2(_01057_),
    .B1_N(_01061_),
    .X(_01062_));
 sky130_fd_sc_hd__and2b_1 _08143_ (.A_N(_01053_),
    .B(_01062_),
    .X(_01063_));
 sky130_fd_sc_hd__a22o_1 _08144_ (.A1(net111),
    .A2(_00461_),
    .B1(_00465_),
    .B2(_00372_),
    .X(_01064_));
 sky130_fd_sc_hd__xnor2_1 _08145_ (.A(_00431_),
    .B(_01064_),
    .Y(_01065_));
 sky130_fd_sc_hd__o22a_1 _08146_ (.A1(net113),
    .A2(net80),
    .B1(net106),
    .B2(net84),
    .X(_01066_));
 sky130_fd_sc_hd__xnor2_1 _08147_ (.A(net116),
    .B(_01066_),
    .Y(_01067_));
 sky130_fd_sc_hd__nand2_1 _08148_ (.A(_01065_),
    .B(_01067_),
    .Y(_01068_));
 sky130_fd_sc_hd__inv_2 _08149_ (.A(_01068_),
    .Y(_01069_));
 sky130_fd_sc_hd__xnor2_1 _08150_ (.A(_01053_),
    .B(_01062_),
    .Y(_01070_));
 sky130_fd_sc_hd__a21o_1 _08151_ (.A1(_01069_),
    .A2(_01070_),
    .B1(_01063_),
    .X(_01071_));
 sky130_fd_sc_hd__xnor2_2 _08152_ (.A(_01037_),
    .B(_01051_),
    .Y(_01072_));
 sky130_fd_sc_hd__a21oi_1 _08153_ (.A1(_01071_),
    .A2(_01072_),
    .B1(_01052_),
    .Y(_01073_));
 sky130_fd_sc_hd__nor2_1 _08154_ (.A(_01031_),
    .B(_01073_),
    .Y(_01074_));
 sky130_fd_sc_hd__xnor2_1 _08155_ (.A(_00963_),
    .B(_00964_),
    .Y(_01075_));
 sky130_fd_sc_hd__xnor2_1 _08156_ (.A(_00987_),
    .B(_00988_),
    .Y(_01076_));
 sky130_fd_sc_hd__nor2_1 _08157_ (.A(_01075_),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__nand2_1 _08158_ (.A(_01075_),
    .B(_01076_),
    .Y(_01078_));
 sky130_fd_sc_hd__and2b_1 _08159_ (.A_N(_01077_),
    .B(_01078_),
    .X(_01079_));
 sky130_fd_sc_hd__xnor2_2 _08160_ (.A(_01007_),
    .B(_01008_),
    .Y(_01080_));
 sky130_fd_sc_hd__a21o_1 _08161_ (.A1(_01078_),
    .A2(_01080_),
    .B1(_01077_),
    .X(_01081_));
 sky130_fd_sc_hd__xnor2_1 _08162_ (.A(_01031_),
    .B(_01073_),
    .Y(_01082_));
 sky130_fd_sc_hd__and2b_1 _08163_ (.A_N(_01082_),
    .B(_01081_),
    .X(_01083_));
 sky130_fd_sc_hd__xor2_1 _08164_ (.A(_01028_),
    .B(_01029_),
    .X(_01084_));
 sky130_fd_sc_hd__o21ai_1 _08165_ (.A1(_01074_),
    .A2(_01083_),
    .B1(_01084_),
    .Y(_01085_));
 sky130_fd_sc_hd__xor2_1 _08166_ (.A(_01020_),
    .B(_01021_),
    .X(_01086_));
 sky130_fd_sc_hd__and3_1 _08167_ (.A(_01030_),
    .B(_01085_),
    .C(_01086_),
    .X(_01087_));
 sky130_fd_sc_hd__xnor2_1 _08168_ (.A(_01015_),
    .B(_01016_),
    .Y(_01088_));
 sky130_fd_sc_hd__xor2_1 _08169_ (.A(_01081_),
    .B(_01082_),
    .X(_01089_));
 sky130_fd_sc_hd__or2_1 _08170_ (.A(_01088_),
    .B(_01089_),
    .X(_01090_));
 sky130_fd_sc_hd__a21o_1 _08171_ (.A1(_01045_),
    .A2(_01046_),
    .B1(_01048_),
    .X(_01091_));
 sky130_fd_sc_hd__or2_1 _08172_ (.A(_01065_),
    .B(_01067_),
    .X(_01092_));
 sky130_fd_sc_hd__and2_1 _08173_ (.A(_01068_),
    .B(_01092_),
    .X(_01093_));
 sky130_fd_sc_hd__and3_1 _08174_ (.A(_01049_),
    .B(_01091_),
    .C(_01093_),
    .X(_01094_));
 sky130_fd_sc_hd__a21oi_2 _08175_ (.A1(_01049_),
    .A2(_01091_),
    .B1(_01093_),
    .Y(_01095_));
 sky130_fd_sc_hd__nand2_1 _08176_ (.A(_01059_),
    .B(_01060_),
    .Y(_01096_));
 sky130_fd_sc_hd__nand2_1 _08177_ (.A(_01061_),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__or3_1 _08178_ (.A(_01094_),
    .B(_01095_),
    .C(_01097_),
    .X(_01098_));
 sky130_fd_sc_hd__o21bai_2 _08179_ (.A1(_01095_),
    .A2(_01097_),
    .B1_N(_01094_),
    .Y(_01099_));
 sky130_fd_sc_hd__o22a_1 _08180_ (.A1(net125),
    .A2(net24),
    .B1(net22),
    .B2(net124),
    .X(_01100_));
 sky130_fd_sc_hd__xnor2_1 _08181_ (.A(net86),
    .B(_01100_),
    .Y(_01101_));
 sky130_fd_sc_hd__o22a_1 _08182_ (.A1(net209),
    .A2(net21),
    .B1(net19),
    .B2(net152),
    .X(_01102_));
 sky130_fd_sc_hd__xnor2_1 _08183_ (.A(net96),
    .B(_01102_),
    .Y(_01103_));
 sky130_fd_sc_hd__o22a_1 _08184_ (.A1(net151),
    .A2(net28),
    .B1(net26),
    .B2(net149),
    .X(_01104_));
 sky130_fd_sc_hd__xor2_1 _08185_ (.A(net88),
    .B(_01104_),
    .X(_01105_));
 sky130_fd_sc_hd__xnor2_1 _08186_ (.A(_01101_),
    .B(_01103_),
    .Y(_01106_));
 sky130_fd_sc_hd__nor2_1 _08187_ (.A(_01105_),
    .B(_01106_),
    .Y(_01107_));
 sky130_fd_sc_hd__a21o_1 _08188_ (.A1(_01101_),
    .A2(_01103_),
    .B1(_01107_),
    .X(_01108_));
 sky130_fd_sc_hd__and2_1 _08189_ (.A(_01099_),
    .B(_01108_),
    .X(_01109_));
 sky130_fd_sc_hd__o22a_1 _08190_ (.A1(net124),
    .A2(net84),
    .B1(net80),
    .B2(net106),
    .X(_01110_));
 sky130_fd_sc_hd__xnor2_1 _08191_ (.A(net116),
    .B(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__a22o_1 _08192_ (.A1(_00412_),
    .A2(_00461_),
    .B1(_00465_),
    .B2(net111),
    .X(_01112_));
 sky130_fd_sc_hd__xnor2_1 _08193_ (.A(_00431_),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__nand2_1 _08194_ (.A(_01111_),
    .B(_01113_),
    .Y(_01114_));
 sky130_fd_sc_hd__a22o_1 _08195_ (.A1(_06702_),
    .A2(_00464_),
    .B1(net71),
    .B2(_06726_),
    .X(_01115_));
 sky130_fd_sc_hd__xnor2_1 _08196_ (.A(net181),
    .B(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__or3_1 _08197_ (.A(net285),
    .B(_00206_),
    .C(_00207_),
    .X(_01117_));
 sky130_fd_sc_hd__a21o_1 _08198_ (.A1(_00200_),
    .A2(_00201_),
    .B1(net236),
    .X(_01118_));
 sky130_fd_sc_hd__nand3_1 _08199_ (.A(net198),
    .B(_01117_),
    .C(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__a21o_1 _08200_ (.A1(_01117_),
    .A2(_01118_),
    .B1(net198),
    .X(_01120_));
 sky130_fd_sc_hd__nand3_1 _08201_ (.A(_01116_),
    .B(_01119_),
    .C(_01120_),
    .Y(_01121_));
 sky130_fd_sc_hd__o22a_1 _08202_ (.A1(_00157_),
    .A2(net103),
    .B1(net100),
    .B2(_00160_),
    .X(_01122_));
 sky130_fd_sc_hd__xnor2_1 _08203_ (.A(_06694_),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__a21o_1 _08204_ (.A1(_01119_),
    .A2(_01120_),
    .B1(_01116_),
    .X(_01124_));
 sky130_fd_sc_hd__nand3_1 _08205_ (.A(_01121_),
    .B(_01123_),
    .C(_01124_),
    .Y(_01125_));
 sky130_fd_sc_hd__a21boi_2 _08206_ (.A1(_01123_),
    .A2(_01124_),
    .B1_N(_01121_),
    .Y(_01126_));
 sky130_fd_sc_hd__o22a_1 _08207_ (.A1(net104),
    .A2(net82),
    .B1(net76),
    .B2(net130),
    .X(_01127_));
 sky130_fd_sc_hd__xnor2_2 _08208_ (.A(net175),
    .B(_01127_),
    .Y(_01128_));
 sky130_fd_sc_hd__o22a_1 _08209_ (.A1(net123),
    .A2(net69),
    .B1(net67),
    .B2(net119),
    .X(_01129_));
 sky130_fd_sc_hd__xnor2_2 _08210_ (.A(net147),
    .B(_01129_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _08211_ (.A(_01128_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__a22o_1 _08212_ (.A1(net128),
    .A2(net114),
    .B1(_00397_),
    .B2(net126),
    .X(_01132_));
 sky130_fd_sc_hd__xor2_2 _08213_ (.A(net156),
    .B(_01132_),
    .X(_01133_));
 sky130_fd_sc_hd__xnor2_2 _08214_ (.A(_01128_),
    .B(_01130_),
    .Y(_01134_));
 sky130_fd_sc_hd__inv_2 _08215_ (.A(_01134_),
    .Y(_01135_));
 sky130_fd_sc_hd__nand2_1 _08216_ (.A(_01133_),
    .B(_01135_),
    .Y(_01136_));
 sky130_fd_sc_hd__xnor2_1 _08217_ (.A(_01114_),
    .B(_01126_),
    .Y(_01137_));
 sky130_fd_sc_hd__a21oi_1 _08218_ (.A1(_01131_),
    .A2(_01136_),
    .B1(_01137_),
    .Y(_01138_));
 sky130_fd_sc_hd__o21bai_2 _08219_ (.A1(_01114_),
    .A2(_01126_),
    .B1_N(_01138_),
    .Y(_01139_));
 sky130_fd_sc_hd__xor2_2 _08220_ (.A(_01099_),
    .B(_01108_),
    .X(_01140_));
 sky130_fd_sc_hd__a21o_1 _08221_ (.A1(_01139_),
    .A2(_01140_),
    .B1(_01109_),
    .X(_01141_));
 sky130_fd_sc_hd__xor2_2 _08222_ (.A(_01071_),
    .B(_01072_),
    .X(_01142_));
 sky130_fd_sc_hd__xor2_1 _08223_ (.A(_01035_),
    .B(_01036_),
    .X(_01143_));
 sky130_fd_sc_hd__xor2_1 _08224_ (.A(_01038_),
    .B(_01050_),
    .X(_01144_));
 sky130_fd_sc_hd__xnor2_1 _08225_ (.A(_01069_),
    .B(_01070_),
    .Y(_01145_));
 sky130_fd_sc_hd__xnor2_1 _08226_ (.A(_01143_),
    .B(_01144_),
    .Y(_01146_));
 sky130_fd_sc_hd__or2_1 _08227_ (.A(_01145_),
    .B(_01146_),
    .X(_01147_));
 sky130_fd_sc_hd__a21bo_1 _08228_ (.A1(_01143_),
    .A2(_01144_),
    .B1_N(_01147_),
    .X(_01148_));
 sky130_fd_sc_hd__xnor2_2 _08229_ (.A(_01141_),
    .B(_01142_),
    .Y(_01149_));
 sky130_fd_sc_hd__and2b_1 _08230_ (.A_N(_01149_),
    .B(_01148_),
    .X(_01150_));
 sky130_fd_sc_hd__a21o_1 _08231_ (.A1(_01141_),
    .A2(_01142_),
    .B1(_01150_),
    .X(_01151_));
 sky130_fd_sc_hd__xor2_1 _08232_ (.A(_01088_),
    .B(_01089_),
    .X(_01152_));
 sky130_fd_sc_hd__nand2_1 _08233_ (.A(_01151_),
    .B(_01152_),
    .Y(_01153_));
 sky130_fd_sc_hd__or3_1 _08234_ (.A(_01074_),
    .B(_01083_),
    .C(_01084_),
    .X(_01154_));
 sky130_fd_sc_hd__nand2_1 _08235_ (.A(_01085_),
    .B(_01154_),
    .Y(_01155_));
 sky130_fd_sc_hd__and3_1 _08236_ (.A(_01090_),
    .B(_01153_),
    .C(_01155_),
    .X(_01156_));
 sky130_fd_sc_hd__a21o_1 _08237_ (.A1(_01090_),
    .A2(_01153_),
    .B1(_01155_),
    .X(_01157_));
 sky130_fd_sc_hd__nand2b_2 _08238_ (.A_N(_01156_),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__xnor2_2 _08239_ (.A(_01079_),
    .B(_01080_),
    .Y(_01159_));
 sky130_fd_sc_hd__xor2_2 _08240_ (.A(_01148_),
    .B(_01149_),
    .X(_01160_));
 sky130_fd_sc_hd__nor2_1 _08241_ (.A(_01159_),
    .B(_01160_),
    .Y(_01161_));
 sky130_fd_sc_hd__xor2_2 _08242_ (.A(_01159_),
    .B(_01160_),
    .X(_01162_));
 sky130_fd_sc_hd__xnor2_2 _08243_ (.A(_01139_),
    .B(_01140_),
    .Y(_01163_));
 sky130_fd_sc_hd__o22a_1 _08244_ (.A1(net149),
    .A2(net24),
    .B1(net22),
    .B2(net125),
    .X(_01164_));
 sky130_fd_sc_hd__xnor2_1 _08245_ (.A(_00359_),
    .B(_01164_),
    .Y(_01165_));
 sky130_fd_sc_hd__nor2_1 _08246_ (.A(net209),
    .B(net19),
    .Y(_01166_));
 sky130_fd_sc_hd__xnor2_1 _08247_ (.A(net96),
    .B(_01166_),
    .Y(_01167_));
 sky130_fd_sc_hd__nor2_1 _08248_ (.A(_01165_),
    .B(_01167_),
    .Y(_01168_));
 sky130_fd_sc_hd__o22a_1 _08249_ (.A1(_00320_),
    .A2(net28),
    .B1(net26),
    .B2(net151),
    .X(_01169_));
 sky130_fd_sc_hd__xnor2_1 _08250_ (.A(net88),
    .B(_01169_),
    .Y(_01170_));
 sky130_fd_sc_hd__and2_1 _08251_ (.A(_01165_),
    .B(_01167_),
    .X(_01171_));
 sky130_fd_sc_hd__nor2_1 _08252_ (.A(_01168_),
    .B(_01171_),
    .Y(_01172_));
 sky130_fd_sc_hd__a21o_1 _08253_ (.A1(_01170_),
    .A2(_01172_),
    .B1(_01168_),
    .X(_01173_));
 sky130_fd_sc_hd__a21o_1 _08254_ (.A1(_01121_),
    .A2(_01124_),
    .B1(_01123_),
    .X(_01174_));
 sky130_fd_sc_hd__or2_1 _08255_ (.A(_01111_),
    .B(_01113_),
    .X(_01175_));
 sky130_fd_sc_hd__and2_1 _08256_ (.A(_01114_),
    .B(_01175_),
    .X(_01176_));
 sky130_fd_sc_hd__and3_1 _08257_ (.A(_01125_),
    .B(_01174_),
    .C(_01176_),
    .X(_01177_));
 sky130_fd_sc_hd__xor2_2 _08258_ (.A(_01133_),
    .B(_01134_),
    .X(_01178_));
 sky130_fd_sc_hd__a21oi_2 _08259_ (.A1(_01125_),
    .A2(_01174_),
    .B1(_01176_),
    .Y(_01179_));
 sky130_fd_sc_hd__or3_1 _08260_ (.A(_01177_),
    .B(_01178_),
    .C(_01179_),
    .X(_01180_));
 sky130_fd_sc_hd__o21bai_2 _08261_ (.A1(_01178_),
    .A2(_01179_),
    .B1_N(_01177_),
    .Y(_01181_));
 sky130_fd_sc_hd__and2_1 _08262_ (.A(_01173_),
    .B(_01181_),
    .X(_01182_));
 sky130_fd_sc_hd__a22o_1 _08263_ (.A1(net128),
    .A2(net121),
    .B1(net114),
    .B2(net126),
    .X(_01183_));
 sky130_fd_sc_hd__xor2_1 _08264_ (.A(net156),
    .B(_01183_),
    .X(_01184_));
 sky130_fd_sc_hd__o22a_1 _08265_ (.A1(net104),
    .A2(net85),
    .B1(net82),
    .B2(net130),
    .X(_01185_));
 sky130_fd_sc_hd__xnor2_1 _08266_ (.A(net175),
    .B(_01185_),
    .Y(_01186_));
 sky130_fd_sc_hd__and2_1 _08267_ (.A(_01184_),
    .B(_01186_),
    .X(_01187_));
 sky130_fd_sc_hd__o22a_1 _08268_ (.A1(net133),
    .A2(net76),
    .B1(net74),
    .B2(net158),
    .X(_01188_));
 sky130_fd_sc_hd__xnor2_1 _08269_ (.A(net181),
    .B(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__a21o_1 _08270_ (.A1(_00200_),
    .A2(_00201_),
    .B1(net286),
    .X(_01190_));
 sky130_fd_sc_hd__nand2_1 _08271_ (.A(_00138_),
    .B(_00229_),
    .Y(_01191_));
 sky130_fd_sc_hd__and3_1 _08272_ (.A(net197),
    .B(_01190_),
    .C(_01191_),
    .X(_01192_));
 sky130_fd_sc_hd__a21oi_1 _08273_ (.A1(_01190_),
    .A2(_01191_),
    .B1(net197),
    .Y(_01193_));
 sky130_fd_sc_hd__or3_2 _08274_ (.A(_01189_),
    .B(_01192_),
    .C(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__a22o_1 _08275_ (.A1(_00159_),
    .A2(_00220_),
    .B1(net71),
    .B2(_00158_),
    .X(_01195_));
 sky130_fd_sc_hd__xnor2_1 _08276_ (.A(net201),
    .B(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__o21ai_1 _08277_ (.A1(_01192_),
    .A2(_01193_),
    .B1(_01189_),
    .Y(_01197_));
 sky130_fd_sc_hd__nand3_2 _08278_ (.A(_01194_),
    .B(_01196_),
    .C(_01197_),
    .Y(_01198_));
 sky130_fd_sc_hd__xnor2_1 _08279_ (.A(net96),
    .B(_01187_),
    .Y(_01199_));
 sky130_fd_sc_hd__a21oi_1 _08280_ (.A1(_01194_),
    .A2(_01198_),
    .B1(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__a21o_1 _08281_ (.A1(net96),
    .A2(_01187_),
    .B1(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__xor2_2 _08282_ (.A(_01173_),
    .B(_01181_),
    .X(_01202_));
 sky130_fd_sc_hd__a21o_1 _08283_ (.A1(_01201_),
    .A2(_01202_),
    .B1(_01182_),
    .X(_01203_));
 sky130_fd_sc_hd__and2b_1 _08284_ (.A_N(_01163_),
    .B(_01203_),
    .X(_01204_));
 sky130_fd_sc_hd__o21ai_1 _08285_ (.A1(_01094_),
    .A2(_01095_),
    .B1(_01097_),
    .Y(_01205_));
 sky130_fd_sc_hd__and2_1 _08286_ (.A(_01105_),
    .B(_01106_),
    .X(_01206_));
 sky130_fd_sc_hd__nor2_1 _08287_ (.A(_01107_),
    .B(_01206_),
    .Y(_01207_));
 sky130_fd_sc_hd__and3_1 _08288_ (.A(_01098_),
    .B(_01205_),
    .C(_01207_),
    .X(_01208_));
 sky130_fd_sc_hd__a21oi_1 _08289_ (.A1(_01098_),
    .A2(_01205_),
    .B1(_01207_),
    .Y(_01209_));
 sky130_fd_sc_hd__and3_1 _08290_ (.A(_01131_),
    .B(_01136_),
    .C(_01137_),
    .X(_01210_));
 sky130_fd_sc_hd__or2_1 _08291_ (.A(_01138_),
    .B(_01210_),
    .X(_01211_));
 sky130_fd_sc_hd__nor3_1 _08292_ (.A(_01208_),
    .B(_01209_),
    .C(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__or2_1 _08293_ (.A(_01208_),
    .B(_01212_),
    .X(_01213_));
 sky130_fd_sc_hd__xnor2_2 _08294_ (.A(_01163_),
    .B(_01203_),
    .Y(_01214_));
 sky130_fd_sc_hd__a21o_1 _08295_ (.A1(_01213_),
    .A2(_01214_),
    .B1(_01204_),
    .X(_01215_));
 sky130_fd_sc_hd__a21oi_1 _08296_ (.A1(_01162_),
    .A2(_01215_),
    .B1(_01161_),
    .Y(_01216_));
 sky130_fd_sc_hd__xnor2_1 _08297_ (.A(_01151_),
    .B(_01152_),
    .Y(_01217_));
 sky130_fd_sc_hd__and2_1 _08298_ (.A(_01216_),
    .B(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__or2_1 _08299_ (.A(_01216_),
    .B(_01217_),
    .X(_01219_));
 sky130_fd_sc_hd__nand2_1 _08300_ (.A(_01145_),
    .B(_01146_),
    .Y(_01220_));
 sky130_fd_sc_hd__nand2_2 _08301_ (.A(_01147_),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__xnor2_2 _08302_ (.A(_01213_),
    .B(_01214_),
    .Y(_01222_));
 sky130_fd_sc_hd__nor2_1 _08303_ (.A(_01221_),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__o22a_1 _08304_ (.A1(net104),
    .A2(net115),
    .B1(net85),
    .B2(net130),
    .X(_01224_));
 sky130_fd_sc_hd__xnor2_2 _08305_ (.A(net175),
    .B(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__a22o_1 _08306_ (.A1(net128),
    .A2(_00372_),
    .B1(net121),
    .B2(net126),
    .X(_01226_));
 sky130_fd_sc_hd__xor2_2 _08307_ (.A(net156),
    .B(_01226_),
    .X(_01227_));
 sky130_fd_sc_hd__nand2_1 _08308_ (.A(_01225_),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__xnor2_1 _08309_ (.A(_01184_),
    .B(_01186_),
    .Y(_01229_));
 sky130_fd_sc_hd__nor2_1 _08310_ (.A(_01228_),
    .B(_01229_),
    .Y(_01230_));
 sky130_fd_sc_hd__xor2_1 _08311_ (.A(_01228_),
    .B(_01229_),
    .X(_01231_));
 sky130_fd_sc_hd__a21o_1 _08312_ (.A1(_01194_),
    .A2(_01197_),
    .B1(_01196_),
    .X(_01232_));
 sky130_fd_sc_hd__and3_1 _08313_ (.A(_01198_),
    .B(_01231_),
    .C(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__a31o_2 _08314_ (.A1(_01198_),
    .A2(_01231_),
    .A3(_01232_),
    .B1(_01230_),
    .X(_01234_));
 sky130_fd_sc_hd__o22a_1 _08315_ (.A1(net125),
    .A2(net84),
    .B1(net80),
    .B2(net124),
    .X(_01235_));
 sky130_fd_sc_hd__xnor2_1 _08316_ (.A(net116),
    .B(_01235_),
    .Y(_01236_));
 sky130_fd_sc_hd__o22a_1 _08317_ (.A1(net110),
    .A2(net69),
    .B1(net67),
    .B2(net123),
    .X(_01237_));
 sky130_fd_sc_hd__xnor2_1 _08318_ (.A(net147),
    .B(_01237_),
    .Y(_01238_));
 sky130_fd_sc_hd__a22o_1 _08319_ (.A1(_00412_),
    .A2(_00465_),
    .B1(_00476_),
    .B2(_00461_),
    .X(_01239_));
 sky130_fd_sc_hd__xnor2_1 _08320_ (.A(_00431_),
    .B(_01239_),
    .Y(_01240_));
 sky130_fd_sc_hd__inv_2 _08321_ (.A(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__xnor2_1 _08322_ (.A(_01236_),
    .B(_01238_),
    .Y(_01242_));
 sky130_fd_sc_hd__nor2_1 _08323_ (.A(_01241_),
    .B(_01242_),
    .Y(_01243_));
 sky130_fd_sc_hd__a21o_2 _08324_ (.A1(_01236_),
    .A2(_01238_),
    .B1(_01243_),
    .X(_01244_));
 sky130_fd_sc_hd__nand2_1 _08325_ (.A(_01234_),
    .B(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__o22a_1 _08326_ (.A1(net133),
    .A2(net82),
    .B1(net76),
    .B2(net158),
    .X(_01246_));
 sky130_fd_sc_hd__xnor2_2 _08327_ (.A(net180),
    .B(_01246_),
    .Y(_01247_));
 sky130_fd_sc_hd__o22a_1 _08328_ (.A1(_00139_),
    .A2(net103),
    .B1(net100),
    .B2(net286),
    .X(_01248_));
 sky130_fd_sc_hd__xnor2_2 _08329_ (.A(net199),
    .B(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__nand2_1 _08330_ (.A(_01247_),
    .B(_01249_),
    .Y(_01250_));
 sky130_fd_sc_hd__a22o_1 _08331_ (.A1(_00158_),
    .A2(_00464_),
    .B1(net71),
    .B2(_00159_),
    .X(_01251_));
 sky130_fd_sc_hd__xnor2_2 _08332_ (.A(net200),
    .B(_01251_),
    .Y(_01252_));
 sky130_fd_sc_hd__xnor2_2 _08333_ (.A(_01247_),
    .B(_01249_),
    .Y(_01253_));
 sky130_fd_sc_hd__o21ai_1 _08334_ (.A1(_01252_),
    .A2(_01253_),
    .B1(_01250_),
    .Y(_01254_));
 sky130_fd_sc_hd__o22a_1 _08335_ (.A1(net151),
    .A2(net24),
    .B1(net22),
    .B2(net149),
    .X(_01255_));
 sky130_fd_sc_hd__xnor2_1 _08336_ (.A(net86),
    .B(_01255_),
    .Y(_01256_));
 sky130_fd_sc_hd__and2_1 _08337_ (.A(_01254_),
    .B(_01256_),
    .X(_01257_));
 sky130_fd_sc_hd__o22a_2 _08338_ (.A1(net209),
    .A2(net28),
    .B1(net26),
    .B2(net152),
    .X(_01258_));
 sky130_fd_sc_hd__xnor2_4 _08339_ (.A(net88),
    .B(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__or2_2 _08340_ (.A(_01254_),
    .B(_01256_),
    .X(_01260_));
 sky130_fd_sc_hd__nand2b_2 _08341_ (.A_N(_01257_),
    .B(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__a21oi_4 _08342_ (.A1(_01259_),
    .A2(_01260_),
    .B1(_01257_),
    .Y(_01262_));
 sky130_fd_sc_hd__xnor2_4 _08343_ (.A(_01234_),
    .B(_01244_),
    .Y(_01263_));
 sky130_fd_sc_hd__o21a_1 _08344_ (.A1(_01262_),
    .A2(_01263_),
    .B1(_01245_),
    .X(_01264_));
 sky130_fd_sc_hd__xor2_2 _08345_ (.A(_01201_),
    .B(_01202_),
    .X(_01265_));
 sky130_fd_sc_hd__and2b_1 _08346_ (.A_N(_01264_),
    .B(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__xor2_1 _08347_ (.A(_01170_),
    .B(_01172_),
    .X(_01267_));
 sky130_fd_sc_hd__o21ai_1 _08348_ (.A1(_01177_),
    .A2(_01179_),
    .B1(_01178_),
    .Y(_01268_));
 sky130_fd_sc_hd__and3_1 _08349_ (.A(_01180_),
    .B(_01267_),
    .C(_01268_),
    .X(_01269_));
 sky130_fd_sc_hd__and3_1 _08350_ (.A(_01194_),
    .B(_01198_),
    .C(_01199_),
    .X(_01270_));
 sky130_fd_sc_hd__or2_1 _08351_ (.A(_01200_),
    .B(_01270_),
    .X(_01271_));
 sky130_fd_sc_hd__a21oi_1 _08352_ (.A1(_01180_),
    .A2(_01268_),
    .B1(_01267_),
    .Y(_01272_));
 sky130_fd_sc_hd__or3_1 _08353_ (.A(_01269_),
    .B(_01271_),
    .C(_01272_),
    .X(_01273_));
 sky130_fd_sc_hd__and2b_1 _08354_ (.A_N(_01269_),
    .B(_01273_),
    .X(_01274_));
 sky130_fd_sc_hd__xnor2_2 _08355_ (.A(_01264_),
    .B(_01265_),
    .Y(_01275_));
 sky130_fd_sc_hd__and2b_1 _08356_ (.A_N(_01274_),
    .B(_01275_),
    .X(_01276_));
 sky130_fd_sc_hd__or2_1 _08357_ (.A(_01266_),
    .B(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__xor2_2 _08358_ (.A(_01221_),
    .B(_01222_),
    .X(_01278_));
 sky130_fd_sc_hd__a21o_1 _08359_ (.A1(_01277_),
    .A2(_01278_),
    .B1(_01223_),
    .X(_01279_));
 sky130_fd_sc_hd__xor2_2 _08360_ (.A(_01162_),
    .B(_01215_),
    .X(_01280_));
 sky130_fd_sc_hd__nand2_1 _08361_ (.A(_01279_),
    .B(_01280_),
    .Y(_01281_));
 sky130_fd_sc_hd__a21o_1 _08362_ (.A1(_01219_),
    .A2(_01281_),
    .B1(_01218_),
    .X(_01282_));
 sky130_fd_sc_hd__nor2_1 _08363_ (.A(_01279_),
    .B(_01280_),
    .Y(_01283_));
 sky130_fd_sc_hd__xnor2_1 _08364_ (.A(_01279_),
    .B(_01280_),
    .Y(_01284_));
 sky130_fd_sc_hd__nand2b_2 _08365_ (.A_N(_01218_),
    .B(_01219_),
    .Y(_01285_));
 sky130_fd_sc_hd__o21a_1 _08366_ (.A1(_01208_),
    .A2(_01209_),
    .B1(_01211_),
    .X(_01286_));
 sky130_fd_sc_hd__nor2_2 _08367_ (.A(_01212_),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__xnor2_2 _08368_ (.A(_01274_),
    .B(_01275_),
    .Y(_01288_));
 sky130_fd_sc_hd__and2_1 _08369_ (.A(_01287_),
    .B(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__xor2_4 _08370_ (.A(_01287_),
    .B(_01288_),
    .X(_01290_));
 sky130_fd_sc_hd__xor2_4 _08371_ (.A(_01262_),
    .B(_01263_),
    .X(_01291_));
 sky130_fd_sc_hd__o22a_1 _08372_ (.A1(net132),
    .A2(net76),
    .B1(net74),
    .B2(net157),
    .X(_01292_));
 sky130_fd_sc_hd__xnor2_1 _08373_ (.A(net201),
    .B(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__a22o_1 _08374_ (.A1(net291),
    .A2(_00220_),
    .B1(net71),
    .B2(_00138_),
    .X(_01294_));
 sky130_fd_sc_hd__xnor2_1 _08375_ (.A(net197),
    .B(_01294_),
    .Y(_01295_));
 sky130_fd_sc_hd__nand2b_1 _08376_ (.A_N(_01293_),
    .B(_01295_),
    .Y(_01296_));
 sky130_fd_sc_hd__xnor2_2 _08377_ (.A(_01225_),
    .B(_01227_),
    .Y(_01297_));
 sky130_fd_sc_hd__nor2_1 _08378_ (.A(_01296_),
    .B(_01297_),
    .Y(_01298_));
 sky130_fd_sc_hd__xor2_2 _08379_ (.A(_01296_),
    .B(_01297_),
    .X(_01299_));
 sky130_fd_sc_hd__xor2_2 _08380_ (.A(_01252_),
    .B(_01253_),
    .X(_01300_));
 sky130_fd_sc_hd__a21o_2 _08381_ (.A1(_01299_),
    .A2(_01300_),
    .B1(_01298_),
    .X(_01301_));
 sky130_fd_sc_hd__o22a_1 _08382_ (.A1(net149),
    .A2(net84),
    .B1(net80),
    .B2(net125),
    .X(_01302_));
 sky130_fd_sc_hd__xnor2_1 _08383_ (.A(_00381_),
    .B(_01302_),
    .Y(_01303_));
 sky130_fd_sc_hd__o22a_1 _08384_ (.A1(net113),
    .A2(net69),
    .B1(net67),
    .B2(net110),
    .X(_01304_));
 sky130_fd_sc_hd__xor2_1 _08385_ (.A(net147),
    .B(_01304_),
    .X(_01305_));
 sky130_fd_sc_hd__nor2_1 _08386_ (.A(_01303_),
    .B(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__a22o_1 _08387_ (.A1(_00287_),
    .A2(_00461_),
    .B1(_00465_),
    .B2(_00476_),
    .X(_01307_));
 sky130_fd_sc_hd__xnor2_1 _08388_ (.A(net109),
    .B(_01307_),
    .Y(_01308_));
 sky130_fd_sc_hd__xnor2_1 _08389_ (.A(_01303_),
    .B(_01305_),
    .Y(_01309_));
 sky130_fd_sc_hd__nor2_1 _08390_ (.A(_01308_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__nor2_2 _08391_ (.A(_01306_),
    .B(_01310_),
    .Y(_01311_));
 sky130_fd_sc_hd__o21a_1 _08392_ (.A1(_01306_),
    .A2(_01310_),
    .B1(_01301_),
    .X(_01312_));
 sky130_fd_sc_hd__o22a_1 _08393_ (.A1(net152),
    .A2(net24),
    .B1(net22),
    .B2(net151),
    .X(_01313_));
 sky130_fd_sc_hd__xnor2_1 _08394_ (.A(net86),
    .B(_01313_),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_1 _08395_ (.A(net209),
    .B(net26),
    .Y(_01315_));
 sky130_fd_sc_hd__mux2_4 _08396_ (.A0(net88),
    .A1(_01314_),
    .S(_01315_),
    .X(_01316_));
 sky130_fd_sc_hd__xnor2_4 _08397_ (.A(_01301_),
    .B(_01311_),
    .Y(_01317_));
 sky130_fd_sc_hd__a21oi_4 _08398_ (.A1(_01316_),
    .A2(_01317_),
    .B1(_01312_),
    .Y(_01318_));
 sky130_fd_sc_hd__and2b_1 _08399_ (.A_N(_01318_),
    .B(_01291_),
    .X(_01319_));
 sky130_fd_sc_hd__a21oi_1 _08400_ (.A1(_01198_),
    .A2(_01232_),
    .B1(_01231_),
    .Y(_01320_));
 sky130_fd_sc_hd__and2_1 _08401_ (.A(_01241_),
    .B(_01242_),
    .X(_01321_));
 sky130_fd_sc_hd__or2_1 _08402_ (.A(_01243_),
    .B(_01321_),
    .X(_01322_));
 sky130_fd_sc_hd__or3_1 _08403_ (.A(_01233_),
    .B(_01320_),
    .C(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__o21ai_1 _08404_ (.A1(_01233_),
    .A2(_01320_),
    .B1(_01322_),
    .Y(_01324_));
 sky130_fd_sc_hd__nand2_2 _08405_ (.A(_01323_),
    .B(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__xnor2_4 _08406_ (.A(_01259_),
    .B(_01261_),
    .Y(_01326_));
 sky130_fd_sc_hd__a21bo_2 _08407_ (.A1(_01324_),
    .A2(_01326_),
    .B1_N(_01323_),
    .X(_01327_));
 sky130_fd_sc_hd__xnor2_4 _08408_ (.A(_01291_),
    .B(_01318_),
    .Y(_01328_));
 sky130_fd_sc_hd__a21o_2 _08409_ (.A1(_01327_),
    .A2(_01328_),
    .B1(_01319_),
    .X(_01329_));
 sky130_fd_sc_hd__a21oi_2 _08410_ (.A1(_01290_),
    .A2(_01329_),
    .B1(_01289_),
    .Y(_01330_));
 sky130_fd_sc_hd__xnor2_2 _08411_ (.A(_01277_),
    .B(_01278_),
    .Y(_01331_));
 sky130_fd_sc_hd__and2_1 _08412_ (.A(_01330_),
    .B(_01331_),
    .X(_01332_));
 sky130_fd_sc_hd__or2_1 _08413_ (.A(_01330_),
    .B(_01331_),
    .X(_01333_));
 sky130_fd_sc_hd__o21ai_1 _08414_ (.A1(_01269_),
    .A2(_01272_),
    .B1(_01271_),
    .Y(_01334_));
 sky130_fd_sc_hd__nand2_2 _08415_ (.A(_01273_),
    .B(_01334_),
    .Y(_01335_));
 sky130_fd_sc_hd__xnor2_4 _08416_ (.A(_01327_),
    .B(_01328_),
    .Y(_01336_));
 sky130_fd_sc_hd__xor2_4 _08417_ (.A(_01316_),
    .B(_01317_),
    .X(_01337_));
 sky130_fd_sc_hd__xnor2_1 _08418_ (.A(_01293_),
    .B(_01295_),
    .Y(_01338_));
 sky130_fd_sc_hd__o22a_1 _08419_ (.A1(net209),
    .A2(net24),
    .B1(net22),
    .B2(net152),
    .X(_01339_));
 sky130_fd_sc_hd__xnor2_1 _08420_ (.A(net86),
    .B(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__nand2_1 _08421_ (.A(_01338_),
    .B(_01340_),
    .Y(_01341_));
 sky130_fd_sc_hd__o22a_1 _08422_ (.A1(net132),
    .A2(net82),
    .B1(net76),
    .B2(net157),
    .X(_01342_));
 sky130_fd_sc_hd__xnor2_1 _08423_ (.A(net201),
    .B(_01342_),
    .Y(_01343_));
 sky130_fd_sc_hd__a22o_1 _08424_ (.A1(_00138_),
    .A2(_00464_),
    .B1(net71),
    .B2(net291),
    .X(_01344_));
 sky130_fd_sc_hd__xnor2_1 _08425_ (.A(net197),
    .B(_01344_),
    .Y(_01345_));
 sky130_fd_sc_hd__nand2b_1 _08426_ (.A_N(_01343_),
    .B(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__xnor2_1 _08427_ (.A(_01338_),
    .B(_01340_),
    .Y(_01347_));
 sky130_fd_sc_hd__o21ai_2 _08428_ (.A1(_01346_),
    .A2(_01347_),
    .B1(_01341_),
    .Y(_01348_));
 sky130_fd_sc_hd__a22o_1 _08429_ (.A1(net126),
    .A2(_00372_),
    .B1(net111),
    .B2(net128),
    .X(_01349_));
 sky130_fd_sc_hd__xor2_1 _08430_ (.A(net156),
    .B(_01349_),
    .X(_01350_));
 sky130_fd_sc_hd__o22a_1 _08431_ (.A1(net133),
    .A2(net85),
    .B1(net82),
    .B2(net158),
    .X(_01351_));
 sky130_fd_sc_hd__xnor2_1 _08432_ (.A(net180),
    .B(_01351_),
    .Y(_01352_));
 sky130_fd_sc_hd__and2_1 _08433_ (.A(_01350_),
    .B(_01352_),
    .X(_01353_));
 sky130_fd_sc_hd__o22a_1 _08434_ (.A1(net104),
    .A2(net119),
    .B1(net115),
    .B2(net130),
    .X(_01354_));
 sky130_fd_sc_hd__xnor2_1 _08435_ (.A(net175),
    .B(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__xor2_1 _08436_ (.A(_01350_),
    .B(_01352_),
    .X(_01356_));
 sky130_fd_sc_hd__and2_1 _08437_ (.A(_01355_),
    .B(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__nor2_1 _08438_ (.A(_01353_),
    .B(_01357_),
    .Y(_01358_));
 sky130_fd_sc_hd__o21a_1 _08439_ (.A1(_01353_),
    .A2(_01357_),
    .B1(_01348_),
    .X(_01359_));
 sky130_fd_sc_hd__o22a_1 _08440_ (.A1(net106),
    .A2(net69),
    .B1(net67),
    .B2(net113),
    .X(_01360_));
 sky130_fd_sc_hd__xnor2_1 _08441_ (.A(net147),
    .B(_01360_),
    .Y(_01361_));
 sky130_fd_sc_hd__o22a_1 _08442_ (.A1(net151),
    .A2(net84),
    .B1(net80),
    .B2(net149),
    .X(_01362_));
 sky130_fd_sc_hd__xnor2_1 _08443_ (.A(net116),
    .B(_01362_),
    .Y(_01363_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(_01361_),
    .B(_01363_),
    .Y(_01364_));
 sky130_fd_sc_hd__o22a_1 _08445_ (.A1(net125),
    .A2(net75),
    .B1(net72),
    .B2(net124),
    .X(_01365_));
 sky130_fd_sc_hd__xnor2_1 _08446_ (.A(net109),
    .B(_01365_),
    .Y(_01366_));
 sky130_fd_sc_hd__inv_2 _08447_ (.A(_01366_),
    .Y(_01367_));
 sky130_fd_sc_hd__or2_1 _08448_ (.A(_01361_),
    .B(_01363_),
    .X(_01368_));
 sky130_fd_sc_hd__nand2_1 _08449_ (.A(_01364_),
    .B(_01368_),
    .Y(_01369_));
 sky130_fd_sc_hd__o21ai_2 _08450_ (.A1(_01367_),
    .A2(_01369_),
    .B1(_01364_),
    .Y(_01370_));
 sky130_fd_sc_hd__xnor2_2 _08451_ (.A(_01348_),
    .B(_01358_),
    .Y(_01371_));
 sky130_fd_sc_hd__a21o_2 _08452_ (.A1(_01370_),
    .A2(_01371_),
    .B1(_01359_),
    .X(_01372_));
 sky130_fd_sc_hd__xnor2_2 _08453_ (.A(_01299_),
    .B(_01300_),
    .Y(_01373_));
 sky130_fd_sc_hd__and2_1 _08454_ (.A(_01308_),
    .B(_01309_),
    .X(_01374_));
 sky130_fd_sc_hd__or2_1 _08455_ (.A(_01310_),
    .B(_01374_),
    .X(_01375_));
 sky130_fd_sc_hd__xor2_1 _08456_ (.A(_01373_),
    .B(_01375_),
    .X(_01376_));
 sky130_fd_sc_hd__xnor2_1 _08457_ (.A(_01314_),
    .B(_01315_),
    .Y(_01377_));
 sky130_fd_sc_hd__and2b_1 _08458_ (.A_N(_01377_),
    .B(_01376_),
    .X(_01378_));
 sky130_fd_sc_hd__o21ba_2 _08459_ (.A1(_01373_),
    .A2(_01375_),
    .B1_N(_01378_),
    .X(_01379_));
 sky130_fd_sc_hd__xor2_4 _08460_ (.A(_01337_),
    .B(_01372_),
    .X(_01380_));
 sky130_fd_sc_hd__nand2b_1 _08461_ (.A_N(_01379_),
    .B(_01380_),
    .Y(_01381_));
 sky130_fd_sc_hd__a21bo_1 _08462_ (.A1(_01337_),
    .A2(_01372_),
    .B1_N(_01381_),
    .X(_01382_));
 sky130_fd_sc_hd__xnor2_2 _08463_ (.A(_01335_),
    .B(_01336_),
    .Y(_01383_));
 sky130_fd_sc_hd__nand2b_1 _08464_ (.A_N(_01383_),
    .B(_01382_),
    .Y(_01384_));
 sky130_fd_sc_hd__o21ai_4 _08465_ (.A1(_01335_),
    .A2(_01336_),
    .B1(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__xor2_4 _08466_ (.A(_01290_),
    .B(_01329_),
    .X(_01386_));
 sky130_fd_sc_hd__nand2_1 _08467_ (.A(_01385_),
    .B(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__a21o_1 _08468_ (.A1(_01333_),
    .A2(_01387_),
    .B1(_01332_),
    .X(_01388_));
 sky130_fd_sc_hd__nor2_1 _08469_ (.A(_01385_),
    .B(_01386_),
    .Y(_01389_));
 sky130_fd_sc_hd__xnor2_4 _08470_ (.A(_01385_),
    .B(_01386_),
    .Y(_01390_));
 sky130_fd_sc_hd__xnor2_2 _08471_ (.A(_01330_),
    .B(_01331_),
    .Y(_01391_));
 sky130_fd_sc_hd__xnor2_4 _08472_ (.A(_01325_),
    .B(_01326_),
    .Y(_01392_));
 sky130_fd_sc_hd__xnor2_4 _08473_ (.A(_01379_),
    .B(_01380_),
    .Y(_01393_));
 sky130_fd_sc_hd__and2_1 _08474_ (.A(_01392_),
    .B(_01393_),
    .X(_01394_));
 sky130_fd_sc_hd__xor2_4 _08475_ (.A(_01392_),
    .B(_01393_),
    .X(_01395_));
 sky130_fd_sc_hd__a22o_1 _08476_ (.A1(net128),
    .A2(_00412_),
    .B1(net111),
    .B2(net126),
    .X(_01396_));
 sky130_fd_sc_hd__xor2_1 _08477_ (.A(net156),
    .B(_01396_),
    .X(_01397_));
 sky130_fd_sc_hd__a32o_1 _08478_ (.A1(_06726_),
    .A2(_00395_),
    .A3(_00396_),
    .B1(net114),
    .B2(_06702_),
    .X(_01398_));
 sky130_fd_sc_hd__xnor2_2 _08479_ (.A(net181),
    .B(_01398_),
    .Y(_01399_));
 sky130_fd_sc_hd__xnor2_1 _08480_ (.A(_01397_),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__o22a_1 _08481_ (.A1(net104),
    .A2(net123),
    .B1(net119),
    .B2(net130),
    .X(_01401_));
 sky130_fd_sc_hd__xnor2_1 _08482_ (.A(_00188_),
    .B(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__nor2_1 _08483_ (.A(_01400_),
    .B(_01402_),
    .Y(_01403_));
 sky130_fd_sc_hd__a21o_1 _08484_ (.A1(_01397_),
    .A2(_01399_),
    .B1(_01403_),
    .X(_01404_));
 sky130_fd_sc_hd__xnor2_1 _08485_ (.A(_01343_),
    .B(_01345_),
    .Y(_01405_));
 sky130_fd_sc_hd__nor2_1 _08486_ (.A(net209),
    .B(net22),
    .Y(_01406_));
 sky130_fd_sc_hd__mux2_1 _08487_ (.A0(net86),
    .A1(_01405_),
    .S(_01406_),
    .X(_01407_));
 sky130_fd_sc_hd__o22a_1 _08488_ (.A1(net152),
    .A2(net84),
    .B1(net80),
    .B2(net151),
    .X(_01408_));
 sky130_fd_sc_hd__xnor2_1 _08489_ (.A(net116),
    .B(_01408_),
    .Y(_01409_));
 sky130_fd_sc_hd__o22a_1 _08490_ (.A1(net124),
    .A2(net69),
    .B1(net67),
    .B2(net106),
    .X(_01410_));
 sky130_fd_sc_hd__xnor2_1 _08491_ (.A(net147),
    .B(_01410_),
    .Y(_01411_));
 sky130_fd_sc_hd__o22a_1 _08492_ (.A1(net149),
    .A2(net75),
    .B1(net72),
    .B2(net125),
    .X(_01412_));
 sky130_fd_sc_hd__xnor2_1 _08493_ (.A(net109),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__inv_2 _08494_ (.A(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hd__xnor2_1 _08495_ (.A(_01409_),
    .B(_01411_),
    .Y(_01415_));
 sky130_fd_sc_hd__or2_1 _08496_ (.A(_01414_),
    .B(_01415_),
    .X(_01416_));
 sky130_fd_sc_hd__a21bo_1 _08497_ (.A1(_01409_),
    .A2(_01411_),
    .B1_N(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__xnor2_1 _08498_ (.A(_01404_),
    .B(_01407_),
    .Y(_01418_));
 sky130_fd_sc_hd__nand2b_1 _08499_ (.A_N(_01418_),
    .B(_01417_),
    .Y(_01419_));
 sky130_fd_sc_hd__a21bo_1 _08500_ (.A1(_01404_),
    .A2(_01407_),
    .B1_N(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__xnor2_2 _08501_ (.A(_01370_),
    .B(_01371_),
    .Y(_01421_));
 sky130_fd_sc_hd__nand2b_1 _08502_ (.A_N(_01421_),
    .B(_01420_),
    .Y(_01422_));
 sky130_fd_sc_hd__xnor2_1 _08503_ (.A(_01346_),
    .B(_01347_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_1 _08504_ (.A(_01355_),
    .B(_01356_),
    .Y(_01424_));
 sky130_fd_sc_hd__or2_1 _08505_ (.A(_01357_),
    .B(_01424_),
    .X(_01425_));
 sky130_fd_sc_hd__xnor2_1 _08506_ (.A(_01367_),
    .B(_01369_),
    .Y(_01426_));
 sky130_fd_sc_hd__xnor2_1 _08507_ (.A(_01423_),
    .B(_01425_),
    .Y(_01427_));
 sky130_fd_sc_hd__nor2_1 _08508_ (.A(_01426_),
    .B(_01427_),
    .Y(_01428_));
 sky130_fd_sc_hd__o21ba_1 _08509_ (.A1(_01423_),
    .A2(_01425_),
    .B1_N(_01428_),
    .X(_01429_));
 sky130_fd_sc_hd__xnor2_2 _08510_ (.A(_01420_),
    .B(_01421_),
    .Y(_01430_));
 sky130_fd_sc_hd__nand2b_1 _08511_ (.A_N(_01429_),
    .B(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__nand2_2 _08512_ (.A(_01422_),
    .B(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__a21oi_2 _08513_ (.A1(_01395_),
    .A2(_01432_),
    .B1(_01394_),
    .Y(_01433_));
 sky130_fd_sc_hd__xor2_2 _08514_ (.A(_01382_),
    .B(_01383_),
    .X(_01434_));
 sky130_fd_sc_hd__and2_1 _08515_ (.A(_01433_),
    .B(_01434_),
    .X(_01435_));
 sky130_fd_sc_hd__and2b_1 _08516_ (.A_N(_01376_),
    .B(_01377_),
    .X(_01436_));
 sky130_fd_sc_hd__nor2_1 _08517_ (.A(_01378_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__xnor2_2 _08518_ (.A(_01429_),
    .B(_01430_),
    .Y(_01438_));
 sky130_fd_sc_hd__nand2_1 _08519_ (.A(_01437_),
    .B(_01438_),
    .Y(_01439_));
 sky130_fd_sc_hd__xnor2_2 _08520_ (.A(_01437_),
    .B(_01438_),
    .Y(_01440_));
 sky130_fd_sc_hd__xnor2_1 _08521_ (.A(_01417_),
    .B(_01418_),
    .Y(_01441_));
 sky130_fd_sc_hd__a22o_1 _08522_ (.A1(net150),
    .A2(_00461_),
    .B1(_00465_),
    .B2(_00340_),
    .X(_01442_));
 sky130_fd_sc_hd__xnor2_1 _08523_ (.A(_00431_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__o22a_1 _08524_ (.A1(net208),
    .A2(net84),
    .B1(net80),
    .B2(net152),
    .X(_01444_));
 sky130_fd_sc_hd__xnor2_1 _08525_ (.A(net116),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__nand2_1 _08526_ (.A(_01443_),
    .B(_01445_),
    .Y(_01446_));
 sky130_fd_sc_hd__o22a_1 _08527_ (.A1(net133),
    .A2(net119),
    .B1(net115),
    .B2(net158),
    .X(_01447_));
 sky130_fd_sc_hd__xnor2_1 _08528_ (.A(net180),
    .B(_01447_),
    .Y(_01448_));
 sky130_fd_sc_hd__o22a_1 _08529_ (.A1(net236),
    .A2(net76),
    .B1(net74),
    .B2(net285),
    .X(_01449_));
 sky130_fd_sc_hd__xnor2_1 _08530_ (.A(net199),
    .B(_01449_),
    .Y(_01450_));
 sky130_fd_sc_hd__nand2_1 _08531_ (.A(_01448_),
    .B(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__xnor2_1 _08532_ (.A(_01448_),
    .B(_01450_),
    .Y(_01452_));
 sky130_fd_sc_hd__o22a_1 _08533_ (.A1(net132),
    .A2(net85),
    .B1(net82),
    .B2(net157),
    .X(_01453_));
 sky130_fd_sc_hd__xnor2_1 _08534_ (.A(net201),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__o21a_1 _08535_ (.A1(_01452_),
    .A2(_01454_),
    .B1(_01451_),
    .X(_01455_));
 sky130_fd_sc_hd__nor2_1 _08536_ (.A(_01446_),
    .B(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__o22a_1 _08537_ (.A1(net125),
    .A2(net69),
    .B1(net67),
    .B2(net124),
    .X(_01457_));
 sky130_fd_sc_hd__xnor2_1 _08538_ (.A(net147),
    .B(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__o22a_1 _08539_ (.A1(net130),
    .A2(net123),
    .B1(net110),
    .B2(net104),
    .X(_01459_));
 sky130_fd_sc_hd__xnor2_1 _08540_ (.A(net175),
    .B(_01459_),
    .Y(_01460_));
 sky130_fd_sc_hd__nand2_1 _08541_ (.A(_01458_),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__a22o_1 _08542_ (.A1(net126),
    .A2(_00412_),
    .B1(_00476_),
    .B2(net128),
    .X(_01462_));
 sky130_fd_sc_hd__xnor2_1 _08543_ (.A(net156),
    .B(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__or2_1 _08544_ (.A(_01458_),
    .B(_01460_),
    .X(_01464_));
 sky130_fd_sc_hd__nand2_1 _08545_ (.A(_01461_),
    .B(_01464_),
    .Y(_01465_));
 sky130_fd_sc_hd__o21ai_1 _08546_ (.A1(_01463_),
    .A2(_01465_),
    .B1(_01461_),
    .Y(_01466_));
 sky130_fd_sc_hd__nand2_1 _08547_ (.A(_01446_),
    .B(_01455_),
    .Y(_01467_));
 sky130_fd_sc_hd__xnor2_1 _08548_ (.A(_01446_),
    .B(_01455_),
    .Y(_01468_));
 sky130_fd_sc_hd__a21oi_1 _08549_ (.A1(_01466_),
    .A2(_01467_),
    .B1(_01456_),
    .Y(_01469_));
 sky130_fd_sc_hd__nand2b_1 _08550_ (.A_N(_01469_),
    .B(_01441_),
    .Y(_01470_));
 sky130_fd_sc_hd__and2_1 _08551_ (.A(_01400_),
    .B(_01402_),
    .X(_01471_));
 sky130_fd_sc_hd__nor2_1 _08552_ (.A(_01403_),
    .B(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__xnor2_1 _08553_ (.A(_01405_),
    .B(_01406_),
    .Y(_01473_));
 sky130_fd_sc_hd__nand2b_1 _08554_ (.A_N(_01473_),
    .B(_01472_),
    .Y(_01474_));
 sky130_fd_sc_hd__xor2_1 _08555_ (.A(_01472_),
    .B(_01473_),
    .X(_01475_));
 sky130_fd_sc_hd__nand2_1 _08556_ (.A(_01414_),
    .B(_01415_),
    .Y(_01476_));
 sky130_fd_sc_hd__nand2_1 _08557_ (.A(_01416_),
    .B(_01476_),
    .Y(_01477_));
 sky130_fd_sc_hd__or2_1 _08558_ (.A(_01475_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__nand2_1 _08559_ (.A(_01474_),
    .B(_01478_),
    .Y(_01479_));
 sky130_fd_sc_hd__xor2_1 _08560_ (.A(_01441_),
    .B(_01469_),
    .X(_01480_));
 sky130_fd_sc_hd__nand2b_1 _08561_ (.A_N(_01480_),
    .B(_01479_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand2_2 _08562_ (.A(_01470_),
    .B(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__inv_2 _08563_ (.A(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__o21a_2 _08564_ (.A1(_01440_),
    .A2(_01483_),
    .B1(_01439_),
    .X(_01484_));
 sky130_fd_sc_hd__xnor2_4 _08565_ (.A(_01395_),
    .B(_01432_),
    .Y(_01485_));
 sky130_fd_sc_hd__or2_1 _08566_ (.A(_01484_),
    .B(_01485_),
    .X(_01486_));
 sky130_fd_sc_hd__or2_1 _08567_ (.A(_01433_),
    .B(_01434_),
    .X(_01487_));
 sky130_fd_sc_hd__a21oi_1 _08568_ (.A1(_01486_),
    .A2(_01487_),
    .B1(_01435_),
    .Y(_01488_));
 sky130_fd_sc_hd__xnor2_1 _08569_ (.A(_01433_),
    .B(_01434_),
    .Y(_01489_));
 sky130_fd_sc_hd__and2_1 _08570_ (.A(_01484_),
    .B(_01485_),
    .X(_01490_));
 sky130_fd_sc_hd__xnor2_4 _08571_ (.A(_01484_),
    .B(_01485_),
    .Y(_01491_));
 sky130_fd_sc_hd__nor2_1 _08572_ (.A(_01489_),
    .B(_01491_),
    .Y(_01492_));
 sky130_fd_sc_hd__xnor2_2 _08573_ (.A(_01440_),
    .B(_01482_),
    .Y(_01493_));
 sky130_fd_sc_hd__and2_1 _08574_ (.A(_01426_),
    .B(_01427_),
    .X(_01494_));
 sky130_fd_sc_hd__nor2_1 _08575_ (.A(_01428_),
    .B(_01494_),
    .Y(_01495_));
 sky130_fd_sc_hd__xnor2_1 _08576_ (.A(_01479_),
    .B(_01480_),
    .Y(_01496_));
 sky130_fd_sc_hd__xnor2_1 _08577_ (.A(_01466_),
    .B(_01468_),
    .Y(_01497_));
 sky130_fd_sc_hd__a22o_1 _08578_ (.A1(_00319_),
    .A2(_00461_),
    .B1(_00465_),
    .B2(net150),
    .X(_01498_));
 sky130_fd_sc_hd__xnor2_1 _08579_ (.A(_00431_),
    .B(_01498_),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _08580_ (.A(net208),
    .B(net80),
    .Y(_01500_));
 sky130_fd_sc_hd__xnor2_1 _08581_ (.A(net116),
    .B(_01500_),
    .Y(_01501_));
 sky130_fd_sc_hd__and2b_1 _08582_ (.A_N(_01501_),
    .B(_01499_),
    .X(_01502_));
 sky130_fd_sc_hd__o22a_1 _08583_ (.A1(net133),
    .A2(net123),
    .B1(net119),
    .B2(net158),
    .X(_01503_));
 sky130_fd_sc_hd__xnor2_2 _08584_ (.A(net180),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__a22o_1 _08585_ (.A1(_00138_),
    .A2(net81),
    .B1(net78),
    .B2(net291),
    .X(_01505_));
 sky130_fd_sc_hd__xnor2_2 _08586_ (.A(net197),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__nand2_1 _08587_ (.A(_01504_),
    .B(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__xnor2_2 _08588_ (.A(_01504_),
    .B(_01506_),
    .Y(_01508_));
 sky130_fd_sc_hd__a22o_1 _08589_ (.A1(_00158_),
    .A2(net114),
    .B1(_00397_),
    .B2(_00159_),
    .X(_01509_));
 sky130_fd_sc_hd__xnor2_2 _08590_ (.A(net200),
    .B(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__o21ai_2 _08591_ (.A1(_01508_),
    .A2(_01510_),
    .B1(_01507_),
    .Y(_01511_));
 sky130_fd_sc_hd__nand2_1 _08592_ (.A(_01502_),
    .B(_01511_),
    .Y(_01512_));
 sky130_fd_sc_hd__o22a_1 _08593_ (.A1(net149),
    .A2(net69),
    .B1(net67),
    .B2(net125),
    .X(_01513_));
 sky130_fd_sc_hd__xnor2_1 _08594_ (.A(net147),
    .B(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__o22a_1 _08595_ (.A1(net104),
    .A2(net113),
    .B1(net110),
    .B2(net130),
    .X(_01515_));
 sky130_fd_sc_hd__xnor2_1 _08596_ (.A(net175),
    .B(_01515_),
    .Y(_01516_));
 sky130_fd_sc_hd__nand2_1 _08597_ (.A(_01514_),
    .B(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__a22o_1 _08598_ (.A1(net128),
    .A2(_00287_),
    .B1(_00476_),
    .B2(net126),
    .X(_01518_));
 sky130_fd_sc_hd__xnor2_2 _08599_ (.A(net156),
    .B(_01518_),
    .Y(_01519_));
 sky130_fd_sc_hd__xnor2_1 _08600_ (.A(_01514_),
    .B(_01516_),
    .Y(_01520_));
 sky130_fd_sc_hd__o21ai_2 _08601_ (.A1(_01519_),
    .A2(_01520_),
    .B1(_01517_),
    .Y(_01521_));
 sky130_fd_sc_hd__inv_2 _08602_ (.A(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__xnor2_2 _08603_ (.A(_01502_),
    .B(_01511_),
    .Y(_01523_));
 sky130_fd_sc_hd__o21a_1 _08604_ (.A1(_01522_),
    .A2(_01523_),
    .B1(_01512_),
    .X(_01524_));
 sky130_fd_sc_hd__nand2b_1 _08605_ (.A_N(_01524_),
    .B(_01497_),
    .Y(_01525_));
 sky130_fd_sc_hd__xnor2_1 _08606_ (.A(_01452_),
    .B(_01454_),
    .Y(_01526_));
 sky130_fd_sc_hd__or2_1 _08607_ (.A(_01443_),
    .B(_01445_),
    .X(_01527_));
 sky130_fd_sc_hd__nand2_1 _08608_ (.A(_01446_),
    .B(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__xnor2_1 _08609_ (.A(_01526_),
    .B(_01528_),
    .Y(_01529_));
 sky130_fd_sc_hd__xnor2_1 _08610_ (.A(_01463_),
    .B(_01465_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_1 _08611_ (.A(_01529_),
    .B(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__o21bai_1 _08612_ (.A1(_01526_),
    .A2(_01528_),
    .B1_N(_01531_),
    .Y(_01532_));
 sky130_fd_sc_hd__xnor2_1 _08613_ (.A(_01497_),
    .B(_01524_),
    .Y(_01533_));
 sky130_fd_sc_hd__a21bo_1 _08614_ (.A1(_01532_),
    .A2(_01533_),
    .B1_N(_01525_),
    .X(_01534_));
 sky130_fd_sc_hd__xnor2_1 _08615_ (.A(_01495_),
    .B(_01496_),
    .Y(_01535_));
 sky130_fd_sc_hd__nand2b_1 _08616_ (.A_N(_01535_),
    .B(_01534_),
    .Y(_01536_));
 sky130_fd_sc_hd__a21bo_1 _08617_ (.A1(_01495_),
    .A2(_01496_),
    .B1_N(_01536_),
    .X(_01537_));
 sky130_fd_sc_hd__or2_1 _08618_ (.A(_01493_),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__nand2_1 _08619_ (.A(_01493_),
    .B(_01537_),
    .Y(_01539_));
 sky130_fd_sc_hd__nand2_1 _08620_ (.A(_01475_),
    .B(_01477_),
    .Y(_01540_));
 sky130_fd_sc_hd__nand2_1 _08621_ (.A(_01478_),
    .B(_01540_),
    .Y(_01541_));
 sky130_fd_sc_hd__xnor2_1 _08622_ (.A(_01532_),
    .B(_01533_),
    .Y(_01542_));
 sky130_fd_sc_hd__or2_1 _08623_ (.A(_01541_),
    .B(_01542_),
    .X(_01543_));
 sky130_fd_sc_hd__o22a_1 _08624_ (.A1(net130),
    .A2(net113),
    .B1(net106),
    .B2(net104),
    .X(_01544_));
 sky130_fd_sc_hd__xnor2_2 _08625_ (.A(net175),
    .B(_01544_),
    .Y(_01545_));
 sky130_fd_sc_hd__a22o_1 _08626_ (.A1(net128),
    .A2(_00266_),
    .B1(_00287_),
    .B2(net126),
    .X(_01546_));
 sky130_fd_sc_hd__xor2_2 _08627_ (.A(net156),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__nand2_2 _08628_ (.A(_01545_),
    .B(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _08629_ (.A(_00381_),
    .B(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__a22o_1 _08630_ (.A1(_06726_),
    .A2(_00372_),
    .B1(net111),
    .B2(_06702_),
    .X(_01550_));
 sky130_fd_sc_hd__xnor2_2 _08631_ (.A(net181),
    .B(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__a22o_1 _08632_ (.A1(_00138_),
    .A2(_00397_),
    .B1(net81),
    .B2(net291),
    .X(_01552_));
 sky130_fd_sc_hd__xnor2_2 _08633_ (.A(net197),
    .B(_01552_),
    .Y(_01553_));
 sky130_fd_sc_hd__nand2_1 _08634_ (.A(_01551_),
    .B(_01553_),
    .Y(_01554_));
 sky130_fd_sc_hd__o22a_1 _08635_ (.A1(net132),
    .A2(net119),
    .B1(net115),
    .B2(net157),
    .X(_01555_));
 sky130_fd_sc_hd__xnor2_2 _08636_ (.A(net201),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__xnor2_2 _08637_ (.A(_01551_),
    .B(_01553_),
    .Y(_01557_));
 sky130_fd_sc_hd__o21ai_4 _08638_ (.A1(_01556_),
    .A2(_01557_),
    .B1(_01554_),
    .Y(_01558_));
 sky130_fd_sc_hd__nand2_1 _08639_ (.A(_00381_),
    .B(_01548_),
    .Y(_01559_));
 sky130_fd_sc_hd__xnor2_2 _08640_ (.A(_00381_),
    .B(_01548_),
    .Y(_01560_));
 sky130_fd_sc_hd__a21o_1 _08641_ (.A1(_01558_),
    .A2(_01559_),
    .B1(_01549_),
    .X(_01561_));
 sky130_fd_sc_hd__xnor2_2 _08642_ (.A(_01521_),
    .B(_01523_),
    .Y(_01562_));
 sky130_fd_sc_hd__xor2_1 _08643_ (.A(_01508_),
    .B(_01510_),
    .X(_01563_));
 sky130_fd_sc_hd__and2b_1 _08644_ (.A_N(_01499_),
    .B(_01501_),
    .X(_01564_));
 sky130_fd_sc_hd__nor2_1 _08645_ (.A(_01502_),
    .B(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__xnor2_1 _08646_ (.A(_01563_),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__xnor2_1 _08647_ (.A(_01519_),
    .B(_01520_),
    .Y(_01567_));
 sky130_fd_sc_hd__or2_1 _08648_ (.A(_01566_),
    .B(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__a21bo_1 _08649_ (.A1(_01563_),
    .A2(_01565_),
    .B1_N(_01568_),
    .X(_01569_));
 sky130_fd_sc_hd__xnor2_2 _08650_ (.A(_01561_),
    .B(_01562_),
    .Y(_01570_));
 sky130_fd_sc_hd__and2b_1 _08651_ (.A_N(_01570_),
    .B(_01569_),
    .X(_01571_));
 sky130_fd_sc_hd__a21oi_2 _08652_ (.A1(_01561_),
    .A2(_01562_),
    .B1(_01571_),
    .Y(_01572_));
 sky130_fd_sc_hd__xor2_2 _08653_ (.A(_01541_),
    .B(_01542_),
    .X(_01573_));
 sky130_fd_sc_hd__nand2b_1 _08654_ (.A_N(_01572_),
    .B(_01573_),
    .Y(_01574_));
 sky130_fd_sc_hd__xor2_1 _08655_ (.A(_01534_),
    .B(_01535_),
    .X(_01575_));
 sky130_fd_sc_hd__a21oi_2 _08656_ (.A1(_01543_),
    .A2(_01574_),
    .B1(_01575_),
    .Y(_01576_));
 sky130_fd_sc_hd__a21o_1 _08657_ (.A1(_01493_),
    .A2(_01537_),
    .B1(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__and2_1 _08658_ (.A(_01529_),
    .B(_01530_),
    .X(_01578_));
 sky130_fd_sc_hd__nor2_2 _08659_ (.A(_01531_),
    .B(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__xnor2_2 _08660_ (.A(_01569_),
    .B(_01570_),
    .Y(_01580_));
 sky130_fd_sc_hd__and2_1 _08661_ (.A(_01579_),
    .B(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__xnor2_4 _08662_ (.A(_01558_),
    .B(_01560_),
    .Y(_01582_));
 sky130_fd_sc_hd__a22o_1 _08663_ (.A1(_06702_),
    .A2(_00412_),
    .B1(net111),
    .B2(_06726_),
    .X(_01583_));
 sky130_fd_sc_hd__xnor2_2 _08664_ (.A(net181),
    .B(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__a32o_1 _08665_ (.A1(net292),
    .A2(_00395_),
    .A3(_00396_),
    .B1(_00138_),
    .B2(net114),
    .X(_01585_));
 sky130_fd_sc_hd__xnor2_2 _08666_ (.A(net197),
    .B(_01585_),
    .Y(_01586_));
 sky130_fd_sc_hd__nand2_1 _08667_ (.A(_01584_),
    .B(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__o22a_1 _08668_ (.A1(net132),
    .A2(net123),
    .B1(net119),
    .B2(net157),
    .X(_01588_));
 sky130_fd_sc_hd__xnor2_2 _08669_ (.A(net201),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__xnor2_2 _08670_ (.A(_01584_),
    .B(_01586_),
    .Y(_01590_));
 sky130_fd_sc_hd__o21ai_2 _08671_ (.A1(_01589_),
    .A2(_01590_),
    .B1(_01587_),
    .Y(_01591_));
 sky130_fd_sc_hd__o22a_1 _08672_ (.A1(net151),
    .A2(net69),
    .B1(net67),
    .B2(net149),
    .X(_01592_));
 sky130_fd_sc_hd__xnor2_2 _08673_ (.A(net147),
    .B(_01592_),
    .Y(_01593_));
 sky130_fd_sc_hd__and2_1 _08674_ (.A(_01591_),
    .B(_01593_),
    .X(_01594_));
 sky130_fd_sc_hd__o22a_1 _08675_ (.A1(net208),
    .A2(net75),
    .B1(net72),
    .B2(net152),
    .X(_01595_));
 sky130_fd_sc_hd__xnor2_2 _08676_ (.A(net109),
    .B(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__xor2_2 _08677_ (.A(_01591_),
    .B(_01593_),
    .X(_01597_));
 sky130_fd_sc_hd__a21o_1 _08678_ (.A1(_01596_),
    .A2(_01597_),
    .B1(_01594_),
    .X(_01598_));
 sky130_fd_sc_hd__and2_1 _08679_ (.A(_01582_),
    .B(_01598_),
    .X(_01599_));
 sky130_fd_sc_hd__a22o_1 _08680_ (.A1(net126),
    .A2(_00266_),
    .B1(_00340_),
    .B2(net128),
    .X(_01600_));
 sky130_fd_sc_hd__xor2_1 _08681_ (.A(net156),
    .B(_01600_),
    .X(_01601_));
 sky130_fd_sc_hd__o22a_1 _08682_ (.A1(net104),
    .A2(net124),
    .B1(net106),
    .B2(net130),
    .X(_01602_));
 sky130_fd_sc_hd__xnor2_1 _08683_ (.A(net175),
    .B(_01602_),
    .Y(_01603_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_01601_),
    .B(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__xnor2_2 _08685_ (.A(_01545_),
    .B(_01547_),
    .Y(_01605_));
 sky130_fd_sc_hd__xor2_1 _08686_ (.A(_01556_),
    .B(_01557_),
    .X(_01606_));
 sky130_fd_sc_hd__xor2_1 _08687_ (.A(_01604_),
    .B(_01605_),
    .X(_01607_));
 sky130_fd_sc_hd__and2_1 _08688_ (.A(_01606_),
    .B(_01607_),
    .X(_01608_));
 sky130_fd_sc_hd__o21bai_4 _08689_ (.A1(_01604_),
    .A2(_01605_),
    .B1_N(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__xor2_4 _08690_ (.A(_01582_),
    .B(_01598_),
    .X(_01610_));
 sky130_fd_sc_hd__a21o_2 _08691_ (.A1(_01609_),
    .A2(_01610_),
    .B1(_01599_),
    .X(_01611_));
 sky130_fd_sc_hd__xor2_4 _08692_ (.A(_01579_),
    .B(_01580_),
    .X(_01612_));
 sky130_fd_sc_hd__a21o_1 _08693_ (.A1(_01611_),
    .A2(_01612_),
    .B1(_01581_),
    .X(_01613_));
 sky130_fd_sc_hd__xnor2_2 _08694_ (.A(_01572_),
    .B(_01573_),
    .Y(_01614_));
 sky130_fd_sc_hd__or2_1 _08695_ (.A(_01613_),
    .B(_01614_),
    .X(_01615_));
 sky130_fd_sc_hd__nand2_1 _08696_ (.A(_01613_),
    .B(_01614_),
    .Y(_01616_));
 sky130_fd_sc_hd__nand2_1 _08697_ (.A(_01566_),
    .B(_01567_),
    .Y(_01617_));
 sky130_fd_sc_hd__nand2_4 _08698_ (.A(_01568_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__xnor2_4 _08699_ (.A(_01609_),
    .B(_01610_),
    .Y(_01619_));
 sky130_fd_sc_hd__xnor2_4 _08700_ (.A(_01618_),
    .B(_01619_),
    .Y(_01620_));
 sky130_fd_sc_hd__xnor2_2 _08701_ (.A(_01596_),
    .B(_01597_),
    .Y(_01621_));
 sky130_fd_sc_hd__o22a_1 _08702_ (.A1(net152),
    .A2(net69),
    .B1(net67),
    .B2(net151),
    .X(_01622_));
 sky130_fd_sc_hd__xnor2_2 _08703_ (.A(net147),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_1 _08704_ (.A(net208),
    .B(net72),
    .Y(_01624_));
 sky130_fd_sc_hd__mux2_1 _08705_ (.A0(net109),
    .A1(_01623_),
    .S(_01624_),
    .X(_01625_));
 sky130_fd_sc_hd__nand2b_1 _08706_ (.A_N(_01621_),
    .B(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hd__a22o_1 _08707_ (.A1(_00159_),
    .A2(_00372_),
    .B1(net111),
    .B2(_00158_),
    .X(_01627_));
 sky130_fd_sc_hd__xnor2_1 _08708_ (.A(net200),
    .B(_01627_),
    .Y(_01628_));
 sky130_fd_sc_hd__o22a_1 _08709_ (.A1(net236),
    .A2(net119),
    .B1(net115),
    .B2(net285),
    .X(_01629_));
 sky130_fd_sc_hd__xnor2_2 _08710_ (.A(net199),
    .B(_01629_),
    .Y(_01630_));
 sky130_fd_sc_hd__nand2b_1 _08711_ (.A_N(_01628_),
    .B(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__xnor2_1 _08712_ (.A(_01601_),
    .B(_01603_),
    .Y(_01632_));
 sky130_fd_sc_hd__or2_1 _08713_ (.A(_01631_),
    .B(_01632_),
    .X(_01633_));
 sky130_fd_sc_hd__xnor2_1 _08714_ (.A(_01631_),
    .B(_01632_),
    .Y(_01634_));
 sky130_fd_sc_hd__xnor2_2 _08715_ (.A(_01589_),
    .B(_01590_),
    .Y(_01635_));
 sky130_fd_sc_hd__o21a_1 _08716_ (.A1(_01634_),
    .A2(_01635_),
    .B1(_01633_),
    .X(_01636_));
 sky130_fd_sc_hd__xnor2_2 _08717_ (.A(_01621_),
    .B(_01625_),
    .Y(_01637_));
 sky130_fd_sc_hd__nand2b_1 _08718_ (.A_N(_01636_),
    .B(_01637_),
    .Y(_01638_));
 sky130_fd_sc_hd__nand2_2 _08719_ (.A(_01626_),
    .B(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__nand2b_1 _08720_ (.A_N(_01620_),
    .B(_01639_),
    .Y(_01640_));
 sky130_fd_sc_hd__o21ai_4 _08721_ (.A1(_01618_),
    .A2(_01619_),
    .B1(_01640_),
    .Y(_01641_));
 sky130_fd_sc_hd__xor2_4 _08722_ (.A(_01611_),
    .B(_01612_),
    .X(_01642_));
 sky130_fd_sc_hd__a22o_1 _08723_ (.A1(_01613_),
    .A2(_01614_),
    .B1(_01641_),
    .B2(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__xor2_1 _08724_ (.A(_01613_),
    .B(_01614_),
    .X(_01644_));
 sky130_fd_sc_hd__nand2_1 _08725_ (.A(_01615_),
    .B(_01616_),
    .Y(_01645_));
 sky130_fd_sc_hd__xor2_4 _08726_ (.A(_01641_),
    .B(_01642_),
    .X(_01646_));
 sky130_fd_sc_hd__xor2_4 _08727_ (.A(_01620_),
    .B(_01639_),
    .X(_01647_));
 sky130_fd_sc_hd__nor2_1 _08728_ (.A(_01606_),
    .B(_01607_),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_2 _08729_ (.A(_01608_),
    .B(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__xnor2_2 _08730_ (.A(_01636_),
    .B(_01637_),
    .Y(_01650_));
 sky130_fd_sc_hd__and2_1 _08731_ (.A(_01649_),
    .B(_01650_),
    .X(_01651_));
 sky130_fd_sc_hd__a22o_1 _08732_ (.A1(net128),
    .A2(net150),
    .B1(_00340_),
    .B2(net126),
    .X(_01652_));
 sky130_fd_sc_hd__xor2_2 _08733_ (.A(net156),
    .B(_01652_),
    .X(_01653_));
 sky130_fd_sc_hd__o22a_1 _08734_ (.A1(net158),
    .A2(net113),
    .B1(net106),
    .B2(net133),
    .X(_01654_));
 sky130_fd_sc_hd__xnor2_2 _08735_ (.A(net180),
    .B(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__nand2_1 _08736_ (.A(_01653_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__o22a_1 _08737_ (.A1(net104),
    .A2(net125),
    .B1(net124),
    .B2(net130),
    .X(_01657_));
 sky130_fd_sc_hd__xnor2_2 _08738_ (.A(_00188_),
    .B(_01657_),
    .Y(_01658_));
 sky130_fd_sc_hd__xnor2_2 _08739_ (.A(_01653_),
    .B(_01655_),
    .Y(_01659_));
 sky130_fd_sc_hd__or2_1 _08740_ (.A(_01658_),
    .B(_01659_),
    .X(_01660_));
 sky130_fd_sc_hd__o21ai_1 _08741_ (.A1(_01658_),
    .A2(_01659_),
    .B1(_01656_),
    .Y(_01661_));
 sky130_fd_sc_hd__xnor2_2 _08742_ (.A(_01623_),
    .B(_01624_),
    .Y(_01662_));
 sky130_fd_sc_hd__a21o_1 _08743_ (.A1(_01656_),
    .A2(_01660_),
    .B1(_01662_),
    .X(_01663_));
 sky130_fd_sc_hd__xnor2_1 _08744_ (.A(_01628_),
    .B(_01630_),
    .Y(_01664_));
 sky130_fd_sc_hd__o22a_1 _08745_ (.A1(net208),
    .A2(net69),
    .B1(net67),
    .B2(net152),
    .X(_01665_));
 sky130_fd_sc_hd__xnor2_1 _08746_ (.A(net147),
    .B(_01665_),
    .Y(_01666_));
 sky130_fd_sc_hd__nand2_1 _08747_ (.A(_01664_),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__a22o_1 _08748_ (.A1(_00158_),
    .A2(_00412_),
    .B1(net111),
    .B2(_00159_),
    .X(_01668_));
 sky130_fd_sc_hd__xnor2_2 _08749_ (.A(net200),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__o22a_1 _08750_ (.A1(net236),
    .A2(net123),
    .B1(net119),
    .B2(net285),
    .X(_01670_));
 sky130_fd_sc_hd__xnor2_2 _08751_ (.A(net199),
    .B(_01670_),
    .Y(_01671_));
 sky130_fd_sc_hd__nand2b_1 _08752_ (.A_N(_01669_),
    .B(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__xnor2_1 _08753_ (.A(_01664_),
    .B(_01666_),
    .Y(_01673_));
 sky130_fd_sc_hd__o21a_1 _08754_ (.A1(_01672_),
    .A2(_01673_),
    .B1(_01667_),
    .X(_01674_));
 sky130_fd_sc_hd__and3_1 _08755_ (.A(_01656_),
    .B(_01660_),
    .C(_01662_),
    .X(_01675_));
 sky130_fd_sc_hd__xnor2_1 _08756_ (.A(_01661_),
    .B(_01662_),
    .Y(_01676_));
 sky130_fd_sc_hd__o21ai_4 _08757_ (.A1(_01674_),
    .A2(_01675_),
    .B1(_01663_),
    .Y(_01677_));
 sky130_fd_sc_hd__xor2_4 _08758_ (.A(_01649_),
    .B(_01650_),
    .X(_01678_));
 sky130_fd_sc_hd__a21oi_2 _08759_ (.A1(_01677_),
    .A2(_01678_),
    .B1(_01651_),
    .Y(_01679_));
 sky130_fd_sc_hd__nand2_1 _08760_ (.A(_01647_),
    .B(_01679_),
    .Y(_01680_));
 sky130_fd_sc_hd__xnor2_1 _08761_ (.A(_01634_),
    .B(_01635_),
    .Y(_01681_));
 sky130_fd_sc_hd__xor2_1 _08762_ (.A(_01674_),
    .B(_01676_),
    .X(_01682_));
 sky130_fd_sc_hd__nor2_1 _08763_ (.A(_01681_),
    .B(_01682_),
    .Y(_01683_));
 sky130_fd_sc_hd__xor2_1 _08764_ (.A(_01681_),
    .B(_01682_),
    .X(_01684_));
 sky130_fd_sc_hd__nand2_1 _08765_ (.A(_01658_),
    .B(_01659_),
    .Y(_01685_));
 sky130_fd_sc_hd__xnor2_1 _08766_ (.A(_01658_),
    .B(_01659_),
    .Y(_01686_));
 sky130_fd_sc_hd__a22o_1 _08767_ (.A1(net128),
    .A2(_00319_),
    .B1(net150),
    .B2(net126),
    .X(_01687_));
 sky130_fd_sc_hd__xor2_1 _08768_ (.A(net156),
    .B(_01687_),
    .X(_01688_));
 sky130_fd_sc_hd__o22a_1 _08769_ (.A1(net133),
    .A2(net124),
    .B1(net106),
    .B2(net158),
    .X(_01689_));
 sky130_fd_sc_hd__xnor2_1 _08770_ (.A(net180),
    .B(_01689_),
    .Y(_01690_));
 sky130_fd_sc_hd__and2_1 _08771_ (.A(_01688_),
    .B(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__o22a_1 _08772_ (.A1(net130),
    .A2(net125),
    .B1(net149),
    .B2(net104),
    .X(_01692_));
 sky130_fd_sc_hd__xnor2_1 _08773_ (.A(net175),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__xor2_1 _08774_ (.A(_01688_),
    .B(_01690_),
    .X(_01694_));
 sky130_fd_sc_hd__a21o_1 _08775_ (.A1(_01693_),
    .A2(_01694_),
    .B1(_01691_),
    .X(_01695_));
 sky130_fd_sc_hd__xnor2_1 _08776_ (.A(_01686_),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__xnor2_1 _08777_ (.A(_01669_),
    .B(_01671_),
    .Y(_01697_));
 sky130_fd_sc_hd__or3_1 _08778_ (.A(net208),
    .B(net67),
    .C(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__o21bai_1 _08779_ (.A1(net209),
    .A2(net67),
    .B1_N(net147),
    .Y(_01699_));
 sky130_fd_sc_hd__nand2_1 _08780_ (.A(_01698_),
    .B(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__and3_1 _08781_ (.A(_01696_),
    .B(_01698_),
    .C(_01699_),
    .X(_01701_));
 sky130_fd_sc_hd__a31o_1 _08782_ (.A1(_01660_),
    .A2(_01685_),
    .A3(_01695_),
    .B1(_01701_),
    .X(_01702_));
 sky130_fd_sc_hd__a21o_1 _08783_ (.A1(_01684_),
    .A2(_01702_),
    .B1(_01683_),
    .X(_01703_));
 sky130_fd_sc_hd__xor2_4 _08784_ (.A(_01677_),
    .B(_01678_),
    .X(_01704_));
 sky130_fd_sc_hd__a2bb2o_1 _08785_ (.A1_N(_01647_),
    .A2_N(_01679_),
    .B1(_01703_),
    .B2(_01704_),
    .X(_01705_));
 sky130_fd_sc_hd__xor2_2 _08786_ (.A(_01647_),
    .B(_01679_),
    .X(_01706_));
 sky130_fd_sc_hd__or2_2 _08787_ (.A(_01703_),
    .B(_01704_),
    .X(_01707_));
 sky130_fd_sc_hd__xor2_2 _08788_ (.A(_01703_),
    .B(_01704_),
    .X(_01708_));
 sky130_fd_sc_hd__xnor2_1 _08789_ (.A(_01684_),
    .B(_01702_),
    .Y(_01709_));
 sky130_fd_sc_hd__xor2_1 _08790_ (.A(_01672_),
    .B(_01673_),
    .X(_01710_));
 sky130_fd_sc_hd__xnor2_1 _08791_ (.A(_01696_),
    .B(_01700_),
    .Y(_01711_));
 sky130_fd_sc_hd__nand2_1 _08792_ (.A(_01710_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__xnor2_1 _08793_ (.A(_01710_),
    .B(_01711_),
    .Y(_01713_));
 sky130_fd_sc_hd__o22a_1 _08794_ (.A1(net133),
    .A2(net125),
    .B1(net124),
    .B2(net158),
    .X(_01714_));
 sky130_fd_sc_hd__xnor2_1 _08795_ (.A(net180),
    .B(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__a22o_1 _08796_ (.A1(net291),
    .A2(_00372_),
    .B1(net111),
    .B2(_00138_),
    .X(_01716_));
 sky130_fd_sc_hd__xnor2_1 _08797_ (.A(net197),
    .B(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__nand2_1 _08798_ (.A(_01715_),
    .B(_01717_),
    .Y(_01718_));
 sky130_fd_sc_hd__xnor2_1 _08799_ (.A(_01715_),
    .B(_01717_),
    .Y(_01719_));
 sky130_fd_sc_hd__o22a_1 _08800_ (.A1(net157),
    .A2(net113),
    .B1(net106),
    .B2(net132),
    .X(_01720_));
 sky130_fd_sc_hd__xnor2_2 _08801_ (.A(net200),
    .B(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__inv_2 _08802_ (.A(_01721_),
    .Y(_01722_));
 sky130_fd_sc_hd__o21ai_1 _08803_ (.A1(_01719_),
    .A2(_01722_),
    .B1(_01718_),
    .Y(_01723_));
 sky130_fd_sc_hd__xnor2_1 _08804_ (.A(_01693_),
    .B(_01694_),
    .Y(_01724_));
 sky130_fd_sc_hd__nand2b_1 _08805_ (.A_N(_01724_),
    .B(_01723_),
    .Y(_01725_));
 sky130_fd_sc_hd__a22o_1 _08806_ (.A1(net206),
    .A2(net128),
    .B1(net126),
    .B2(_00319_),
    .X(_01726_));
 sky130_fd_sc_hd__xor2_1 _08807_ (.A(net156),
    .B(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__o22a_1 _08808_ (.A1(net104),
    .A2(net151),
    .B1(net149),
    .B2(net130),
    .X(_01728_));
 sky130_fd_sc_hd__xnor2_1 _08809_ (.A(net175),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__and2_1 _08810_ (.A(_01727_),
    .B(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__xnor2_1 _08811_ (.A(_01723_),
    .B(_01724_),
    .Y(_01731_));
 sky130_fd_sc_hd__a21bo_1 _08812_ (.A1(_01730_),
    .A2(_01731_),
    .B1_N(_01725_),
    .X(_01732_));
 sky130_fd_sc_hd__nand2b_1 _08813_ (.A_N(_01713_),
    .B(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__and3_1 _08814_ (.A(_01709_),
    .B(_01712_),
    .C(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__xnor2_1 _08815_ (.A(_01713_),
    .B(_01732_),
    .Y(_01735_));
 sky130_fd_sc_hd__xnor2_1 _08816_ (.A(_01730_),
    .B(_01731_),
    .Y(_01736_));
 sky130_fd_sc_hd__o21ai_1 _08817_ (.A1(net209),
    .A2(net67),
    .B1(_01697_),
    .Y(_01737_));
 sky130_fd_sc_hd__and2_1 _08818_ (.A(_01698_),
    .B(_01737_),
    .X(_01738_));
 sky130_fd_sc_hd__nor2_1 _08819_ (.A(_01736_),
    .B(_01738_),
    .Y(_01739_));
 sky130_fd_sc_hd__xnor2_1 _08820_ (.A(_01719_),
    .B(_01721_),
    .Y(_01740_));
 sky130_fd_sc_hd__o22a_1 _08821_ (.A1(net158),
    .A2(net125),
    .B1(net149),
    .B2(net133),
    .X(_01741_));
 sky130_fd_sc_hd__xnor2_2 _08822_ (.A(net180),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__a22o_1 _08823_ (.A1(_00138_),
    .A2(_00412_),
    .B1(net111),
    .B2(net291),
    .X(_01743_));
 sky130_fd_sc_hd__xnor2_2 _08824_ (.A(net197),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__nand2_1 _08825_ (.A(_01742_),
    .B(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__o22a_1 _08826_ (.A1(net132),
    .A2(net124),
    .B1(net106),
    .B2(net157),
    .X(_01746_));
 sky130_fd_sc_hd__xnor2_2 _08827_ (.A(net201),
    .B(_01746_),
    .Y(_01747_));
 sky130_fd_sc_hd__xnor2_2 _08828_ (.A(_01742_),
    .B(_01744_),
    .Y(_01748_));
 sky130_fd_sc_hd__o21a_1 _08829_ (.A1(_01747_),
    .A2(_01748_),
    .B1(_01745_),
    .X(_01749_));
 sky130_fd_sc_hd__nand2b_1 _08830_ (.A_N(_01749_),
    .B(_01740_),
    .Y(_01750_));
 sky130_fd_sc_hd__o22a_1 _08831_ (.A1(net104),
    .A2(net152),
    .B1(net151),
    .B2(net130),
    .X(_01751_));
 sky130_fd_sc_hd__xnor2_1 _08832_ (.A(_00188_),
    .B(_01751_),
    .Y(_01752_));
 sky130_fd_sc_hd__nor2_1 _08833_ (.A(net212),
    .B(_00232_),
    .Y(_01753_));
 sky130_fd_sc_hd__xnor2_2 _08834_ (.A(net154),
    .B(_01753_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_1 _08835_ (.A(_01752_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__xnor2_1 _08836_ (.A(_01740_),
    .B(_01749_),
    .Y(_01756_));
 sky130_fd_sc_hd__a21bo_1 _08837_ (.A1(_01755_),
    .A2(_01756_),
    .B1_N(_01750_),
    .X(_01757_));
 sky130_fd_sc_hd__xnor2_1 _08838_ (.A(_01736_),
    .B(_01738_),
    .Y(_01758_));
 sky130_fd_sc_hd__and2b_1 _08839_ (.A_N(_01758_),
    .B(_01757_),
    .X(_01759_));
 sky130_fd_sc_hd__o21ai_1 _08840_ (.A1(_01739_),
    .A2(_01759_),
    .B1(_01735_),
    .Y(_01760_));
 sky130_fd_sc_hd__a21oi_1 _08841_ (.A1(_01712_),
    .A2(_01733_),
    .B1(_01709_),
    .Y(_01761_));
 sky130_fd_sc_hd__a21o_1 _08842_ (.A1(_01712_),
    .A2(_01733_),
    .B1(_01709_),
    .X(_01762_));
 sky130_fd_sc_hd__or3_1 _08843_ (.A(_01735_),
    .B(_01739_),
    .C(_01759_),
    .X(_01763_));
 sky130_fd_sc_hd__and2_1 _08844_ (.A(_01760_),
    .B(_01763_),
    .X(_01764_));
 sky130_fd_sc_hd__nor2_1 _08845_ (.A(_01727_),
    .B(_01729_),
    .Y(_01765_));
 sky130_fd_sc_hd__or2_1 _08846_ (.A(_01730_),
    .B(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__xnor2_1 _08847_ (.A(_01755_),
    .B(_01756_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _08848_ (.A(_01766_),
    .B(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__xor2_1 _08849_ (.A(_01766_),
    .B(_01767_),
    .X(_01769_));
 sky130_fd_sc_hd__xor2_2 _08850_ (.A(_01747_),
    .B(_01748_),
    .X(_01770_));
 sky130_fd_sc_hd__nand2_1 _08851_ (.A(net156),
    .B(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__a22o_1 _08852_ (.A1(_00158_),
    .A2(_00266_),
    .B1(_00287_),
    .B2(_00159_),
    .X(_01772_));
 sky130_fd_sc_hd__xnor2_1 _08853_ (.A(net200),
    .B(_01772_),
    .Y(_01773_));
 sky130_fd_sc_hd__o22a_1 _08854_ (.A1(net285),
    .A2(net113),
    .B1(net106),
    .B2(net236),
    .X(_01774_));
 sky130_fd_sc_hd__xnor2_1 _08855_ (.A(net199),
    .B(_01774_),
    .Y(_01775_));
 sky130_fd_sc_hd__nand2b_1 _08856_ (.A_N(_01773_),
    .B(_01775_),
    .Y(_01776_));
 sky130_fd_sc_hd__xnor2_2 _08857_ (.A(net156),
    .B(_01770_),
    .Y(_01777_));
 sky130_fd_sc_hd__o21ai_1 _08858_ (.A1(_01776_),
    .A2(_01777_),
    .B1(_01771_),
    .Y(_01778_));
 sky130_fd_sc_hd__and2_1 _08859_ (.A(_01769_),
    .B(_01778_),
    .X(_01779_));
 sky130_fd_sc_hd__xnor2_1 _08860_ (.A(_01757_),
    .B(_01758_),
    .Y(_01780_));
 sky130_fd_sc_hd__or3_1 _08861_ (.A(_01768_),
    .B(_01779_),
    .C(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__and2_1 _08862_ (.A(_01752_),
    .B(_01754_),
    .X(_01782_));
 sky130_fd_sc_hd__nor2_1 _08863_ (.A(_01755_),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__xor2_2 _08864_ (.A(_01776_),
    .B(_01777_),
    .X(_01784_));
 sky130_fd_sc_hd__nand2_1 _08865_ (.A(_01783_),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__o22a_1 _08866_ (.A1(net157),
    .A2(net125),
    .B1(net149),
    .B2(net132),
    .X(_01786_));
 sky130_fd_sc_hd__xnor2_2 _08867_ (.A(net200),
    .B(_01786_),
    .Y(_01787_));
 sky130_fd_sc_hd__o22a_1 _08868_ (.A1(net236),
    .A2(net124),
    .B1(net106),
    .B2(net285),
    .X(_01788_));
 sky130_fd_sc_hd__xnor2_2 _08869_ (.A(net199),
    .B(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__a22o_1 _08870_ (.A1(_06702_),
    .A2(net150),
    .B1(_00340_),
    .B2(_06726_),
    .X(_01790_));
 sky130_fd_sc_hd__xnor2_1 _08871_ (.A(net181),
    .B(_01790_),
    .Y(_01791_));
 sky130_fd_sc_hd__nand3_2 _08872_ (.A(_01787_),
    .B(_01789_),
    .C(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__o22a_1 _08873_ (.A1(net208),
    .A2(net104),
    .B1(net130),
    .B2(net152),
    .X(_01793_));
 sky130_fd_sc_hd__xnor2_1 _08874_ (.A(net175),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__a21o_1 _08875_ (.A1(_01787_),
    .A2(_01789_),
    .B1(_01791_),
    .X(_01795_));
 sky130_fd_sc_hd__nand3_1 _08876_ (.A(_01792_),
    .B(_01794_),
    .C(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__nand2_2 _08877_ (.A(_01792_),
    .B(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__inv_2 _08878_ (.A(_01797_),
    .Y(_01798_));
 sky130_fd_sc_hd__xnor2_2 _08879_ (.A(_01783_),
    .B(_01784_),
    .Y(_01799_));
 sky130_fd_sc_hd__o21ai_1 _08880_ (.A1(_01798_),
    .A2(_01799_),
    .B1(_01785_),
    .Y(_01800_));
 sky130_fd_sc_hd__xor2_1 _08881_ (.A(_01769_),
    .B(_01778_),
    .X(_01801_));
 sky130_fd_sc_hd__and2_1 _08882_ (.A(_01800_),
    .B(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__o21a_1 _08883_ (.A1(_01768_),
    .A2(_01779_),
    .B1(_01780_),
    .X(_01803_));
 sky130_fd_sc_hd__o21ai_1 _08884_ (.A1(_01768_),
    .A2(_01779_),
    .B1(_01780_),
    .Y(_01804_));
 sky130_fd_sc_hd__or2_1 _08885_ (.A(_01800_),
    .B(_01801_),
    .X(_01805_));
 sky130_fd_sc_hd__and2b_1 _08886_ (.A_N(_01802_),
    .B(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__xnor2_1 _08887_ (.A(_01773_),
    .B(_01775_),
    .Y(_01807_));
 sky130_fd_sc_hd__a21o_1 _08888_ (.A1(_01792_),
    .A2(_01795_),
    .B1(_01794_),
    .X(_01808_));
 sky130_fd_sc_hd__and3_1 _08889_ (.A(_01796_),
    .B(_01807_),
    .C(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__a21oi_1 _08890_ (.A1(_01796_),
    .A2(_01808_),
    .B1(_01807_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _08891_ (.A(net208),
    .B(net130),
    .Y(_01811_));
 sky130_fd_sc_hd__a22o_1 _08892_ (.A1(_06702_),
    .A2(_00319_),
    .B1(net150),
    .B2(_06726_),
    .X(_01812_));
 sky130_fd_sc_hd__xnor2_1 _08893_ (.A(net181),
    .B(_01812_),
    .Y(_01813_));
 sky130_fd_sc_hd__and2b_1 _08894_ (.A_N(_01813_),
    .B(_01811_),
    .X(_01814_));
 sky130_fd_sc_hd__nor2_1 _08895_ (.A(net175),
    .B(_01811_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor4_1 _08896_ (.A(_01809_),
    .B(_01810_),
    .C(_01814_),
    .D(_01815_),
    .Y(_01816_));
 sky130_fd_sc_hd__or2_1 _08897_ (.A(_01809_),
    .B(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__xnor2_2 _08898_ (.A(_01797_),
    .B(_01799_),
    .Y(_01818_));
 sky130_fd_sc_hd__or2_1 _08899_ (.A(_01817_),
    .B(_01818_),
    .X(_01819_));
 sky130_fd_sc_hd__and2_1 _08900_ (.A(_01817_),
    .B(_01818_),
    .X(_01820_));
 sky130_fd_sc_hd__xor2_1 _08901_ (.A(_01787_),
    .B(_01789_),
    .X(_01821_));
 sky130_fd_sc_hd__xnor2_1 _08902_ (.A(_01811_),
    .B(_01813_),
    .Y(_01822_));
 sky130_fd_sc_hd__nand2b_1 _08903_ (.A_N(_01822_),
    .B(_01821_),
    .Y(_01823_));
 sky130_fd_sc_hd__a22o_1 _08904_ (.A1(_00158_),
    .A2(net150),
    .B1(_00340_),
    .B2(_00159_),
    .X(_01824_));
 sky130_fd_sc_hd__xnor2_1 _08905_ (.A(net200),
    .B(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__a21o_1 _08906_ (.A1(_00284_),
    .A2(_00285_),
    .B1(net285),
    .X(_01826_));
 sky130_fd_sc_hd__or3_1 _08907_ (.A(net236),
    .B(_00264_),
    .C(_00265_),
    .X(_01827_));
 sky130_fd_sc_hd__and3_1 _08908_ (.A(net197),
    .B(_01826_),
    .C(_01827_),
    .X(_01828_));
 sky130_fd_sc_hd__a21oi_1 _08909_ (.A1(_01826_),
    .A2(_01827_),
    .B1(net197),
    .Y(_01829_));
 sky130_fd_sc_hd__or3_2 _08910_ (.A(_01825_),
    .B(_01828_),
    .C(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__xor2_1 _08911_ (.A(_01821_),
    .B(_01822_),
    .X(_01831_));
 sky130_fd_sc_hd__or2_1 _08912_ (.A(_01830_),
    .B(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__o22a_1 _08913_ (.A1(_01809_),
    .A2(_01810_),
    .B1(_01814_),
    .B2(_01815_),
    .X(_01833_));
 sky130_fd_sc_hd__a211o_1 _08914_ (.A1(_01823_),
    .A2(_01832_),
    .B1(_01833_),
    .C1(_01816_),
    .X(_01834_));
 sky130_fd_sc_hd__o211ai_2 _08915_ (.A1(_01816_),
    .A2(_01833_),
    .B1(_01832_),
    .C1(_01823_),
    .Y(_01835_));
 sky130_fd_sc_hd__xor2_1 _08916_ (.A(_01830_),
    .B(_01831_),
    .X(_01836_));
 sky130_fd_sc_hd__o21ai_1 _08917_ (.A1(_01828_),
    .A2(_01829_),
    .B1(_01825_),
    .Y(_01837_));
 sky130_fd_sc_hd__a22o_1 _08918_ (.A1(net206),
    .A2(_06702_),
    .B1(_06726_),
    .B2(_00319_),
    .X(_01838_));
 sky130_fd_sc_hd__xnor2_1 _08919_ (.A(net181),
    .B(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__nand3_2 _08920_ (.A(_01830_),
    .B(_01837_),
    .C(_01839_),
    .Y(_01840_));
 sky130_fd_sc_hd__a22o_1 _08921_ (.A1(_00158_),
    .A2(_00319_),
    .B1(net150),
    .B2(_00159_),
    .X(_01841_));
 sky130_fd_sc_hd__xnor2_1 _08922_ (.A(net200),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__o32ai_2 _08923_ (.A1(net285),
    .A2(_00264_),
    .A3(_00265_),
    .B1(net149),
    .B2(net236),
    .Y(_01843_));
 sky130_fd_sc_hd__xnor2_1 _08924_ (.A(net197),
    .B(_01843_),
    .Y(_01844_));
 sky130_fd_sc_hd__nand2b_1 _08925_ (.A_N(_01842_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__inv_2 _08926_ (.A(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__a21o_1 _08927_ (.A1(_01830_),
    .A2(_01837_),
    .B1(_01839_),
    .X(_01847_));
 sky130_fd_sc_hd__nand3_2 _08928_ (.A(_01840_),
    .B(_01846_),
    .C(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__and3b_1 _08929_ (.A_N(_01836_),
    .B(_01840_),
    .C(_01848_),
    .X(_01849_));
 sky130_fd_sc_hd__a21bo_1 _08930_ (.A1(_01840_),
    .A2(_01848_),
    .B1_N(_01836_),
    .X(_01850_));
 sky130_fd_sc_hd__xor2_1 _08931_ (.A(_01842_),
    .B(_01844_),
    .X(_01851_));
 sky130_fd_sc_hd__nand2_1 _08932_ (.A(net206),
    .B(_06726_),
    .Y(_01852_));
 sky130_fd_sc_hd__and3_1 _08933_ (.A(net207),
    .B(_06726_),
    .C(_01851_),
    .X(_01853_));
 sky130_fd_sc_hd__a21oi_1 _08934_ (.A1(net181),
    .A2(_01852_),
    .B1(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__a21o_1 _08935_ (.A1(_01840_),
    .A2(_01847_),
    .B1(_01846_),
    .X(_01855_));
 sky130_fd_sc_hd__a21oi_1 _08936_ (.A1(_01848_),
    .A2(_01855_),
    .B1(_01854_),
    .Y(_01856_));
 sky130_fd_sc_hd__a21o_1 _08937_ (.A1(_01848_),
    .A2(_01855_),
    .B1(_01854_),
    .X(_01857_));
 sky130_fd_sc_hd__and3_1 _08938_ (.A(_01848_),
    .B(_01854_),
    .C(_01855_),
    .X(_01858_));
 sky130_fd_sc_hd__a22o_1 _08939_ (.A1(net207),
    .A2(_00158_),
    .B1(_00159_),
    .B2(_00319_),
    .X(_01859_));
 sky130_fd_sc_hd__xnor2_1 _08940_ (.A(net200),
    .B(_01859_),
    .Y(_01860_));
 sky130_fd_sc_hd__a22o_1 _08941_ (.A1(_00138_),
    .A2(net150),
    .B1(_00340_),
    .B2(net291),
    .X(_01861_));
 sky130_fd_sc_hd__xnor2_1 _08942_ (.A(net197),
    .B(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2b_1 _08943_ (.A_N(_01860_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__xnor2_1 _08944_ (.A(_01851_),
    .B(_01852_),
    .Y(_01864_));
 sky130_fd_sc_hd__nor2_1 _08945_ (.A(_01863_),
    .B(_01864_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _08946_ (.A(_01863_),
    .B(_01864_),
    .Y(_01866_));
 sky130_fd_sc_hd__nand2b_1 _08947_ (.A_N(_01865_),
    .B(_01866_),
    .Y(_01867_));
 sky130_fd_sc_hd__a22o_1 _08948_ (.A1(_00138_),
    .A2(_00319_),
    .B1(net150),
    .B2(net291),
    .X(_01868_));
 sky130_fd_sc_hd__xnor2_2 _08949_ (.A(net197),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_1 _08950_ (.A(net209),
    .B(net157),
    .Y(_01870_));
 sky130_fd_sc_hd__xnor2_1 _08951_ (.A(net201),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__nand2_1 _08952_ (.A(_01869_),
    .B(_01871_),
    .Y(_01872_));
 sky130_fd_sc_hd__xnor2_1 _08953_ (.A(_01869_),
    .B(_01871_),
    .Y(_01873_));
 sky130_fd_sc_hd__xnor2_1 _08954_ (.A(_01869_),
    .B(_01870_),
    .Y(_01874_));
 sky130_fd_sc_hd__o2bb2a_1 _08955_ (.A1_N(net289),
    .A2_N(_06578_),
    .B1(_00320_),
    .B2(net285),
    .X(_01875_));
 sky130_fd_sc_hd__and2_1 _08956_ (.A(_06637_),
    .B(_01875_),
    .X(_01876_));
 sky130_fd_sc_hd__nand2_1 _08957_ (.A(net199),
    .B(_01876_),
    .Y(_01877_));
 sky130_fd_sc_hd__nor2_1 _08958_ (.A(_01874_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__xnor2_1 _08959_ (.A(_01860_),
    .B(_01862_),
    .Y(_01879_));
 sky130_fd_sc_hd__xnor2_1 _08960_ (.A(_01872_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__o21ai_1 _08961_ (.A1(net201),
    .A2(_01873_),
    .B1(_01872_),
    .Y(_01881_));
 sky130_fd_sc_hd__a22o_1 _08962_ (.A1(_01878_),
    .A2(_01880_),
    .B1(_01881_),
    .B2(_01879_),
    .X(_01882_));
 sky130_fd_sc_hd__a21o_1 _08963_ (.A1(_01866_),
    .A2(_01882_),
    .B1(_01865_),
    .X(_01883_));
 sky130_fd_sc_hd__nor2_1 _08964_ (.A(_01856_),
    .B(_01858_),
    .Y(_01884_));
 sky130_fd_sc_hd__a21oi_1 _08965_ (.A1(_01857_),
    .A2(_01883_),
    .B1(_01858_),
    .Y(_01885_));
 sky130_fd_sc_hd__a21o_1 _08966_ (.A1(_01850_),
    .A2(_01885_),
    .B1(_01849_),
    .X(_01886_));
 sky130_fd_sc_hd__and2b_1 _08967_ (.A_N(_01849_),
    .B(_01850_),
    .X(_01887_));
 sky130_fd_sc_hd__a21boi_2 _08968_ (.A1(_01834_),
    .A2(_01886_),
    .B1_N(_01835_),
    .Y(_01888_));
 sky130_fd_sc_hd__a21o_1 _08969_ (.A1(_01817_),
    .A2(_01818_),
    .B1(_01888_),
    .X(_01889_));
 sky130_fd_sc_hd__xor2_1 _08970_ (.A(_01817_),
    .B(_01818_),
    .X(_01890_));
 sky130_fd_sc_hd__nand2_1 _08971_ (.A(_01819_),
    .B(_01889_),
    .Y(_01891_));
 sky130_fd_sc_hd__a311o_1 _08972_ (.A1(_01805_),
    .A2(_01819_),
    .A3(_01889_),
    .B1(_01803_),
    .C1(_01802_),
    .X(_01892_));
 sky130_fd_sc_hd__and2_1 _08973_ (.A(_01781_),
    .B(_01804_),
    .X(_01893_));
 sky130_fd_sc_hd__nand2_1 _08974_ (.A(_01781_),
    .B(_01892_),
    .Y(_01894_));
 sky130_fd_sc_hd__a21oi_1 _08975_ (.A1(_01760_),
    .A2(_01762_),
    .B1(_01734_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_2 _08976_ (.A(_01734_),
    .B(_01761_),
    .Y(_01896_));
 sky130_fd_sc_hd__a41o_1 _08977_ (.A1(_01764_),
    .A2(_01781_),
    .A3(_01892_),
    .A4(_01896_),
    .B1(_01895_),
    .X(_01897_));
 sky130_fd_sc_hd__a32o_2 _08978_ (.A1(_01706_),
    .A2(_01708_),
    .A3(_01897_),
    .B1(_01705_),
    .B2(_01680_),
    .X(_01898_));
 sky130_fd_sc_hd__a32o_1 _08979_ (.A1(_01644_),
    .A2(_01646_),
    .A3(_01898_),
    .B1(_01643_),
    .B2(_01615_),
    .X(_01899_));
 sky130_fd_sc_hd__xor2_1 _08980_ (.A(_01493_),
    .B(_01537_),
    .X(_01900_));
 sky130_fd_sc_hd__nand2_1 _08981_ (.A(_01538_),
    .B(_01539_),
    .Y(_01901_));
 sky130_fd_sc_hd__and3_1 _08982_ (.A(_01543_),
    .B(_01574_),
    .C(_01575_),
    .X(_01902_));
 sky130_fd_sc_hd__nor2_1 _08983_ (.A(_01576_),
    .B(_01902_),
    .Y(_01903_));
 sky130_fd_sc_hd__a32o_2 _08984_ (.A1(_01899_),
    .A2(_01900_),
    .A3(_01903_),
    .B1(_01577_),
    .B2(_01538_),
    .X(_01904_));
 sky130_fd_sc_hd__a21o_1 _08985_ (.A1(_01492_),
    .A2(_01904_),
    .B1(_01488_),
    .X(_01905_));
 sky130_fd_sc_hd__or3b_1 _08986_ (.A(_01390_),
    .B(_01391_),
    .C_N(_01488_),
    .X(_01906_));
 sky130_fd_sc_hd__or4bb_1 _08987_ (.A(_01390_),
    .B(_01391_),
    .C_N(_01492_),
    .D_N(_01904_),
    .X(_01907_));
 sky130_fd_sc_hd__and3_1 _08988_ (.A(_01388_),
    .B(_01906_),
    .C(_01907_),
    .X(_01908_));
 sky130_fd_sc_hd__a311o_1 _08989_ (.A1(_01388_),
    .A2(_01906_),
    .A3(_01907_),
    .B1(_01285_),
    .C1(_01284_),
    .X(_01909_));
 sky130_fd_sc_hd__nand2_2 _08990_ (.A(_01282_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__a21o_1 _08991_ (.A1(_01282_),
    .A2(_01909_),
    .B1(_01158_),
    .X(_01911_));
 sky130_fd_sc_hd__a21o_1 _08992_ (.A1(_01030_),
    .A2(_01085_),
    .B1(_01086_),
    .X(_01912_));
 sky130_fd_sc_hd__and2_1 _08993_ (.A(_01157_),
    .B(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__nand2b_1 _08994_ (.A_N(_01087_),
    .B(_01912_),
    .Y(_01914_));
 sky130_fd_sc_hd__a21oi_4 _08995_ (.A1(_01911_),
    .A2(_01913_),
    .B1(_01087_),
    .Y(_01915_));
 sky130_fd_sc_hd__nor2_1 _08996_ (.A(_01023_),
    .B(_01024_),
    .Y(_01916_));
 sky130_fd_sc_hd__xnor2_4 _08997_ (.A(_01023_),
    .B(_01024_),
    .Y(_01917_));
 sky130_fd_sc_hd__and2b_1 _08998_ (.A_N(_00955_),
    .B(_01026_),
    .X(_01918_));
 sky130_fd_sc_hd__xnor2_2 _08999_ (.A(_00883_),
    .B(_00954_),
    .Y(_01919_));
 sky130_fd_sc_hd__a2111o_1 _09000_ (.A1(_01911_),
    .A2(_01913_),
    .B1(_01917_),
    .C1(_01919_),
    .D1(_01087_),
    .X(_01920_));
 sky130_fd_sc_hd__nand2_1 _09001_ (.A(_01027_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__xnor2_2 _09002_ (.A(_00882_),
    .B(_01921_),
    .Y(_01922_));
 sky130_fd_sc_hd__xnor2_4 _09003_ (.A(_01158_),
    .B(_01910_),
    .Y(_01923_));
 sky130_fd_sc_hd__and2_1 _09004_ (.A(_01874_),
    .B(_01877_),
    .X(_01924_));
 sky130_fd_sc_hd__nor2_1 _09005_ (.A(_01878_),
    .B(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__nand2b_1 _09006_ (.A_N(_01925_),
    .B(_01876_),
    .Y(_01926_));
 sky130_fd_sc_hd__o21ba_1 _09007_ (.A1(net201),
    .A2(_01873_),
    .B1_N(_01878_),
    .X(_01927_));
 sky130_fd_sc_hd__xnor2_1 _09008_ (.A(_01880_),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__nor2_1 _09009_ (.A(_01926_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__xor2_2 _09010_ (.A(_01867_),
    .B(_01882_),
    .X(_01930_));
 sky130_fd_sc_hd__nand2_1 _09011_ (.A(_01929_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__xor2_2 _09012_ (.A(_01883_),
    .B(_01884_),
    .X(_01932_));
 sky130_fd_sc_hd__xor2_1 _09013_ (.A(_01885_),
    .B(_01887_),
    .X(_01933_));
 sky130_fd_sc_hd__and4b_1 _09014_ (.A_N(_01932_),
    .B(_01929_),
    .C(_01930_),
    .D(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__a21oi_1 _09015_ (.A1(_01834_),
    .A2(_01835_),
    .B1(_01886_),
    .Y(_01935_));
 sky130_fd_sc_hd__and3_1 _09016_ (.A(_01834_),
    .B(_01835_),
    .C(_01886_),
    .X(_01936_));
 sky130_fd_sc_hd__nor2_1 _09017_ (.A(_01935_),
    .B(_01936_),
    .Y(_01937_));
 sky130_fd_sc_hd__and2_1 _09018_ (.A(_01934_),
    .B(_01937_),
    .X(_01938_));
 sky130_fd_sc_hd__xnor2_1 _09019_ (.A(_01888_),
    .B(_01890_),
    .Y(_01939_));
 sky130_fd_sc_hd__and2_1 _09020_ (.A(_01938_),
    .B(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__xor2_2 _09021_ (.A(_01806_),
    .B(_01891_),
    .X(_01941_));
 sky130_fd_sc_hd__a211o_1 _09022_ (.A1(_01888_),
    .A2(_01890_),
    .B1(_01802_),
    .C1(_01820_),
    .X(_01942_));
 sky130_fd_sc_hd__and3_1 _09023_ (.A(_01805_),
    .B(_01893_),
    .C(_01942_),
    .X(_01943_));
 sky130_fd_sc_hd__a21oi_1 _09024_ (.A1(_01805_),
    .A2(_01942_),
    .B1(_01893_),
    .Y(_01944_));
 sky130_fd_sc_hd__or2_1 _09025_ (.A(_01943_),
    .B(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__o211a_1 _09026_ (.A1(_01943_),
    .A2(_01944_),
    .B1(_01940_),
    .C1(_01941_),
    .X(_01946_));
 sky130_fd_sc_hd__xnor2_1 _09027_ (.A(_01764_),
    .B(_01894_),
    .Y(_01947_));
 sky130_fd_sc_hd__xor2_1 _09028_ (.A(_01764_),
    .B(_01894_),
    .X(_01948_));
 sky130_fd_sc_hd__a21boi_1 _09029_ (.A1(_01760_),
    .A2(_01804_),
    .B1_N(_01763_),
    .Y(_01949_));
 sky130_fd_sc_hd__a41o_1 _09030_ (.A1(_01764_),
    .A2(_01805_),
    .A3(_01893_),
    .A4(_01942_),
    .B1(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__xor2_2 _09031_ (.A(_01896_),
    .B(_01950_),
    .X(_01951_));
 sky130_fd_sc_hd__or3b_1 _09032_ (.A(_01947_),
    .B(_01951_),
    .C_N(_01946_),
    .X(_01952_));
 sky130_fd_sc_hd__xor2_2 _09033_ (.A(_01708_),
    .B(_01897_),
    .X(_01953_));
 sky130_fd_sc_hd__or4b_1 _09034_ (.A(_01947_),
    .B(_01951_),
    .C(_01953_),
    .D_N(_01946_),
    .X(_01954_));
 sky130_fd_sc_hd__a21o_1 _09035_ (.A1(_01703_),
    .A2(_01704_),
    .B1(_01761_),
    .X(_01955_));
 sky130_fd_sc_hd__a21o_1 _09036_ (.A1(_01896_),
    .A2(_01950_),
    .B1(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__a21oi_1 _09037_ (.A1(_01707_),
    .A2(_01956_),
    .B1(_01706_),
    .Y(_01957_));
 sky130_fd_sc_hd__and3_1 _09038_ (.A(_01706_),
    .B(_01707_),
    .C(_01956_),
    .X(_01958_));
 sky130_fd_sc_hd__or2_1 _09039_ (.A(_01957_),
    .B(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__o21ba_2 _09040_ (.A1(_01957_),
    .A2(_01958_),
    .B1_N(_01954_),
    .X(_01960_));
 sky130_fd_sc_hd__xnor2_4 _09041_ (.A(_01646_),
    .B(_01898_),
    .Y(_01961_));
 sky130_fd_sc_hd__a2bb2o_1 _09042_ (.A1_N(_01647_),
    .A2_N(_01679_),
    .B1(_01641_),
    .B2(_01642_),
    .X(_01962_));
 sky130_fd_sc_hd__o21ai_2 _09043_ (.A1(_01641_),
    .A2(_01642_),
    .B1(_01962_),
    .Y(_01963_));
 sky130_fd_sc_hd__nand4_4 _09044_ (.A(_01646_),
    .B(_01706_),
    .C(_01707_),
    .D(_01956_),
    .Y(_01964_));
 sky130_fd_sc_hd__a21oi_2 _09045_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01645_),
    .Y(_01965_));
 sky130_fd_sc_hd__and3_1 _09046_ (.A(_01645_),
    .B(_01963_),
    .C(_01964_),
    .X(_01966_));
 sky130_fd_sc_hd__or2_1 _09047_ (.A(_01965_),
    .B(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__and3_1 _09048_ (.A(_01960_),
    .B(_01961_),
    .C(_01967_),
    .X(_01968_));
 sky130_fd_sc_hd__xnor2_2 _09049_ (.A(_01899_),
    .B(_01903_),
    .Y(_01969_));
 sky130_fd_sc_hd__o2111ai_4 _09050_ (.A1(_01965_),
    .A2(_01966_),
    .B1(_01969_),
    .C1(_01961_),
    .D1(_01960_),
    .Y(_01970_));
 sky130_fd_sc_hd__and2b_1 _09051_ (.A_N(_01576_),
    .B(_01616_),
    .X(_01971_));
 sky130_fd_sc_hd__or2_1 _09052_ (.A(_01902_),
    .B(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__a2111o_1 _09053_ (.A1(_01963_),
    .A2(_01964_),
    .B1(_01576_),
    .C1(_01645_),
    .D1(_01902_),
    .X(_01973_));
 sky130_fd_sc_hd__a21o_1 _09054_ (.A1(_01972_),
    .A2(_01973_),
    .B1(_01901_),
    .X(_01974_));
 sky130_fd_sc_hd__nand3_2 _09055_ (.A(_01901_),
    .B(_01972_),
    .C(_01973_),
    .Y(_01975_));
 sky130_fd_sc_hd__a21oi_4 _09056_ (.A1(_01974_),
    .A2(_01975_),
    .B1(_01970_),
    .Y(_01976_));
 sky130_fd_sc_hd__xor2_4 _09057_ (.A(_01491_),
    .B(_01904_),
    .X(_01977_));
 sky130_fd_sc_hd__a21o_1 _09058_ (.A1(_01486_),
    .A2(_01539_),
    .B1(_01490_),
    .X(_01978_));
 sky130_fd_sc_hd__a211o_1 _09059_ (.A1(_01972_),
    .A2(_01973_),
    .B1(_01491_),
    .C1(_01901_),
    .X(_01979_));
 sky130_fd_sc_hd__and3_1 _09060_ (.A(_01489_),
    .B(_01978_),
    .C(_01979_),
    .X(_01980_));
 sky130_fd_sc_hd__a21oi_1 _09061_ (.A1(_01978_),
    .A2(_01979_),
    .B1(_01489_),
    .Y(_01981_));
 sky130_fd_sc_hd__nor2_1 _09062_ (.A(_01980_),
    .B(_01981_),
    .Y(_01982_));
 sky130_fd_sc_hd__nand3b_1 _09063_ (.A_N(_01982_),
    .B(_01976_),
    .C(_01977_),
    .Y(_01983_));
 sky130_fd_sc_hd__xnor2_2 _09064_ (.A(_01390_),
    .B(_01905_),
    .Y(_01984_));
 sky130_fd_sc_hd__xor2_1 _09065_ (.A(_01390_),
    .B(_01905_),
    .X(_01985_));
 sky130_fd_sc_hd__nor2_1 _09066_ (.A(_01983_),
    .B(_01984_),
    .Y(_01986_));
 sky130_fd_sc_hd__o2111ai_2 _09067_ (.A1(_01980_),
    .A2(_01981_),
    .B1(_01985_),
    .C1(_01977_),
    .D1(_01976_),
    .Y(_01987_));
 sky130_fd_sc_hd__or2_1 _09068_ (.A(_01390_),
    .B(_01489_),
    .X(_01988_));
 sky130_fd_sc_hd__a21o_1 _09069_ (.A1(_01978_),
    .A2(_01979_),
    .B1(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__a21o_1 _09070_ (.A1(_01387_),
    .A2(_01487_),
    .B1(_01389_),
    .X(_01990_));
 sky130_fd_sc_hd__nand3_1 _09071_ (.A(_01391_),
    .B(_01989_),
    .C(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__a21o_1 _09072_ (.A1(_01989_),
    .A2(_01990_),
    .B1(_01391_),
    .X(_01992_));
 sky130_fd_sc_hd__nand2_1 _09073_ (.A(_01991_),
    .B(_01992_),
    .Y(_01993_));
 sky130_fd_sc_hd__xor2_1 _09074_ (.A(_01284_),
    .B(_01908_),
    .X(_01994_));
 sky130_fd_sc_hd__a211o_1 _09075_ (.A1(_01991_),
    .A2(_01992_),
    .B1(_01994_),
    .C1(_01987_),
    .X(_01995_));
 sky130_fd_sc_hd__a21o_1 _09076_ (.A1(_01281_),
    .A2(_01333_),
    .B1(_01283_),
    .X(_01996_));
 sky130_fd_sc_hd__or2_1 _09077_ (.A(_01284_),
    .B(_01391_),
    .X(_01997_));
 sky130_fd_sc_hd__a211o_1 _09078_ (.A1(_01978_),
    .A2(_01979_),
    .B1(_01988_),
    .C1(_01997_),
    .X(_01998_));
 sky130_fd_sc_hd__or2_1 _09079_ (.A(_01990_),
    .B(_01997_),
    .X(_01999_));
 sky130_fd_sc_hd__and3_1 _09080_ (.A(_01996_),
    .B(_01998_),
    .C(_01999_),
    .X(_02000_));
 sky130_fd_sc_hd__xor2_2 _09081_ (.A(_01285_),
    .B(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__or3_1 _09082_ (.A(_01923_),
    .B(_01995_),
    .C(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__a21o_1 _09083_ (.A1(_01157_),
    .A2(_01219_),
    .B1(_01156_),
    .X(_02003_));
 sky130_fd_sc_hd__a311o_2 _09084_ (.A1(_01996_),
    .A2(_01998_),
    .A3(_01999_),
    .B1(_01285_),
    .C1(_01158_),
    .X(_02004_));
 sky130_fd_sc_hd__a21o_1 _09085_ (.A1(_02003_),
    .A2(_02004_),
    .B1(_01914_),
    .X(_02005_));
 sky130_fd_sc_hd__nand3_1 _09086_ (.A(_01914_),
    .B(_02003_),
    .C(_02004_),
    .Y(_02006_));
 sky130_fd_sc_hd__and2_1 _09087_ (.A(_02005_),
    .B(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__a2111o_1 _09088_ (.A1(_02005_),
    .A2(_02006_),
    .B1(_01923_),
    .C1(_01995_),
    .D1(_02001_),
    .X(_02008_));
 sky130_fd_sc_hd__xor2_2 _09089_ (.A(_01915_),
    .B(_01917_),
    .X(_02009_));
 sky130_fd_sc_hd__nand2b_1 _09090_ (.A_N(_02008_),
    .B(_02009_),
    .Y(_02010_));
 sky130_fd_sc_hd__a21o_1 _09091_ (.A1(_01025_),
    .A2(_01912_),
    .B1(_01916_),
    .X(_02011_));
 sky130_fd_sc_hd__or2_1 _09092_ (.A(_01914_),
    .B(_01917_),
    .X(_02012_));
 sky130_fd_sc_hd__a211o_1 _09093_ (.A1(_02003_),
    .A2(_02004_),
    .B1(_01914_),
    .C1(_01917_),
    .X(_02013_));
 sky130_fd_sc_hd__and3_1 _09094_ (.A(_01918_),
    .B(_02011_),
    .C(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__a21oi_1 _09095_ (.A1(_02011_),
    .A2(_02013_),
    .B1(_01918_),
    .Y(_02015_));
 sky130_fd_sc_hd__a21o_1 _09096_ (.A1(_02011_),
    .A2(_02013_),
    .B1(_01918_),
    .X(_02016_));
 sky130_fd_sc_hd__or4bb_1 _09097_ (.A(_02014_),
    .B(_02008_),
    .C_N(_02009_),
    .D_N(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__nor2_1 _09098_ (.A(_01922_),
    .B(_02017_),
    .Y(_02018_));
 sky130_fd_sc_hd__a21oi_4 _09099_ (.A1(_00773_),
    .A2(_00878_),
    .B1(_00877_),
    .Y(_02019_));
 sky130_fd_sc_hd__o21ai_4 _09100_ (.A1(_00872_),
    .A2(_00873_),
    .B1(_00875_),
    .Y(_02020_));
 sky130_fd_sc_hd__a21oi_2 _09101_ (.A1(_00820_),
    .A2(_00831_),
    .B1(_00830_),
    .Y(_02021_));
 sky130_fd_sc_hd__a22o_1 _09102_ (.A1(_00287_),
    .A2(net14),
    .B1(net30),
    .B2(net107),
    .X(_02022_));
 sky130_fd_sc_hd__xnor2_1 _09103_ (.A(net92),
    .B(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__o22a_1 _09104_ (.A1(net39),
    .A2(net113),
    .B1(net110),
    .B2(net37),
    .X(_02024_));
 sky130_fd_sc_hd__xnor2_1 _09105_ (.A(net99),
    .B(_02024_),
    .Y(_02025_));
 sky130_fd_sc_hd__o22a_1 _09106_ (.A1(_00267_),
    .A2(net33),
    .B1(_00339_),
    .B2(net35),
    .X(_02026_));
 sky130_fd_sc_hd__xnor2_1 _09107_ (.A(net95),
    .B(_02026_),
    .Y(_02027_));
 sky130_fd_sc_hd__xnor2_1 _09108_ (.A(_02025_),
    .B(_02027_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor2_1 _09109_ (.A(_02023_),
    .B(_02028_),
    .Y(_02029_));
 sky130_fd_sc_hd__and2_1 _09110_ (.A(_02023_),
    .B(_02028_),
    .X(_02030_));
 sky130_fd_sc_hd__or2_1 _09111_ (.A(_02029_),
    .B(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__a21oi_1 _09112_ (.A1(_00801_),
    .A2(_00803_),
    .B1(_02031_),
    .Y(_02032_));
 sky130_fd_sc_hd__and3_1 _09113_ (.A(_00801_),
    .B(_00803_),
    .C(_02031_),
    .X(_02033_));
 sky130_fd_sc_hd__nor2_1 _09114_ (.A(_02032_),
    .B(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__and2b_1 _09115_ (.A_N(_02021_),
    .B(_02034_),
    .X(_02035_));
 sky130_fd_sc_hd__xnor2_2 _09116_ (.A(_02021_),
    .B(_02034_),
    .Y(_02036_));
 sky130_fd_sc_hd__o21ai_2 _09117_ (.A1(_00822_),
    .A2(_00828_),
    .B1(_00827_),
    .Y(_02037_));
 sky130_fd_sc_hd__o21ba_1 _09118_ (.A1(_00806_),
    .A2(_00818_),
    .B1_N(_00817_),
    .X(_02038_));
 sky130_fd_sc_hd__xnor2_1 _09119_ (.A(_00856_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__nand2b_1 _09120_ (.A_N(_02039_),
    .B(_02037_),
    .Y(_02040_));
 sky130_fd_sc_hd__xnor2_1 _09121_ (.A(_02037_),
    .B(_02039_),
    .Y(_02041_));
 sky130_fd_sc_hd__a22o_1 _09122_ (.A1(_06725_),
    .A2(net129),
    .B1(net127),
    .B2(_06730_),
    .X(_02042_));
 sky130_fd_sc_hd__xnor2_2 _09123_ (.A(net154),
    .B(_02042_),
    .Y(_02043_));
 sky130_fd_sc_hd__o22a_1 _09124_ (.A1(net42),
    .A2(net68),
    .B1(net66),
    .B2(net40),
    .X(_02044_));
 sky130_fd_sc_hd__xnor2_2 _09125_ (.A(net146),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__o22a_1 _09126_ (.A1(net47),
    .A2(net105),
    .B1(net131),
    .B2(net45),
    .X(_02046_));
 sky130_fd_sc_hd__xnor2_2 _09127_ (.A(net174),
    .B(_02046_),
    .Y(_02047_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(_02045_),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__xnor2_2 _09129_ (.A(_02045_),
    .B(_02047_),
    .Y(_02049_));
 sky130_fd_sc_hd__xnor2_2 _09130_ (.A(_02043_),
    .B(_02049_),
    .Y(_02050_));
 sky130_fd_sc_hd__o22a_1 _09131_ (.A1(net24),
    .A2(net82),
    .B1(net76),
    .B2(net22),
    .X(_02051_));
 sky130_fd_sc_hd__xnor2_2 _09132_ (.A(net86),
    .B(_02051_),
    .Y(_02052_));
 sky130_fd_sc_hd__a22o_1 _09133_ (.A1(_00220_),
    .A2(_00461_),
    .B1(_00465_),
    .B2(_00229_),
    .X(_02053_));
 sky130_fd_sc_hd__xnor2_2 _09134_ (.A(_00431_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__xnor2_2 _09135_ (.A(_02052_),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__o22a_1 _09136_ (.A1(net83),
    .A2(net74),
    .B1(net70),
    .B2(net79),
    .X(_02056_));
 sky130_fd_sc_hd__xnor2_2 _09137_ (.A(net116),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2b_1 _09138_ (.A_N(_02055_),
    .B(_02057_),
    .Y(_02058_));
 sky130_fd_sc_hd__xnor2_2 _09139_ (.A(_02055_),
    .B(_02057_),
    .Y(_02059_));
 sky130_fd_sc_hd__o22a_2 _09140_ (.A1(_00157_),
    .A2(net44),
    .B1(_00517_),
    .B2(net157),
    .X(_02060_));
 sky130_fd_sc_hd__xnor2_4 _09141_ (.A(net202),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__o22a_2 _09142_ (.A1(_06727_),
    .A2(net51),
    .B1(net49),
    .B2(_06701_),
    .X(_02062_));
 sky130_fd_sc_hd__xnor2_4 _09143_ (.A(net179),
    .B(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__a31o_4 _09144_ (.A1(_05134_),
    .A2(_05211_),
    .A3(_00173_),
    .B1(net177),
    .X(_02064_));
 sky130_fd_sc_hd__xnor2_4 _09145_ (.A(_05069_),
    .B(_02064_),
    .Y(_02065_));
 sky130_fd_sc_hd__xnor2_4 _09146_ (.A(_05080_),
    .B(_02064_),
    .Y(_02066_));
 sky130_fd_sc_hd__a22o_1 _09147_ (.A1(_00138_),
    .A2(_00812_),
    .B1(net11),
    .B2(net291),
    .X(_02067_));
 sky130_fd_sc_hd__xnor2_4 _09148_ (.A(net198),
    .B(_02067_),
    .Y(_02068_));
 sky130_fd_sc_hd__nand2_1 _09149_ (.A(_02063_),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__xnor2_4 _09150_ (.A(_02063_),
    .B(_02068_),
    .Y(_02070_));
 sky130_fd_sc_hd__xor2_4 _09151_ (.A(_02061_),
    .B(_02070_),
    .X(_02071_));
 sky130_fd_sc_hd__nand2_1 _09152_ (.A(_02059_),
    .B(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__xnor2_2 _09153_ (.A(_02059_),
    .B(_02071_),
    .Y(_02073_));
 sky130_fd_sc_hd__xor2_1 _09154_ (.A(_02050_),
    .B(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__or3_4 _09155_ (.A(reg1_val[29]),
    .B(net288),
    .C(_00554_),
    .X(_02075_));
 sky130_fd_sc_hd__o21ai_1 _09156_ (.A1(reg1_val[29]),
    .A2(_00554_),
    .B1(net288),
    .Y(_02076_));
 sky130_fd_sc_hd__a21o_1 _09157_ (.A1(_02075_),
    .A2(_02076_),
    .B1(net258),
    .X(_02077_));
 sky130_fd_sc_hd__o21a_2 _09158_ (.A1(net288),
    .A2(net261),
    .B1(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__o211ai_2 _09159_ (.A1(net288),
    .A2(net261),
    .B1(_00787_),
    .C1(_02077_),
    .Y(_02079_));
 sky130_fd_sc_hd__xnor2_4 _09160_ (.A(net64),
    .B(_02078_),
    .Y(_02080_));
 sky130_fd_sc_hd__nand2_1 _09161_ (.A(net207),
    .B(net9),
    .Y(_02081_));
 sky130_fd_sc_hd__a22o_1 _09162_ (.A1(net150),
    .A2(net17),
    .B1(net13),
    .B2(net153),
    .X(_02082_));
 sky130_fd_sc_hd__xnor2_1 _09163_ (.A(net65),
    .B(_02082_),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_1 _09164_ (.A(_02081_),
    .B(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__and2_1 _09165_ (.A(_02081_),
    .B(_02083_),
    .X(_02085_));
 sky130_fd_sc_hd__or2_1 _09166_ (.A(_02084_),
    .B(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__and2_1 _09167_ (.A(_02074_),
    .B(_02086_),
    .X(_02087_));
 sky130_fd_sc_hd__xor2_1 _09168_ (.A(_02074_),
    .B(_02086_),
    .X(_02088_));
 sky130_fd_sc_hd__xor2_1 _09169_ (.A(_02041_),
    .B(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__a21o_1 _09170_ (.A1(_00776_),
    .A2(_00782_),
    .B1(_00781_),
    .X(_02090_));
 sky130_fd_sc_hd__o22a_1 _09171_ (.A1(net28),
    .A2(net115),
    .B1(net85),
    .B2(net26),
    .X(_02091_));
 sky130_fd_sc_hd__xnor2_1 _09172_ (.A(net90),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__o22a_1 _09173_ (.A1(net123),
    .A2(net21),
    .B1(net19),
    .B2(net119),
    .X(_02093_));
 sky130_fd_sc_hd__xnor2_1 _09174_ (.A(net96),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__nand2_2 _09175_ (.A(_02092_),
    .B(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__or2_1 _09176_ (.A(_02092_),
    .B(_02094_),
    .X(_02096_));
 sky130_fd_sc_hd__nand2_1 _09177_ (.A(_02095_),
    .B(_02096_),
    .Y(_02097_));
 sky130_fd_sc_hd__a21oi_1 _09178_ (.A1(_00840_),
    .A2(_00843_),
    .B1(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__and3_1 _09179_ (.A(_00840_),
    .B(_00843_),
    .C(_02097_),
    .X(_02099_));
 sky130_fd_sc_hd__or2_1 _09180_ (.A(_02098_),
    .B(_02099_),
    .X(_02100_));
 sky130_fd_sc_hd__and2b_1 _09181_ (.A_N(_02100_),
    .B(_02090_),
    .X(_02101_));
 sky130_fd_sc_hd__xnor2_1 _09182_ (.A(_02090_),
    .B(_02100_),
    .Y(_02102_));
 sky130_fd_sc_hd__and2_1 _09183_ (.A(_02089_),
    .B(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__nor2_1 _09184_ (.A(_02089_),
    .B(_02102_),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _09185_ (.A(_02103_),
    .B(_02104_),
    .Y(_02105_));
 sky130_fd_sc_hd__xor2_2 _09186_ (.A(_02036_),
    .B(_02105_),
    .X(_02106_));
 sky130_fd_sc_hd__a32o_1 _09187_ (.A1(_00848_),
    .A2(_00849_),
    .A3(_00863_),
    .B1(_00864_),
    .B2(_00793_),
    .X(_02107_));
 sky130_fd_sc_hd__o21bai_4 _09188_ (.A1(_00774_),
    .A2(_00791_),
    .B1_N(_00790_),
    .Y(_02108_));
 sky130_fd_sc_hd__a21o_2 _09189_ (.A1(_00804_),
    .A2(_00847_),
    .B1(_00846_),
    .X(_02109_));
 sky130_fd_sc_hd__nor2_2 _09190_ (.A(_00859_),
    .B(_00862_),
    .Y(_02110_));
 sky130_fd_sc_hd__o21ai_1 _09191_ (.A1(_00859_),
    .A2(_00862_),
    .B1(_02109_),
    .Y(_02111_));
 sky130_fd_sc_hd__xnor2_4 _09192_ (.A(_02109_),
    .B(_02110_),
    .Y(_02112_));
 sky130_fd_sc_hd__xnor2_2 _09193_ (.A(_02108_),
    .B(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__a21oi_2 _09194_ (.A1(_00867_),
    .A2(_00871_),
    .B1(_00870_),
    .Y(_02114_));
 sky130_fd_sc_hd__xnor2_1 _09195_ (.A(_02113_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__nand2b_1 _09196_ (.A_N(_02115_),
    .B(_02107_),
    .Y(_02116_));
 sky130_fd_sc_hd__xnor2_2 _09197_ (.A(_02107_),
    .B(_02115_),
    .Y(_02117_));
 sky130_fd_sc_hd__xnor2_2 _09198_ (.A(_02106_),
    .B(_02117_),
    .Y(_02118_));
 sky130_fd_sc_hd__and2b_1 _09199_ (.A_N(_02118_),
    .B(_02020_),
    .X(_02119_));
 sky130_fd_sc_hd__xor2_4 _09200_ (.A(_02020_),
    .B(_02118_),
    .X(_02120_));
 sky130_fd_sc_hd__or2_1 _09201_ (.A(_02019_),
    .B(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__and2_1 _09202_ (.A(_02019_),
    .B(_02120_),
    .X(_02122_));
 sky130_fd_sc_hd__xnor2_4 _09203_ (.A(_02019_),
    .B(_02120_),
    .Y(_02123_));
 sky130_fd_sc_hd__a21o_1 _09204_ (.A1(_00881_),
    .A2(_01026_),
    .B1(_00880_),
    .X(_02124_));
 sky130_fd_sc_hd__or2_1 _09205_ (.A(_00882_),
    .B(_01919_),
    .X(_02125_));
 sky130_fd_sc_hd__a211o_1 _09206_ (.A1(_02003_),
    .A2(_02004_),
    .B1(_00882_),
    .C1(_01919_),
    .X(_02126_));
 sky130_fd_sc_hd__o221a_2 _09207_ (.A1(_02011_),
    .A2(_02125_),
    .B1(_02126_),
    .B2(_02012_),
    .C1(_02124_),
    .X(_02127_));
 sky130_fd_sc_hd__xnor2_2 _09208_ (.A(_02123_),
    .B(_02127_),
    .Y(_02128_));
 sky130_fd_sc_hd__a21o_2 _09209_ (.A1(_02106_),
    .A2(_02117_),
    .B1(_02119_),
    .X(_02129_));
 sky130_fd_sc_hd__o21ai_4 _09210_ (.A1(_02113_),
    .A2(_02114_),
    .B1(_02116_),
    .Y(_02130_));
 sky130_fd_sc_hd__o21ai_4 _09211_ (.A1(_02050_),
    .A2(_02073_),
    .B1(_02072_),
    .Y(_02131_));
 sky130_fd_sc_hd__a22o_1 _09212_ (.A1(net30),
    .A2(net112),
    .B1(net107),
    .B2(net14),
    .X(_02132_));
 sky130_fd_sc_hd__xnor2_4 _09213_ (.A(net92),
    .B(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__o22a_1 _09214_ (.A1(net37),
    .A2(_00371_),
    .B1(net110),
    .B2(net39),
    .X(_02134_));
 sky130_fd_sc_hd__xnor2_1 _09215_ (.A(net99),
    .B(_02134_),
    .Y(_02135_));
 sky130_fd_sc_hd__o22a_1 _09216_ (.A1(_00267_),
    .A2(net35),
    .B1(net33),
    .B2(net124),
    .X(_02136_));
 sky130_fd_sc_hd__xnor2_1 _09217_ (.A(net95),
    .B(_02136_),
    .Y(_02137_));
 sky130_fd_sc_hd__nand2_1 _09218_ (.A(_02135_),
    .B(_02137_),
    .Y(_02138_));
 sky130_fd_sc_hd__or2_1 _09219_ (.A(_02135_),
    .B(_02137_),
    .X(_02139_));
 sky130_fd_sc_hd__nand2_2 _09220_ (.A(_02138_),
    .B(_02139_),
    .Y(_02140_));
 sky130_fd_sc_hd__xnor2_4 _09221_ (.A(_02133_),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__o21a_2 _09222_ (.A1(_00856_),
    .A2(_02038_),
    .B1(_02040_),
    .X(_02142_));
 sky130_fd_sc_hd__xnor2_2 _09223_ (.A(_02141_),
    .B(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__and2b_1 _09224_ (.A_N(_02143_),
    .B(_02131_),
    .X(_02144_));
 sky130_fd_sc_hd__xnor2_4 _09225_ (.A(_02131_),
    .B(_02143_),
    .Y(_02145_));
 sky130_fd_sc_hd__a21bo_1 _09226_ (.A1(_02052_),
    .A2(_02054_),
    .B1_N(_02058_),
    .X(_02146_));
 sky130_fd_sc_hd__o21a_1 _09227_ (.A1(_02043_),
    .A2(_02049_),
    .B1(_02048_),
    .X(_02147_));
 sky130_fd_sc_hd__xnor2_2 _09228_ (.A(_02095_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__nand2b_1 _09229_ (.A_N(_02148_),
    .B(_02146_),
    .Y(_02149_));
 sky130_fd_sc_hd__xor2_2 _09230_ (.A(_02146_),
    .B(_02148_),
    .X(_02150_));
 sky130_fd_sc_hd__a22o_1 _09231_ (.A1(_06730_),
    .A2(net129),
    .B1(net127),
    .B2(_00150_),
    .X(_02151_));
 sky130_fd_sc_hd__xnor2_2 _09232_ (.A(net154),
    .B(_02151_),
    .Y(_02152_));
 sky130_fd_sc_hd__o22a_1 _09233_ (.A1(net40),
    .A2(net68),
    .B1(net66),
    .B2(net56),
    .X(_02153_));
 sky130_fd_sc_hd__xnor2_2 _09234_ (.A(net146),
    .B(_02153_),
    .Y(_02154_));
 sky130_fd_sc_hd__o22a_1 _09235_ (.A1(net45),
    .A2(net105),
    .B1(net131),
    .B2(net49),
    .X(_02155_));
 sky130_fd_sc_hd__xnor2_2 _09236_ (.A(net174),
    .B(_02155_),
    .Y(_02156_));
 sky130_fd_sc_hd__nand2_1 _09237_ (.A(_02154_),
    .B(_02156_),
    .Y(_02157_));
 sky130_fd_sc_hd__xnor2_2 _09238_ (.A(_02154_),
    .B(_02156_),
    .Y(_02158_));
 sky130_fd_sc_hd__xnor2_2 _09239_ (.A(_02152_),
    .B(_02158_),
    .Y(_02159_));
 sky130_fd_sc_hd__o22a_1 _09240_ (.A1(net103),
    .A2(net79),
    .B1(net70),
    .B2(net83),
    .X(_02160_));
 sky130_fd_sc_hd__xnor2_1 _09241_ (.A(_00381_),
    .B(_02160_),
    .Y(_02161_));
 sky130_fd_sc_hd__o22a_1 _09242_ (.A1(net24),
    .A2(net76),
    .B1(net74),
    .B2(net23),
    .X(_02162_));
 sky130_fd_sc_hd__xnor2_1 _09243_ (.A(net86),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__o22a_1 _09244_ (.A1(net100),
    .A2(net75),
    .B1(net72),
    .B2(net42),
    .X(_02164_));
 sky130_fd_sc_hd__xnor2_1 _09245_ (.A(net108),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__xnor2_1 _09246_ (.A(_02163_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__or2_1 _09247_ (.A(_02161_),
    .B(_02166_),
    .X(_02167_));
 sky130_fd_sc_hd__nand2_1 _09248_ (.A(_02161_),
    .B(_02166_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _09249_ (.A(_02167_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__a22o_1 _09250_ (.A1(_00158_),
    .A2(_00516_),
    .B1(_00812_),
    .B2(_00159_),
    .X(_02170_));
 sky130_fd_sc_hd__xnor2_4 _09251_ (.A(net200),
    .B(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__o22a_2 _09252_ (.A1(_06701_),
    .A2(net51),
    .B1(net44),
    .B2(_06727_),
    .X(_02172_));
 sky130_fd_sc_hd__xnor2_4 _09253_ (.A(net179),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__or4_2 _09254_ (.A(_05069_),
    .B(_05123_),
    .C(_05221_),
    .D(_00174_),
    .X(_02174_));
 sky130_fd_sc_hd__a21oi_2 _09255_ (.A1(net294),
    .A2(_02174_),
    .B1(_04906_),
    .Y(_02175_));
 sky130_fd_sc_hd__a21o_2 _09256_ (.A1(net294),
    .A2(_02174_),
    .B1(_04906_),
    .X(_02176_));
 sky130_fd_sc_hd__a22o_1 _09257_ (.A1(_00138_),
    .A2(net11),
    .B1(net6),
    .B2(net292),
    .X(_02177_));
 sky130_fd_sc_hd__xnor2_4 _09258_ (.A(net198),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__nand2_1 _09259_ (.A(_02173_),
    .B(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__xnor2_4 _09260_ (.A(_02173_),
    .B(_02178_),
    .Y(_02180_));
 sky130_fd_sc_hd__xor2_4 _09261_ (.A(_02171_),
    .B(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__xnor2_2 _09262_ (.A(_02169_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__and2b_1 _09263_ (.A_N(_02159_),
    .B(_02182_),
    .X(_02183_));
 sky130_fd_sc_hd__xor2_2 _09264_ (.A(_02159_),
    .B(_02182_),
    .X(_02184_));
 sky130_fd_sc_hd__a21oi_1 _09265_ (.A1(net294),
    .A2(_02075_),
    .B1(_04598_),
    .Y(_02185_));
 sky130_fd_sc_hd__a21o_1 _09266_ (.A1(net294),
    .A2(_02075_),
    .B1(_04598_),
    .X(_02186_));
 sky130_fd_sc_hd__a2111o_1 _09267_ (.A1(net294),
    .A2(_00554_),
    .B1(reg1_val[29]),
    .C1(net288),
    .D1(_04598_),
    .X(_02187_));
 sky130_fd_sc_hd__o21ai_2 _09268_ (.A1(_02079_),
    .A2(net61),
    .B1(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__a22o_1 _09269_ (.A1(net153),
    .A2(net9),
    .B1(net4),
    .B2(net207),
    .X(_02189_));
 sky130_fd_sc_hd__xnor2_2 _09270_ (.A(net60),
    .B(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__o21ai_4 _09271_ (.A1(_02061_),
    .A2(_02070_),
    .B1(_02069_),
    .Y(_02191_));
 sky130_fd_sc_hd__a22o_1 _09272_ (.A1(net148),
    .A2(net17),
    .B1(net13),
    .B2(net150),
    .X(_02192_));
 sky130_fd_sc_hd__xnor2_2 _09273_ (.A(net65),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__nand2_1 _09274_ (.A(_02191_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__xor2_2 _09275_ (.A(_02191_),
    .B(_02193_),
    .X(_02195_));
 sky130_fd_sc_hd__xnor2_2 _09276_ (.A(_02190_),
    .B(_02195_),
    .Y(_02196_));
 sky130_fd_sc_hd__or2_1 _09277_ (.A(_02184_),
    .B(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__xnor2_2 _09278_ (.A(_02184_),
    .B(_02196_),
    .Y(_02198_));
 sky130_fd_sc_hd__xor2_1 _09279_ (.A(_02150_),
    .B(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__a21oi_1 _09280_ (.A1(_02025_),
    .A2(_02027_),
    .B1(_02029_),
    .Y(_02200_));
 sky130_fd_sc_hd__o22a_1 _09281_ (.A1(net120),
    .A2(net21),
    .B1(net19),
    .B2(net115),
    .X(_02201_));
 sky130_fd_sc_hd__xnor2_1 _09282_ (.A(net96),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__o22a_1 _09283_ (.A1(net28),
    .A2(net85),
    .B1(net82),
    .B2(net26),
    .X(_02203_));
 sky130_fd_sc_hd__xnor2_1 _09284_ (.A(net90),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__nand2_1 _09285_ (.A(_02202_),
    .B(_02204_),
    .Y(_02205_));
 sky130_fd_sc_hd__or2_1 _09286_ (.A(_02202_),
    .B(_02204_),
    .X(_02206_));
 sky130_fd_sc_hd__nand2_1 _09287_ (.A(_02205_),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__and2_1 _09288_ (.A(_02081_),
    .B(net60),
    .X(_02208_));
 sky130_fd_sc_hd__nor3_1 _09289_ (.A(_02084_),
    .B(_02207_),
    .C(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__o21a_1 _09290_ (.A1(_02084_),
    .A2(_02208_),
    .B1(_02207_),
    .X(_02210_));
 sky130_fd_sc_hd__nor2_1 _09291_ (.A(_02209_),
    .B(_02210_),
    .Y(_02211_));
 sky130_fd_sc_hd__and2b_1 _09292_ (.A_N(_02200_),
    .B(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__xnor2_1 _09293_ (.A(_02200_),
    .B(_02211_),
    .Y(_02213_));
 sky130_fd_sc_hd__and2_1 _09294_ (.A(_02199_),
    .B(_02213_),
    .X(_02214_));
 sky130_fd_sc_hd__nor2_1 _09295_ (.A(_02199_),
    .B(_02213_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_2 _09296_ (.A(_02214_),
    .B(_02215_),
    .Y(_02216_));
 sky130_fd_sc_hd__xor2_4 _09297_ (.A(_02145_),
    .B(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__a21o_2 _09298_ (.A1(_02036_),
    .A2(_02105_),
    .B1(_02103_),
    .X(_02218_));
 sky130_fd_sc_hd__or2_4 _09299_ (.A(_02032_),
    .B(_02035_),
    .X(_02219_));
 sky130_fd_sc_hd__a21o_2 _09300_ (.A1(_02041_),
    .A2(_02088_),
    .B1(_02087_),
    .X(_02220_));
 sky130_fd_sc_hd__nor2_2 _09301_ (.A(_02098_),
    .B(_02101_),
    .Y(_02221_));
 sky130_fd_sc_hd__o21ai_1 _09302_ (.A1(_02098_),
    .A2(_02101_),
    .B1(_02220_),
    .Y(_02222_));
 sky130_fd_sc_hd__xnor2_4 _09303_ (.A(_02220_),
    .B(_02221_),
    .Y(_02223_));
 sky130_fd_sc_hd__xnor2_4 _09304_ (.A(_02219_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__a21boi_4 _09305_ (.A1(_02108_),
    .A2(_02112_),
    .B1_N(_02111_),
    .Y(_02225_));
 sky130_fd_sc_hd__xnor2_4 _09306_ (.A(_02224_),
    .B(_02225_),
    .Y(_02226_));
 sky130_fd_sc_hd__nand2b_1 _09307_ (.A_N(_02226_),
    .B(_02218_),
    .Y(_02227_));
 sky130_fd_sc_hd__xnor2_4 _09308_ (.A(_02218_),
    .B(_02226_),
    .Y(_02228_));
 sky130_fd_sc_hd__and2_1 _09309_ (.A(_02217_),
    .B(_02228_),
    .X(_02229_));
 sky130_fd_sc_hd__xor2_4 _09310_ (.A(_02217_),
    .B(_02228_),
    .X(_02230_));
 sky130_fd_sc_hd__xor2_4 _09311_ (.A(_02130_),
    .B(_02230_),
    .X(_02231_));
 sky130_fd_sc_hd__nor2_1 _09312_ (.A(_02129_),
    .B(_02231_),
    .Y(_02232_));
 sky130_fd_sc_hd__xnor2_4 _09313_ (.A(_02129_),
    .B(_02231_),
    .Y(_02233_));
 sky130_fd_sc_hd__a21oi_2 _09314_ (.A1(_00881_),
    .A2(_02121_),
    .B1(_02122_),
    .Y(_02234_));
 sky130_fd_sc_hd__a21o_1 _09315_ (.A1(_00881_),
    .A2(_02121_),
    .B1(_02122_),
    .X(_02235_));
 sky130_fd_sc_hd__or2_1 _09316_ (.A(_00882_),
    .B(_02123_),
    .X(_02236_));
 sky130_fd_sc_hd__a2111oi_2 _09317_ (.A1(_01025_),
    .A2(_01026_),
    .B1(_02123_),
    .C1(_00955_),
    .D1(_00882_),
    .Y(_02237_));
 sky130_fd_sc_hd__nor4_1 _09318_ (.A(_00882_),
    .B(_01917_),
    .C(_01919_),
    .D(_02123_),
    .Y(_02238_));
 sky130_fd_sc_hd__a211oi_4 _09319_ (.A1(_01915_),
    .A2(_02238_),
    .B1(_02237_),
    .C1(_02234_),
    .Y(_02239_));
 sky130_fd_sc_hd__xor2_2 _09320_ (.A(_02233_),
    .B(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__or4b_4 _09321_ (.A(_01922_),
    .B(_02240_),
    .C(_02017_),
    .D_N(_02128_),
    .X(_02241_));
 sky130_fd_sc_hd__a2111o_1 _09322_ (.A1(_02011_),
    .A2(_02013_),
    .B1(_02123_),
    .C1(_02125_),
    .D1(_02233_),
    .X(_02242_));
 sky130_fd_sc_hd__a21boi_1 _09323_ (.A1(_02129_),
    .A2(_02231_),
    .B1_N(_02121_),
    .Y(_02243_));
 sky130_fd_sc_hd__o32a_1 _09324_ (.A1(_02123_),
    .A2(_02124_),
    .A3(_02233_),
    .B1(_02243_),
    .B2(_02232_),
    .X(_02244_));
 sky130_fd_sc_hd__nand2_1 _09325_ (.A(_02242_),
    .B(_02244_),
    .Y(_02245_));
 sky130_fd_sc_hd__a21oi_4 _09326_ (.A1(_02130_),
    .A2(_02230_),
    .B1(_02229_),
    .Y(_02246_));
 sky130_fd_sc_hd__o21ai_4 _09327_ (.A1(_02224_),
    .A2(_02225_),
    .B1(_02227_),
    .Y(_02247_));
 sky130_fd_sc_hd__a31o_2 _09328_ (.A1(_02167_),
    .A2(_02168_),
    .A3(_02181_),
    .B1(_02183_),
    .X(_02248_));
 sky130_fd_sc_hd__o22a_1 _09329_ (.A1(_00286_),
    .A2(net35),
    .B1(net33),
    .B2(_00477_),
    .X(_02249_));
 sky130_fd_sc_hd__xnor2_1 _09330_ (.A(net95),
    .B(_02249_),
    .Y(_02250_));
 sky130_fd_sc_hd__inv_2 _09331_ (.A(_02250_),
    .Y(_02251_));
 sky130_fd_sc_hd__a22o_1 _09332_ (.A1(_00266_),
    .A2(net17),
    .B1(net13),
    .B2(net148),
    .X(_02252_));
 sky130_fd_sc_hd__xnor2_2 _09333_ (.A(net65),
    .B(_02252_),
    .Y(_02253_));
 sky130_fd_sc_hd__a22o_1 _09334_ (.A1(net14),
    .A2(net112),
    .B1(net111),
    .B2(net30),
    .X(_02254_));
 sky130_fd_sc_hd__xnor2_2 _09335_ (.A(net91),
    .B(_02254_),
    .Y(_02255_));
 sky130_fd_sc_hd__nand2_1 _09336_ (.A(_02253_),
    .B(_02255_),
    .Y(_02256_));
 sky130_fd_sc_hd__xnor2_2 _09337_ (.A(_02253_),
    .B(_02255_),
    .Y(_02257_));
 sky130_fd_sc_hd__xnor2_2 _09338_ (.A(_02251_),
    .B(_02257_),
    .Y(_02258_));
 sky130_fd_sc_hd__o21a_1 _09339_ (.A1(_02095_),
    .A2(_02147_),
    .B1(_02149_),
    .X(_02259_));
 sky130_fd_sc_hd__xnor2_2 _09340_ (.A(_02258_),
    .B(_02259_),
    .Y(_02260_));
 sky130_fd_sc_hd__and2b_1 _09341_ (.A_N(_02260_),
    .B(_02248_),
    .X(_02261_));
 sky130_fd_sc_hd__xnor2_4 _09342_ (.A(_02248_),
    .B(_02260_),
    .Y(_02262_));
 sky130_fd_sc_hd__a21bo_1 _09343_ (.A1(_02163_),
    .A2(_02165_),
    .B1_N(_02167_),
    .X(_02263_));
 sky130_fd_sc_hd__o21a_1 _09344_ (.A1(_02152_),
    .A2(_02158_),
    .B1(_02157_),
    .X(_02264_));
 sky130_fd_sc_hd__or2_1 _09345_ (.A(_02205_),
    .B(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__xnor2_1 _09346_ (.A(_02205_),
    .B(_02264_),
    .Y(_02266_));
 sky130_fd_sc_hd__nand2b_1 _09347_ (.A_N(_02266_),
    .B(_02263_),
    .Y(_02267_));
 sky130_fd_sc_hd__nand2b_1 _09348_ (.A_N(_02263_),
    .B(_02266_),
    .Y(_02268_));
 sky130_fd_sc_hd__nand2_1 _09349_ (.A(_02267_),
    .B(_02268_),
    .Y(_02269_));
 sky130_fd_sc_hd__a22o_1 _09350_ (.A1(_00150_),
    .A2(net129),
    .B1(net127),
    .B2(_00161_),
    .X(_02270_));
 sky130_fd_sc_hd__xnor2_2 _09351_ (.A(net154),
    .B(_02270_),
    .Y(_02271_));
 sky130_fd_sc_hd__o22a_1 _09352_ (.A1(net49),
    .A2(net105),
    .B1(net131),
    .B2(net51),
    .X(_02272_));
 sky130_fd_sc_hd__xnor2_1 _09353_ (.A(net174),
    .B(_02272_),
    .Y(_02273_));
 sky130_fd_sc_hd__o22a_1 _09354_ (.A1(net56),
    .A2(net68),
    .B1(net66),
    .B2(net53),
    .X(_02274_));
 sky130_fd_sc_hd__xnor2_1 _09355_ (.A(net146),
    .B(_02274_),
    .Y(_02275_));
 sky130_fd_sc_hd__nand2_1 _09356_ (.A(_02273_),
    .B(_02275_),
    .Y(_02276_));
 sky130_fd_sc_hd__or2_1 _09357_ (.A(_02273_),
    .B(_02275_),
    .X(_02277_));
 sky130_fd_sc_hd__nand2_1 _09358_ (.A(_02276_),
    .B(_02277_),
    .Y(_02278_));
 sky130_fd_sc_hd__xnor2_2 _09359_ (.A(_02271_),
    .B(_02278_),
    .Y(_02279_));
 sky130_fd_sc_hd__o22a_1 _09360_ (.A1(net103),
    .A2(net83),
    .B1(net79),
    .B2(net100),
    .X(_02280_));
 sky130_fd_sc_hd__xnor2_1 _09361_ (.A(net116),
    .B(_02280_),
    .Y(_02281_));
 sky130_fd_sc_hd__o22a_1 _09362_ (.A1(net25),
    .A2(net74),
    .B1(net70),
    .B2(net23),
    .X(_02282_));
 sky130_fd_sc_hd__xnor2_1 _09363_ (.A(net86),
    .B(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__o22a_1 _09364_ (.A1(net42),
    .A2(net75),
    .B1(net72),
    .B2(net40),
    .X(_02284_));
 sky130_fd_sc_hd__xnor2_1 _09365_ (.A(net108),
    .B(_02284_),
    .Y(_02285_));
 sky130_fd_sc_hd__and2_1 _09366_ (.A(_02283_),
    .B(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__nor2_1 _09367_ (.A(_02283_),
    .B(_02285_),
    .Y(_02287_));
 sky130_fd_sc_hd__nor2_1 _09368_ (.A(_02286_),
    .B(_02287_),
    .Y(_02288_));
 sky130_fd_sc_hd__xnor2_1 _09369_ (.A(_02281_),
    .B(_02288_),
    .Y(_02289_));
 sky130_fd_sc_hd__a22o_1 _09370_ (.A1(_00158_),
    .A2(_00812_),
    .B1(net11),
    .B2(_00159_),
    .X(_02290_));
 sky130_fd_sc_hd__xnor2_2 _09371_ (.A(net200),
    .B(_02290_),
    .Y(_02291_));
 sky130_fd_sc_hd__o32a_1 _09372_ (.A1(_06727_),
    .A2(_00513_),
    .A3(_00515_),
    .B1(net44),
    .B2(_06701_),
    .X(_02292_));
 sky130_fd_sc_hd__xnor2_2 _09373_ (.A(net180),
    .B(_02292_),
    .Y(_02293_));
 sky130_fd_sc_hd__a21oi_2 _09374_ (.A1(_00138_),
    .A2(net6),
    .B1(net198),
    .Y(_02294_));
 sky130_fd_sc_hd__nand2_1 _09375_ (.A(_02293_),
    .B(_02294_),
    .Y(_02295_));
 sky130_fd_sc_hd__xnor2_2 _09376_ (.A(_02293_),
    .B(_02294_),
    .Y(_02296_));
 sky130_fd_sc_hd__xor2_2 _09377_ (.A(_02291_),
    .B(_02296_),
    .X(_02297_));
 sky130_fd_sc_hd__and2b_1 _09378_ (.A_N(_02289_),
    .B(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__xor2_1 _09379_ (.A(_02289_),
    .B(_02297_),
    .X(_02299_));
 sky130_fd_sc_hd__xor2_1 _09380_ (.A(_02279_),
    .B(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__nor2_1 _09381_ (.A(net212),
    .B(net60),
    .Y(_02301_));
 sky130_fd_sc_hd__o21a_1 _09382_ (.A1(_02171_),
    .A2(_02180_),
    .B1(_02179_),
    .X(_02302_));
 sky130_fd_sc_hd__a22o_1 _09383_ (.A1(net150),
    .A2(net9),
    .B1(net4),
    .B2(net153),
    .X(_02303_));
 sky130_fd_sc_hd__xnor2_1 _09384_ (.A(net60),
    .B(_02303_),
    .Y(_02304_));
 sky130_fd_sc_hd__and2b_1 _09385_ (.A_N(_02302_),
    .B(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__xnor2_1 _09386_ (.A(_02302_),
    .B(_02304_),
    .Y(_02306_));
 sky130_fd_sc_hd__xor2_1 _09387_ (.A(_02301_),
    .B(_02306_),
    .X(_02307_));
 sky130_fd_sc_hd__nand2_1 _09388_ (.A(_02300_),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__xnor2_1 _09389_ (.A(_02300_),
    .B(_02307_),
    .Y(_02309_));
 sky130_fd_sc_hd__xor2_1 _09390_ (.A(_02269_),
    .B(_02309_),
    .X(_02310_));
 sky130_fd_sc_hd__o21ai_2 _09391_ (.A1(_02133_),
    .A2(_02140_),
    .B1(_02138_),
    .Y(_02311_));
 sky130_fd_sc_hd__inv_2 _09392_ (.A(_02311_),
    .Y(_02312_));
 sky130_fd_sc_hd__o22a_1 _09393_ (.A1(_00391_),
    .A2(net21),
    .B1(net19),
    .B2(net85),
    .X(_02313_));
 sky130_fd_sc_hd__xnor2_1 _09394_ (.A(net97),
    .B(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__inv_2 _09395_ (.A(_02314_),
    .Y(_02315_));
 sky130_fd_sc_hd__o22a_1 _09396_ (.A1(net28),
    .A2(_00442_),
    .B1(net76),
    .B2(net27),
    .X(_02316_));
 sky130_fd_sc_hd__xnor2_1 _09397_ (.A(net88),
    .B(_02316_),
    .Y(_02317_));
 sky130_fd_sc_hd__o22a_1 _09398_ (.A1(net39),
    .A2(_00371_),
    .B1(net120),
    .B2(net37),
    .X(_02318_));
 sky130_fd_sc_hd__xnor2_1 _09399_ (.A(net99),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__nand2_1 _09400_ (.A(_02317_),
    .B(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__xnor2_1 _09401_ (.A(_02317_),
    .B(_02319_),
    .Y(_02321_));
 sky130_fd_sc_hd__xnor2_1 _09402_ (.A(_02315_),
    .B(_02321_),
    .Y(_02322_));
 sky130_fd_sc_hd__a21boi_2 _09403_ (.A1(_02190_),
    .A2(_02195_),
    .B1_N(_02194_),
    .Y(_02323_));
 sky130_fd_sc_hd__nor2_1 _09404_ (.A(_02322_),
    .B(_02323_),
    .Y(_02324_));
 sky130_fd_sc_hd__xnor2_1 _09405_ (.A(_02322_),
    .B(_02323_),
    .Y(_02325_));
 sky130_fd_sc_hd__xnor2_1 _09406_ (.A(_02311_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__and2_1 _09407_ (.A(_02310_),
    .B(_02326_),
    .X(_02327_));
 sky130_fd_sc_hd__nor2_1 _09408_ (.A(_02310_),
    .B(_02326_),
    .Y(_02328_));
 sky130_fd_sc_hd__nor2_2 _09409_ (.A(_02327_),
    .B(_02328_),
    .Y(_02329_));
 sky130_fd_sc_hd__xor2_4 _09410_ (.A(_02262_),
    .B(_02329_),
    .X(_02330_));
 sky130_fd_sc_hd__a21o_1 _09411_ (.A1(_02145_),
    .A2(_02216_),
    .B1(_02214_),
    .X(_02331_));
 sky130_fd_sc_hd__o21bai_4 _09412_ (.A1(_02141_),
    .A2(_02142_),
    .B1_N(_02144_),
    .Y(_02332_));
 sky130_fd_sc_hd__o21ai_4 _09413_ (.A1(_02150_),
    .A2(_02198_),
    .B1(_02197_),
    .Y(_02333_));
 sky130_fd_sc_hd__nor2_2 _09414_ (.A(_02209_),
    .B(_02212_),
    .Y(_02334_));
 sky130_fd_sc_hd__o21a_1 _09415_ (.A1(_02209_),
    .A2(_02212_),
    .B1(_02333_),
    .X(_02335_));
 sky130_fd_sc_hd__xnor2_4 _09416_ (.A(_02333_),
    .B(_02334_),
    .Y(_02336_));
 sky130_fd_sc_hd__xnor2_4 _09417_ (.A(_02332_),
    .B(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__a21boi_4 _09418_ (.A1(_02219_),
    .A2(_02223_),
    .B1_N(_02222_),
    .Y(_02338_));
 sky130_fd_sc_hd__xnor2_2 _09419_ (.A(_02337_),
    .B(_02338_),
    .Y(_02339_));
 sky130_fd_sc_hd__nand2b_1 _09420_ (.A_N(_02339_),
    .B(_02331_),
    .Y(_02340_));
 sky130_fd_sc_hd__xnor2_2 _09421_ (.A(_02331_),
    .B(_02339_),
    .Y(_02341_));
 sky130_fd_sc_hd__and2_1 _09422_ (.A(_02330_),
    .B(_02341_),
    .X(_02342_));
 sky130_fd_sc_hd__xor2_4 _09423_ (.A(_02330_),
    .B(_02341_),
    .X(_02343_));
 sky130_fd_sc_hd__xnor2_4 _09424_ (.A(_02247_),
    .B(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__and2_1 _09425_ (.A(_02246_),
    .B(_02344_),
    .X(_02345_));
 sky130_fd_sc_hd__xnor2_4 _09426_ (.A(_02246_),
    .B(_02344_),
    .Y(_02346_));
 sky130_fd_sc_hd__xnor2_2 _09427_ (.A(_02245_),
    .B(_02346_),
    .Y(_02347_));
 sky130_fd_sc_hd__and4b_4 _09428_ (.A_N(net298),
    .B(net297),
    .C(_04434_),
    .D(instruction[3]),
    .X(_02348_));
 sky130_fd_sc_hd__or4b_4 _09429_ (.A(_04423_),
    .B(net298),
    .C(instruction[5]),
    .D_N(net297),
    .X(_02349_));
 sky130_fd_sc_hd__a21oi_1 _09430_ (.A1(net138),
    .A2(_02241_),
    .B1(_02347_),
    .Y(_02350_));
 sky130_fd_sc_hd__a31o_1 _09431_ (.A1(net138),
    .A2(_02241_),
    .A3(_02347_),
    .B1(net235),
    .X(_02351_));
 sky130_fd_sc_hd__or2_1 _09432_ (.A(_02350_),
    .B(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__or4b_2 _09433_ (.A(instruction[3]),
    .B(net298),
    .C(_06676_),
    .D_N(_06634_),
    .X(_02353_));
 sky130_fd_sc_hd__nor2_1 _09434_ (.A(net284),
    .B(_06670_),
    .Y(_02354_));
 sky130_fd_sc_hd__or2_1 _09435_ (.A(net284),
    .B(_06670_),
    .X(_02355_));
 sky130_fd_sc_hd__mux2_1 _09436_ (.A0(net289),
    .A1(net288),
    .S(net170),
    .X(_02356_));
 sky130_fd_sc_hd__mux2_1 _09437_ (.A0(net285),
    .A1(_04598_),
    .S(net170),
    .X(_02357_));
 sky130_fd_sc_hd__nand2_1 _09438_ (.A(net210),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__o211a_1 _09439_ (.A1(net210),
    .A2(_02356_),
    .B1(_02358_),
    .C1(net213),
    .X(_02359_));
 sky130_fd_sc_hd__mux2_1 _09440_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net170),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _09441_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net170),
    .X(_02361_));
 sky130_fd_sc_hd__mux2_1 _09442_ (.A0(_02360_),
    .A1(_02361_),
    .S(net210),
    .X(_02362_));
 sky130_fd_sc_hd__mux2_1 _09443_ (.A0(net287),
    .A1(reg1_val[24]),
    .S(net170),
    .X(_02363_));
 sky130_fd_sc_hd__mux2_1 _09444_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net170),
    .X(_02364_));
 sky130_fd_sc_hd__mux2_1 _09445_ (.A0(_02363_),
    .A1(_02364_),
    .S(net208),
    .X(_02365_));
 sky130_fd_sc_hd__mux2_1 _09446_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net170),
    .X(_02366_));
 sky130_fd_sc_hd__mux2_1 _09447_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net170),
    .X(_02367_));
 sky130_fd_sc_hd__mux2_1 _09448_ (.A0(_02366_),
    .A1(_02367_),
    .S(net208),
    .X(_02368_));
 sky130_fd_sc_hd__mux2_1 _09449_ (.A0(_02365_),
    .A1(_02368_),
    .S(net213),
    .X(_02369_));
 sky130_fd_sc_hd__a211o_1 _09450_ (.A1(_06569_),
    .A2(_02362_),
    .B1(_02359_),
    .C1(net216),
    .X(_02370_));
 sky130_fd_sc_hd__o211a_1 _09451_ (.A1(net217),
    .A2(_02369_),
    .B1(_02370_),
    .C1(_06553_),
    .X(_02371_));
 sky130_fd_sc_hd__mux2_1 _09452_ (.A0(reg1_val[15]),
    .A1(reg1_val[16]),
    .S(net170),
    .X(_02372_));
 sky130_fd_sc_hd__mux2_1 _09453_ (.A0(reg1_val[14]),
    .A1(reg1_val[17]),
    .S(net170),
    .X(_02373_));
 sky130_fd_sc_hd__mux2_1 _09454_ (.A0(_02372_),
    .A1(_02373_),
    .S(net210),
    .X(_02374_));
 sky130_fd_sc_hd__mux2_1 _09455_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net170),
    .X(_02375_));
 sky130_fd_sc_hd__mux2_1 _09456_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net170),
    .X(_02376_));
 sky130_fd_sc_hd__mux2_1 _09457_ (.A0(_02375_),
    .A1(_02376_),
    .S(net208),
    .X(_02377_));
 sky130_fd_sc_hd__mux2_1 _09458_ (.A0(_02374_),
    .A1(_02377_),
    .S(net213),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _09459_ (.A0(net290),
    .A1(reg1_val[20]),
    .S(net170),
    .X(_02379_));
 sky130_fd_sc_hd__mux2_1 _09460_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net170),
    .X(_02380_));
 sky130_fd_sc_hd__mux2_1 _09461_ (.A0(_02379_),
    .A1(_02380_),
    .S(net208),
    .X(_02381_));
 sky130_fd_sc_hd__mux2_1 _09462_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net170),
    .X(_02382_));
 sky130_fd_sc_hd__mux2_1 _09463_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net170),
    .X(_02383_));
 sky130_fd_sc_hd__mux2_1 _09464_ (.A0(_02382_),
    .A1(_02383_),
    .S(net208),
    .X(_02384_));
 sky130_fd_sc_hd__mux2_1 _09465_ (.A0(_02381_),
    .A1(_02384_),
    .S(net213),
    .X(_02385_));
 sky130_fd_sc_hd__mux2_1 _09466_ (.A0(_02378_),
    .A1(_02385_),
    .S(net217),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _09467_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net168),
    .X(_02387_));
 sky130_fd_sc_hd__mux2_1 _09468_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net168),
    .X(_02388_));
 sky130_fd_sc_hd__mux2_1 _09469_ (.A0(_02387_),
    .A1(_02388_),
    .S(net210),
    .X(_02389_));
 sky130_fd_sc_hd__mux2_1 _09470_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net168),
    .X(_02390_));
 sky130_fd_sc_hd__mux2_1 _09471_ (.A0(net290),
    .A1(reg1_val[20]),
    .S(net168),
    .X(_02391_));
 sky130_fd_sc_hd__mux2_1 _09472_ (.A0(_02390_),
    .A1(_02391_),
    .S(net210),
    .X(_02392_));
 sky130_fd_sc_hd__mux2_1 _09473_ (.A0(_02389_),
    .A1(_02392_),
    .S(net213),
    .X(_02393_));
 sky130_fd_sc_hd__mux2_1 _09474_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net168),
    .X(_02394_));
 sky130_fd_sc_hd__mux2_1 _09475_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net168),
    .X(_02395_));
 sky130_fd_sc_hd__mux2_1 _09476_ (.A0(_02394_),
    .A1(_02395_),
    .S(net210),
    .X(_02396_));
 sky130_fd_sc_hd__mux2_1 _09477_ (.A0(reg1_val[14]),
    .A1(reg1_val[17]),
    .S(net168),
    .X(_02397_));
 sky130_fd_sc_hd__mux2_1 _09478_ (.A0(reg1_val[15]),
    .A1(reg1_val[16]),
    .S(net168),
    .X(_02398_));
 sky130_fd_sc_hd__mux2_1 _09479_ (.A0(_02397_),
    .A1(_02398_),
    .S(net210),
    .X(_02399_));
 sky130_fd_sc_hd__mux2_1 _09480_ (.A0(_02396_),
    .A1(_02399_),
    .S(net213),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _09481_ (.A0(_02393_),
    .A1(_02400_),
    .S(net217),
    .X(_02401_));
 sky130_fd_sc_hd__mux2_1 _09482_ (.A0(net291),
    .A1(reg1_val[31]),
    .S(net169),
    .X(_02402_));
 sky130_fd_sc_hd__mux2_1 _09483_ (.A0(net289),
    .A1(net288),
    .S(net169),
    .X(_02403_));
 sky130_fd_sc_hd__mux2_1 _09484_ (.A0(_02402_),
    .A1(_02403_),
    .S(net211),
    .X(_02404_));
 sky130_fd_sc_hd__mux2_1 _09485_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net169),
    .X(_02405_));
 sky130_fd_sc_hd__mux2_1 _09486_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net168),
    .X(_02406_));
 sky130_fd_sc_hd__mux2_1 _09487_ (.A0(_02405_),
    .A1(_02406_),
    .S(net210),
    .X(_02407_));
 sky130_fd_sc_hd__mux2_1 _09488_ (.A0(_02404_),
    .A1(_02407_),
    .S(net214),
    .X(_02408_));
 sky130_fd_sc_hd__mux2_1 _09489_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net168),
    .X(_02409_));
 sky130_fd_sc_hd__mux2_1 _09490_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net168),
    .X(_02410_));
 sky130_fd_sc_hd__mux2_1 _09491_ (.A0(_02409_),
    .A1(_02410_),
    .S(net210),
    .X(_02411_));
 sky130_fd_sc_hd__mux2_1 _09492_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net168),
    .X(_02412_));
 sky130_fd_sc_hd__mux2_1 _09493_ (.A0(net287),
    .A1(reg1_val[24]),
    .S(net168),
    .X(_02413_));
 sky130_fd_sc_hd__mux2_1 _09494_ (.A0(_02412_),
    .A1(_02413_),
    .S(net210),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _09495_ (.A0(_02411_),
    .A1(_02414_),
    .S(net214),
    .X(_02415_));
 sky130_fd_sc_hd__mux2_1 _09496_ (.A0(_02408_),
    .A1(_02415_),
    .S(_06560_),
    .X(_02416_));
 sky130_fd_sc_hd__mux2_1 _09497_ (.A0(_02401_),
    .A1(_02416_),
    .S(net218),
    .X(_02417_));
 sky130_fd_sc_hd__a211o_1 _09498_ (.A1(net219),
    .A2(_02386_),
    .B1(_02371_),
    .C1(net222),
    .X(_02418_));
 sky130_fd_sc_hd__o21ai_2 _09499_ (.A1(net220),
    .A2(_02417_),
    .B1(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__nand2_1 _09500_ (.A(net291),
    .B(curr_PC[0]),
    .Y(_02420_));
 sky130_fd_sc_hd__or2_1 _09501_ (.A(net291),
    .B(curr_PC[0]),
    .X(_02421_));
 sky130_fd_sc_hd__a21oi_1 _09502_ (.A1(_02420_),
    .A2(_02421_),
    .B1(net223),
    .Y(_02422_));
 sky130_fd_sc_hd__a211o_1 _09503_ (.A1(net223),
    .A2(_02419_),
    .B1(_02422_),
    .C1(_06667_),
    .X(_02423_));
 sky130_fd_sc_hd__nor2_2 _09504_ (.A(net295),
    .B(_06670_),
    .Y(_02424_));
 sky130_fd_sc_hd__or2_4 _09505_ (.A(net295),
    .B(_06670_),
    .X(_02425_));
 sky130_fd_sc_hd__and3b_4 _09506_ (.A_N(net297),
    .B(_04434_),
    .C(_06636_),
    .X(_02426_));
 sky130_fd_sc_hd__or3_4 _09507_ (.A(instruction[3]),
    .B(net298),
    .C(_06668_),
    .X(_02427_));
 sky130_fd_sc_hd__nor2_1 _09508_ (.A(_06650_),
    .B(_06676_),
    .Y(_02428_));
 sky130_fd_sc_hd__or2_4 _09509_ (.A(_06650_),
    .B(_06676_),
    .X(_02429_));
 sky130_fd_sc_hd__a21o_1 _09510_ (.A1(_02427_),
    .A2(_02429_),
    .B1(_06639_),
    .X(_02430_));
 sky130_fd_sc_hd__and4b_1 _09511_ (.A_N(net298),
    .B(net297),
    .C(instruction[5]),
    .D(instruction[3]),
    .X(_02431_));
 sky130_fd_sc_hd__or4b_4 _09512_ (.A(_04423_),
    .B(_04434_),
    .C(instruction[4]),
    .D_N(net297),
    .X(_02432_));
 sky130_fd_sc_hd__and3_2 _09513_ (.A(net297),
    .B(_04434_),
    .C(_06636_),
    .X(_02433_));
 sky130_fd_sc_hd__nand2_8 _09514_ (.A(_06636_),
    .B(_06656_),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_4 _09515_ (.A(_04434_),
    .B(_06665_),
    .Y(_02435_));
 sky130_fd_sc_hd__or2_2 _09516_ (.A(_04434_),
    .B(_06665_),
    .X(_02436_));
 sky130_fd_sc_hd__a21o_1 _09517_ (.A1(_02434_),
    .A2(net194),
    .B1(net211),
    .X(_02437_));
 sky130_fd_sc_hd__a21o_1 _09518_ (.A1(_02432_),
    .A2(_02437_),
    .B1(net285),
    .X(_02438_));
 sky130_fd_sc_hd__nor2_2 _09519_ (.A(_06669_),
    .B(_06676_),
    .Y(_02439_));
 sky130_fd_sc_hd__or2_4 _09520_ (.A(_06669_),
    .B(_06676_),
    .X(_02440_));
 sky130_fd_sc_hd__nor2_4 _09521_ (.A(_04423_),
    .B(_06658_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_1 _09522_ (.A(instruction[3]),
    .B(_06657_),
    .Y(_02442_));
 sky130_fd_sc_hd__nor2_4 _09523_ (.A(instruction[3]),
    .B(_06658_),
    .Y(_02443_));
 sky130_fd_sc_hd__nand2_1 _09524_ (.A(_04423_),
    .B(_06657_),
    .Y(_02444_));
 sky130_fd_sc_hd__nand3_2 _09525_ (.A(net297),
    .B(instruction[5]),
    .C(_06636_),
    .Y(_02445_));
 sky130_fd_sc_hd__a2bb2o_1 _09526_ (.A1_N(net291),
    .A2_N(net232),
    .B1(_02441_),
    .B2(\div_shifter[32] ),
    .X(_02446_));
 sky130_fd_sc_hd__a221o_1 _09527_ (.A1(_06638_),
    .A2(net193),
    .B1(_02443_),
    .B2(\div_res[0] ),
    .C1(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__and3b_1 _09528_ (.A_N(_02447_),
    .B(_02438_),
    .C(_02430_),
    .X(_02448_));
 sky130_fd_sc_hd__nor2_2 _09529_ (.A(_04598_),
    .B(_06667_),
    .Y(_02449_));
 sky130_fd_sc_hd__mux2_1 _09530_ (.A0(_02402_),
    .A1(_02449_),
    .S(net206),
    .X(_02450_));
 sky130_fd_sc_hd__o21a_1 _09531_ (.A1(net214),
    .A2(_02449_),
    .B1(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__or2_1 _09532_ (.A(net217),
    .B(_02449_),
    .X(_02452_));
 sky130_fd_sc_hd__or2_4 _09533_ (.A(_06553_),
    .B(_02449_),
    .X(_02453_));
 sky130_fd_sc_hd__and3_1 _09534_ (.A(_02451_),
    .B(_02452_),
    .C(_02453_),
    .X(_02454_));
 sky130_fd_sc_hd__nor2_2 _09535_ (.A(net220),
    .B(_02449_),
    .Y(_02455_));
 sky130_fd_sc_hd__or2_4 _09536_ (.A(net220),
    .B(_02449_),
    .X(_02456_));
 sky130_fd_sc_hd__nand2_2 _09537_ (.A(_02454_),
    .B(_02456_),
    .Y(_02457_));
 sky130_fd_sc_hd__o221a_1 _09538_ (.A1(_02419_),
    .A2(_02425_),
    .B1(_02457_),
    .B2(net169),
    .C1(_02448_),
    .X(_02458_));
 sky130_fd_sc_hd__o311a_1 _09539_ (.A1(instruction[5]),
    .A2(_06623_),
    .A3(_06650_),
    .B1(_02423_),
    .C1(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__a31o_1 _09540_ (.A1(_02352_),
    .A2(_02353_),
    .A3(_02459_),
    .B1(_06679_),
    .X(_02460_));
 sky130_fd_sc_hd__o21a_1 _09541_ (.A1(net211),
    .A2(net203),
    .B1(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__or2_1 _09542_ (.A(curr_PC[0]),
    .B(net237),
    .X(_02462_));
 sky130_fd_sc_hd__o21ai_4 _09543_ (.A1(net242),
    .A2(_02461_),
    .B1(_02462_),
    .Y(dest_val[0]));
 sky130_fd_sc_hd__nor2_1 _09544_ (.A(_02241_),
    .B(_02347_),
    .Y(_02463_));
 sky130_fd_sc_hd__a21oi_4 _09545_ (.A1(_02247_),
    .A2(_02343_),
    .B1(_02342_),
    .Y(_02464_));
 sky130_fd_sc_hd__o21ai_4 _09546_ (.A1(_02337_),
    .A2(_02338_),
    .B1(_02340_),
    .Y(_02465_));
 sky130_fd_sc_hd__o21ba_2 _09547_ (.A1(_02279_),
    .A2(_02299_),
    .B1_N(_02298_),
    .X(_02466_));
 sky130_fd_sc_hd__o22a_1 _09548_ (.A1(net33),
    .A2(net113),
    .B1(_00477_),
    .B2(net35),
    .X(_02467_));
 sky130_fd_sc_hd__xnor2_1 _09549_ (.A(net95),
    .B(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__a22o_1 _09550_ (.A1(_00287_),
    .A2(net17),
    .B1(net13),
    .B2(_00266_),
    .X(_02469_));
 sky130_fd_sc_hd__xnor2_1 _09551_ (.A(net65),
    .B(_02469_),
    .Y(_02470_));
 sky130_fd_sc_hd__a22o_1 _09552_ (.A1(net30),
    .A2(net122),
    .B1(net111),
    .B2(net14),
    .X(_02471_));
 sky130_fd_sc_hd__xnor2_1 _09553_ (.A(net91),
    .B(_02471_),
    .Y(_02472_));
 sky130_fd_sc_hd__nand2_1 _09554_ (.A(_02470_),
    .B(_02472_),
    .Y(_02473_));
 sky130_fd_sc_hd__xnor2_1 _09555_ (.A(_02470_),
    .B(_02472_),
    .Y(_02474_));
 sky130_fd_sc_hd__inv_2 _09556_ (.A(_02474_),
    .Y(_02475_));
 sky130_fd_sc_hd__xor2_1 _09557_ (.A(_02468_),
    .B(_02474_),
    .X(_02476_));
 sky130_fd_sc_hd__a21oi_1 _09558_ (.A1(_02265_),
    .A2(_02267_),
    .B1(_02476_),
    .Y(_02477_));
 sky130_fd_sc_hd__and3_1 _09559_ (.A(_02265_),
    .B(_02267_),
    .C(_02476_),
    .X(_02478_));
 sky130_fd_sc_hd__nor2_2 _09560_ (.A(_02477_),
    .B(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__and2b_1 _09561_ (.A_N(_02466_),
    .B(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__xnor2_4 _09562_ (.A(_02466_),
    .B(_02479_),
    .Y(_02481_));
 sky130_fd_sc_hd__a21o_1 _09563_ (.A1(_02281_),
    .A2(_02288_),
    .B1(_02286_),
    .X(_02482_));
 sky130_fd_sc_hd__o21a_1 _09564_ (.A1(_02315_),
    .A2(_02321_),
    .B1(_02320_),
    .X(_02483_));
 sky130_fd_sc_hd__o21a_1 _09565_ (.A1(_02271_),
    .A2(_02278_),
    .B1(_02276_),
    .X(_02484_));
 sky130_fd_sc_hd__nor2_1 _09566_ (.A(_02483_),
    .B(_02484_),
    .Y(_02485_));
 sky130_fd_sc_hd__xor2_2 _09567_ (.A(_02483_),
    .B(_02484_),
    .X(_02486_));
 sky130_fd_sc_hd__xnor2_1 _09568_ (.A(_02482_),
    .B(_02486_),
    .Y(_02487_));
 sky130_fd_sc_hd__o22a_1 _09569_ (.A1(net45),
    .A2(_00227_),
    .B1(_00232_),
    .B2(net49),
    .X(_02488_));
 sky130_fd_sc_hd__xnor2_1 _09570_ (.A(net154),
    .B(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__inv_2 _09571_ (.A(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__o22a_1 _09572_ (.A1(net51),
    .A2(net105),
    .B1(net131),
    .B2(net44),
    .X(_02491_));
 sky130_fd_sc_hd__xnor2_1 _09573_ (.A(net174),
    .B(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__o22a_1 _09574_ (.A1(net53),
    .A2(net68),
    .B1(net66),
    .B2(net47),
    .X(_02493_));
 sky130_fd_sc_hd__xnor2_1 _09575_ (.A(net146),
    .B(_02493_),
    .Y(_02494_));
 sky130_fd_sc_hd__nand2_1 _09576_ (.A(_02492_),
    .B(_02494_),
    .Y(_02495_));
 sky130_fd_sc_hd__or2_1 _09577_ (.A(_02492_),
    .B(_02494_),
    .X(_02496_));
 sky130_fd_sc_hd__nand2_1 _09578_ (.A(_02495_),
    .B(_02496_),
    .Y(_02497_));
 sky130_fd_sc_hd__xnor2_1 _09579_ (.A(_02489_),
    .B(_02497_),
    .Y(_02498_));
 sky130_fd_sc_hd__a22o_1 _09580_ (.A1(_00158_),
    .A2(net11),
    .B1(net6),
    .B2(_00159_),
    .X(_02499_));
 sky130_fd_sc_hd__xnor2_1 _09581_ (.A(net202),
    .B(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__or3_1 _09582_ (.A(_06701_),
    .B(_00513_),
    .C(_00515_),
    .X(_02501_));
 sky130_fd_sc_hd__a21o_1 _09583_ (.A1(_00809_),
    .A2(_00810_),
    .B1(_06727_),
    .X(_02502_));
 sky130_fd_sc_hd__a21o_1 _09584_ (.A1(_02501_),
    .A2(_02502_),
    .B1(net181),
    .X(_02503_));
 sky130_fd_sc_hd__nand3_1 _09585_ (.A(net181),
    .B(_02501_),
    .C(_02502_),
    .Y(_02504_));
 sky130_fd_sc_hd__nand3_2 _09586_ (.A(_06736_),
    .B(_02503_),
    .C(_02504_),
    .Y(_02505_));
 sky130_fd_sc_hd__a21o_1 _09587_ (.A1(_02503_),
    .A2(_02504_),
    .B1(_06736_),
    .X(_02506_));
 sky130_fd_sc_hd__nand3_2 _09588_ (.A(_02500_),
    .B(_02505_),
    .C(_02506_),
    .Y(_02507_));
 sky130_fd_sc_hd__a21o_1 _09589_ (.A1(_02505_),
    .A2(_02506_),
    .B1(_02500_),
    .X(_02508_));
 sky130_fd_sc_hd__o22a_1 _09590_ (.A1(net100),
    .A2(net83),
    .B1(net79),
    .B2(net42),
    .X(_02509_));
 sky130_fd_sc_hd__xnor2_1 _09591_ (.A(net116),
    .B(_02509_),
    .Y(_02510_));
 sky130_fd_sc_hd__inv_2 _09592_ (.A(_02510_),
    .Y(_02511_));
 sky130_fd_sc_hd__o22a_1 _09593_ (.A1(net103),
    .A2(net23),
    .B1(net70),
    .B2(net25),
    .X(_02512_));
 sky130_fd_sc_hd__xnor2_2 _09594_ (.A(net86),
    .B(_02512_),
    .Y(_02513_));
 sky130_fd_sc_hd__o22a_1 _09595_ (.A1(net40),
    .A2(net75),
    .B1(net72),
    .B2(net56),
    .X(_02514_));
 sky130_fd_sc_hd__xnor2_2 _09596_ (.A(net108),
    .B(_02514_),
    .Y(_02515_));
 sky130_fd_sc_hd__nand2_1 _09597_ (.A(_02513_),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__xnor2_2 _09598_ (.A(_02513_),
    .B(_02515_),
    .Y(_02517_));
 sky130_fd_sc_hd__xnor2_1 _09599_ (.A(_02510_),
    .B(_02517_),
    .Y(_02518_));
 sky130_fd_sc_hd__nand3_2 _09600_ (.A(_02507_),
    .B(_02508_),
    .C(_02518_),
    .Y(_02519_));
 sky130_fd_sc_hd__a21o_1 _09601_ (.A1(_02507_),
    .A2(_02508_),
    .B1(_02518_),
    .X(_02520_));
 sky130_fd_sc_hd__nand3_1 _09602_ (.A(_02498_),
    .B(_02519_),
    .C(_02520_),
    .Y(_02521_));
 sky130_fd_sc_hd__a21o_1 _09603_ (.A1(_02519_),
    .A2(_02520_),
    .B1(_02498_),
    .X(_02522_));
 sky130_fd_sc_hd__nand2_1 _09604_ (.A(net153),
    .B(net63),
    .Y(_02523_));
 sky130_fd_sc_hd__o21a_1 _09605_ (.A1(_02291_),
    .A2(_02296_),
    .B1(_02295_),
    .X(_02524_));
 sky130_fd_sc_hd__a22o_1 _09606_ (.A1(net148),
    .A2(net9),
    .B1(net4),
    .B2(net150),
    .X(_02525_));
 sky130_fd_sc_hd__xnor2_1 _09607_ (.A(net60),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__and2b_1 _09608_ (.A_N(_02524_),
    .B(_02526_),
    .X(_02527_));
 sky130_fd_sc_hd__xnor2_1 _09609_ (.A(_02524_),
    .B(_02526_),
    .Y(_02528_));
 sky130_fd_sc_hd__xnor2_1 _09610_ (.A(_02523_),
    .B(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__and3_1 _09611_ (.A(_02521_),
    .B(_02522_),
    .C(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__a21oi_1 _09612_ (.A1(_02521_),
    .A2(_02522_),
    .B1(_02529_),
    .Y(_02531_));
 sky130_fd_sc_hd__nor3_1 _09613_ (.A(_02487_),
    .B(_02530_),
    .C(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__o21a_1 _09614_ (.A1(_02530_),
    .A2(_02531_),
    .B1(_02487_),
    .X(_02533_));
 sky130_fd_sc_hd__nor2_1 _09615_ (.A(_02532_),
    .B(_02533_),
    .Y(_02534_));
 sky130_fd_sc_hd__o21ai_2 _09616_ (.A1(_02251_),
    .A2(_02257_),
    .B1(_02256_),
    .Y(_02535_));
 sky130_fd_sc_hd__inv_2 _09617_ (.A(_02535_),
    .Y(_02536_));
 sky130_fd_sc_hd__o22a_1 _09618_ (.A1(net85),
    .A2(net21),
    .B1(net19),
    .B2(_00442_),
    .X(_02537_));
 sky130_fd_sc_hd__xnor2_2 _09619_ (.A(net97),
    .B(_02537_),
    .Y(_02538_));
 sky130_fd_sc_hd__o22a_1 _09620_ (.A1(net39),
    .A2(net120),
    .B1(_00391_),
    .B2(net37),
    .X(_02539_));
 sky130_fd_sc_hd__xnor2_1 _09621_ (.A(net99),
    .B(_02539_),
    .Y(_02540_));
 sky130_fd_sc_hd__o22a_1 _09622_ (.A1(net28),
    .A2(net76),
    .B1(net74),
    .B2(net26),
    .X(_02541_));
 sky130_fd_sc_hd__xnor2_1 _09623_ (.A(net88),
    .B(_02541_),
    .Y(_02542_));
 sky130_fd_sc_hd__and2_1 _09624_ (.A(_02540_),
    .B(_02542_),
    .X(_02543_));
 sky130_fd_sc_hd__or2_1 _09625_ (.A(_02540_),
    .B(_02542_),
    .X(_02544_));
 sky130_fd_sc_hd__nand2b_1 _09626_ (.A_N(_02543_),
    .B(_02544_),
    .Y(_02545_));
 sky130_fd_sc_hd__xnor2_2 _09627_ (.A(_02538_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__a21o_1 _09628_ (.A1(_02301_),
    .A2(_02306_),
    .B1(_02305_),
    .X(_02547_));
 sky130_fd_sc_hd__nand2_1 _09629_ (.A(_02546_),
    .B(_02547_),
    .Y(_02548_));
 sky130_fd_sc_hd__xnor2_1 _09630_ (.A(_02546_),
    .B(_02547_),
    .Y(_02549_));
 sky130_fd_sc_hd__xnor2_1 _09631_ (.A(_02535_),
    .B(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__and2_1 _09632_ (.A(_02534_),
    .B(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__nor2_1 _09633_ (.A(_02534_),
    .B(_02550_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_2 _09634_ (.A(_02551_),
    .B(_02552_),
    .Y(_02553_));
 sky130_fd_sc_hd__xor2_4 _09635_ (.A(_02481_),
    .B(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__a21o_1 _09636_ (.A1(_02262_),
    .A2(_02329_),
    .B1(_02327_),
    .X(_02555_));
 sky130_fd_sc_hd__o21bai_2 _09637_ (.A1(_02258_),
    .A2(_02259_),
    .B1_N(_02261_),
    .Y(_02556_));
 sky130_fd_sc_hd__o21a_1 _09638_ (.A1(_02269_),
    .A2(_02309_),
    .B1(_02308_),
    .X(_02557_));
 sky130_fd_sc_hd__o21ba_1 _09639_ (.A1(_02312_),
    .A2(_02325_),
    .B1_N(_02324_),
    .X(_02558_));
 sky130_fd_sc_hd__nor2_1 _09640_ (.A(_02557_),
    .B(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__xor2_2 _09641_ (.A(_02557_),
    .B(_02558_),
    .X(_02560_));
 sky130_fd_sc_hd__xnor2_2 _09642_ (.A(_02556_),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__a21oi_4 _09643_ (.A1(_02332_),
    .A2(_02336_),
    .B1(_02335_),
    .Y(_02562_));
 sky130_fd_sc_hd__xnor2_2 _09644_ (.A(_02561_),
    .B(_02562_),
    .Y(_02563_));
 sky130_fd_sc_hd__nand2b_1 _09645_ (.A_N(_02563_),
    .B(_02555_),
    .Y(_02564_));
 sky130_fd_sc_hd__xnor2_2 _09646_ (.A(_02555_),
    .B(_02563_),
    .Y(_02565_));
 sky130_fd_sc_hd__and2_1 _09647_ (.A(_02554_),
    .B(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__xor2_4 _09648_ (.A(_02554_),
    .B(_02565_),
    .X(_02567_));
 sky130_fd_sc_hd__xnor2_4 _09649_ (.A(_02465_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__xnor2_4 _09650_ (.A(_02464_),
    .B(_02568_),
    .Y(_02569_));
 sky130_fd_sc_hd__a2111o_1 _09651_ (.A1(_01027_),
    .A2(_01920_),
    .B1(_02233_),
    .C1(_02236_),
    .D1(_02346_),
    .X(_02570_));
 sky130_fd_sc_hd__o2bb2a_1 _09652_ (.A1_N(_02129_),
    .A2_N(_02231_),
    .B1(_02246_),
    .B2(_02344_),
    .X(_02571_));
 sky130_fd_sc_hd__o32a_1 _09653_ (.A1(_02233_),
    .A2(_02235_),
    .A3(_02346_),
    .B1(_02571_),
    .B2(_02345_),
    .X(_02572_));
 sky130_fd_sc_hd__nand2_1 _09654_ (.A(_02570_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__xor2_2 _09655_ (.A(_02569_),
    .B(_02573_),
    .X(_02574_));
 sky130_fd_sc_hd__or3_1 _09656_ (.A(net135),
    .B(_02463_),
    .C(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__o21ai_1 _09657_ (.A1(net135),
    .A2(_02463_),
    .B1(_02574_),
    .Y(_02576_));
 sky130_fd_sc_hd__and3_1 _09658_ (.A(_02348_),
    .B(_02575_),
    .C(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__or2_1 _09659_ (.A(_06637_),
    .B(net197),
    .X(_02578_));
 sky130_fd_sc_hd__xnor2_1 _09660_ (.A(_01875_),
    .B(_02578_),
    .Y(_02579_));
 sky130_fd_sc_hd__o21ai_1 _09661_ (.A1(_06637_),
    .A2(net135),
    .B1(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__o311a_1 _09662_ (.A1(_06637_),
    .A2(net134),
    .A3(_02579_),
    .B1(_02580_),
    .C1(net233),
    .X(_02581_));
 sky130_fd_sc_hd__mux2_1 _09663_ (.A0(_02356_),
    .A1(_02361_),
    .S(net206),
    .X(_02582_));
 sky130_fd_sc_hd__mux2_1 _09664_ (.A0(_02360_),
    .A1(_02367_),
    .S(net206),
    .X(_02583_));
 sky130_fd_sc_hd__mux2_1 _09665_ (.A0(_02582_),
    .A1(_02583_),
    .S(_06569_),
    .X(_02584_));
 sky130_fd_sc_hd__mux2_1 _09666_ (.A0(_02363_),
    .A1(_02383_),
    .S(net206),
    .X(_02585_));
 sky130_fd_sc_hd__mux2_1 _09667_ (.A0(_02364_),
    .A1(_02366_),
    .S(net208),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _09668_ (.A0(_02585_),
    .A1(_02586_),
    .S(net213),
    .X(_02587_));
 sky130_fd_sc_hd__mux2_1 _09669_ (.A0(_02584_),
    .A1(_02587_),
    .S(net215),
    .X(_02588_));
 sky130_fd_sc_hd__mux2_1 _09670_ (.A0(_02372_),
    .A1(_02398_),
    .S(net206),
    .X(_02589_));
 sky130_fd_sc_hd__mux2_1 _09671_ (.A0(_02373_),
    .A1(_02375_),
    .S(net209),
    .X(_02590_));
 sky130_fd_sc_hd__mux2_1 _09672_ (.A0(_02589_),
    .A1(_02590_),
    .S(net213),
    .X(_02591_));
 sky130_fd_sc_hd__mux2_1 _09673_ (.A0(_02376_),
    .A1(_02379_),
    .S(net208),
    .X(_02592_));
 sky130_fd_sc_hd__mux2_1 _09674_ (.A0(_02380_),
    .A1(_02382_),
    .S(net208),
    .X(_02593_));
 sky130_fd_sc_hd__mux2_1 _09675_ (.A0(_02592_),
    .A1(_02593_),
    .S(net213),
    .X(_02594_));
 sky130_fd_sc_hd__mux2_1 _09676_ (.A0(_02591_),
    .A1(_02594_),
    .S(net217),
    .X(_02595_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(_02588_),
    .A1(_02595_),
    .S(net218),
    .X(_02596_));
 sky130_fd_sc_hd__mux2_1 _09678_ (.A0(_02387_),
    .A1(_02413_),
    .S(net206),
    .X(_02597_));
 sky130_fd_sc_hd__mux2_1 _09679_ (.A0(_02388_),
    .A1(_02390_),
    .S(net210),
    .X(_02598_));
 sky130_fd_sc_hd__mux2_1 _09680_ (.A0(_02597_),
    .A1(_02598_),
    .S(net213),
    .X(_02599_));
 sky130_fd_sc_hd__mux2_1 _09681_ (.A0(_02391_),
    .A1(_02394_),
    .S(net210),
    .X(_02600_));
 sky130_fd_sc_hd__mux2_1 _09682_ (.A0(_02395_),
    .A1(_02397_),
    .S(net210),
    .X(_02601_));
 sky130_fd_sc_hd__mux2_1 _09683_ (.A0(_02600_),
    .A1(_02601_),
    .S(net213),
    .X(_02602_));
 sky130_fd_sc_hd__mux2_1 _09684_ (.A0(_02599_),
    .A1(_02602_),
    .S(net217),
    .X(_02603_));
 sky130_fd_sc_hd__mux2_1 _09685_ (.A0(_02403_),
    .A1(_02405_),
    .S(net211),
    .X(_02604_));
 sky130_fd_sc_hd__mux2_1 _09686_ (.A0(_02450_),
    .A1(_02604_),
    .S(net214),
    .X(_02605_));
 sky130_fd_sc_hd__mux2_1 _09687_ (.A0(_02406_),
    .A1(_02409_),
    .S(net210),
    .X(_02606_));
 sky130_fd_sc_hd__mux2_1 _09688_ (.A0(_02410_),
    .A1(_02412_),
    .S(net210),
    .X(_02607_));
 sky130_fd_sc_hd__mux2_1 _09689_ (.A0(_02606_),
    .A1(_02607_),
    .S(net213),
    .X(_02608_));
 sky130_fd_sc_hd__mux2_1 _09690_ (.A0(_02605_),
    .A1(_02608_),
    .S(net217),
    .X(_02609_));
 sky130_fd_sc_hd__mux2_1 _09691_ (.A0(_02603_),
    .A1(_02609_),
    .S(net219),
    .X(_02610_));
 sky130_fd_sc_hd__mux2_2 _09692_ (.A0(_02596_),
    .A1(_02610_),
    .S(net221),
    .X(_02611_));
 sky130_fd_sc_hd__nand2_1 _09693_ (.A(net289),
    .B(curr_PC[1]),
    .Y(_02612_));
 sky130_fd_sc_hd__or2_1 _09694_ (.A(net289),
    .B(curr_PC[1]),
    .X(_02613_));
 sky130_fd_sc_hd__nand2_1 _09695_ (.A(_02612_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__xnor2_1 _09696_ (.A(_02420_),
    .B(_02614_),
    .Y(_02615_));
 sky130_fd_sc_hd__nand2_1 _09697_ (.A(net244),
    .B(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__o211a_1 _09698_ (.A1(net244),
    .A2(_02611_),
    .B1(_02616_),
    .C1(net205),
    .X(_02617_));
 sky130_fd_sc_hd__a21oi_1 _09699_ (.A1(\div_res[0] ),
    .A2(net140),
    .B1(\div_res[1] ),
    .Y(_02618_));
 sky130_fd_sc_hd__a31o_1 _09700_ (.A1(\div_res[1] ),
    .A2(\div_res[0] ),
    .A3(net140),
    .B1(net190),
    .X(_02619_));
 sky130_fd_sc_hd__nand2_1 _09701_ (.A(_06574_),
    .B(_06578_),
    .Y(_02620_));
 sky130_fd_sc_hd__a22oi_1 _09702_ (.A1(net283),
    .A2(net206),
    .B1(_06579_),
    .B2(_02620_),
    .Y(_02621_));
 sky130_fd_sc_hd__and4_1 _09703_ (.A(net283),
    .B(net206),
    .C(_06579_),
    .D(_02620_),
    .X(_02622_));
 sky130_fd_sc_hd__o21a_1 _09704_ (.A1(_06571_),
    .A2(_02429_),
    .B1(_02440_),
    .X(_02623_));
 sky130_fd_sc_hd__and2_1 _09705_ (.A(divi1_sign),
    .B(net296),
    .X(_02624_));
 sky130_fd_sc_hd__a21oi_4 _09706_ (.A1(\div_shifter[32] ),
    .A2(net230),
    .B1(\div_shifter[33] ),
    .Y(_02625_));
 sky130_fd_sc_hd__a31o_1 _09707_ (.A1(\div_shifter[33] ),
    .A2(\div_shifter[32] ),
    .A3(net230),
    .B1(net192),
    .X(_02626_));
 sky130_fd_sc_hd__o2bb2a_1 _09708_ (.A1_N(_06734_),
    .A2_N(net256),
    .B1(net231),
    .B2(reg1_val[1]),
    .X(_02627_));
 sky130_fd_sc_hd__o221a_1 _09709_ (.A1(net214),
    .A2(net203),
    .B1(_02625_),
    .B2(_02626_),
    .C1(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__o221a_1 _09710_ (.A1(_06572_),
    .A2(net194),
    .B1(_02623_),
    .B2(_06573_),
    .C1(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__o31a_1 _09711_ (.A1(_02427_),
    .A2(_02621_),
    .A3(_02622_),
    .B1(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _09712_ (.A0(_02404_),
    .A1(_02449_),
    .S(_06569_),
    .X(_02631_));
 sky130_fd_sc_hd__o21a_1 _09713_ (.A1(net215),
    .A2(_02631_),
    .B1(_02452_),
    .X(_02632_));
 sky130_fd_sc_hd__o21a_1 _09714_ (.A1(net219),
    .A2(_02632_),
    .B1(_02453_),
    .X(_02633_));
 sky130_fd_sc_hd__o21ai_2 _09715_ (.A1(net221),
    .A2(_02633_),
    .B1(_02456_),
    .Y(_02634_));
 sky130_fd_sc_hd__inv_2 _09716_ (.A(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__o221ai_1 _09717_ (.A1(_02618_),
    .A2(_02619_),
    .B1(_02634_),
    .B2(net169),
    .C1(_02630_),
    .Y(_02636_));
 sky130_fd_sc_hd__a211o_1 _09718_ (.A1(net167),
    .A2(_02611_),
    .B1(_02617_),
    .C1(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__o31a_1 _09719_ (.A1(_02577_),
    .A2(_02581_),
    .A3(_02637_),
    .B1(net241),
    .X(_02638_));
 sky130_fd_sc_hd__or2_1 _09720_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .X(_02639_));
 sky130_fd_sc_hd__nand2_1 _09721_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .Y(_02640_));
 sky130_fd_sc_hd__a31o_4 _09722_ (.A1(net242),
    .A2(_02639_),
    .A3(_02640_),
    .B1(_02638_),
    .X(dest_val[1]));
 sky130_fd_sc_hd__a21oi_1 _09723_ (.A1(_02463_),
    .A2(_02574_),
    .B1(net135),
    .Y(_02641_));
 sky130_fd_sc_hd__a21oi_4 _09724_ (.A1(_02465_),
    .A2(_02567_),
    .B1(_02566_),
    .Y(_02642_));
 sky130_fd_sc_hd__o21ai_4 _09725_ (.A1(_02561_),
    .A2(_02562_),
    .B1(_02564_),
    .Y(_02643_));
 sky130_fd_sc_hd__nand2_2 _09726_ (.A(_02519_),
    .B(_02521_),
    .Y(_02644_));
 sky130_fd_sc_hd__o22a_2 _09727_ (.A1(net35),
    .A2(net113),
    .B1(net110),
    .B2(net33),
    .X(_02645_));
 sky130_fd_sc_hd__xnor2_4 _09728_ (.A(net95),
    .B(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__a22o_2 _09729_ (.A1(net107),
    .A2(net17),
    .B1(net13),
    .B2(_00287_),
    .X(_02647_));
 sky130_fd_sc_hd__xnor2_4 _09730_ (.A(net65),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__a22o_1 _09731_ (.A1(net14),
    .A2(net122),
    .B1(_00375_),
    .B2(net30),
    .X(_02649_));
 sky130_fd_sc_hd__xnor2_4 _09732_ (.A(net91),
    .B(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__nand2_1 _09733_ (.A(_02648_),
    .B(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__xnor2_4 _09734_ (.A(_02648_),
    .B(_02650_),
    .Y(_02652_));
 sky130_fd_sc_hd__inv_2 _09735_ (.A(_02652_),
    .Y(_02653_));
 sky130_fd_sc_hd__xor2_4 _09736_ (.A(_02646_),
    .B(_02652_),
    .X(_02654_));
 sky130_fd_sc_hd__a21oi_4 _09737_ (.A1(_02482_),
    .A2(_02486_),
    .B1(_02485_),
    .Y(_02655_));
 sky130_fd_sc_hd__xnor2_4 _09738_ (.A(_02654_),
    .B(_02655_),
    .Y(_02656_));
 sky130_fd_sc_hd__nand2b_1 _09739_ (.A_N(_02656_),
    .B(_02644_),
    .Y(_02657_));
 sky130_fd_sc_hd__xnor2_4 _09740_ (.A(_02644_),
    .B(_02656_),
    .Y(_02658_));
 sky130_fd_sc_hd__o21ai_2 _09741_ (.A1(_02511_),
    .A2(_02517_),
    .B1(_02516_),
    .Y(_02659_));
 sky130_fd_sc_hd__a21oi_2 _09742_ (.A1(_02538_),
    .A2(_02544_),
    .B1(_02543_),
    .Y(_02660_));
 sky130_fd_sc_hd__o21a_1 _09743_ (.A1(_02490_),
    .A2(_02497_),
    .B1(_02495_),
    .X(_02661_));
 sky130_fd_sc_hd__or2_1 _09744_ (.A(_02660_),
    .B(_02661_),
    .X(_02662_));
 sky130_fd_sc_hd__xor2_1 _09745_ (.A(_02660_),
    .B(_02661_),
    .X(_02663_));
 sky130_fd_sc_hd__nand2_1 _09746_ (.A(_02659_),
    .B(_02663_),
    .Y(_02664_));
 sky130_fd_sc_hd__xnor2_1 _09747_ (.A(_02659_),
    .B(_02663_),
    .Y(_02665_));
 sky130_fd_sc_hd__nand2_1 _09748_ (.A(_00327_),
    .B(net63),
    .Y(_02666_));
 sky130_fd_sc_hd__a22o_1 _09749_ (.A1(_00266_),
    .A2(net9),
    .B1(net4),
    .B2(net148),
    .X(_02667_));
 sky130_fd_sc_hd__xnor2_1 _09750_ (.A(net60),
    .B(_02667_),
    .Y(_02668_));
 sky130_fd_sc_hd__inv_2 _09751_ (.A(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__a21oi_1 _09752_ (.A1(_02505_),
    .A2(_02507_),
    .B1(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__nand3_1 _09753_ (.A(_02505_),
    .B(_02507_),
    .C(_02669_),
    .Y(_02671_));
 sky130_fd_sc_hd__and2b_1 _09754_ (.A_N(_02670_),
    .B(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__xnor2_1 _09755_ (.A(_02666_),
    .B(_02672_),
    .Y(_02673_));
 sky130_fd_sc_hd__a22o_1 _09756_ (.A1(_00144_),
    .A2(net129),
    .B1(net127),
    .B2(_00136_),
    .X(_02674_));
 sky130_fd_sc_hd__xnor2_1 _09757_ (.A(net155),
    .B(_02674_),
    .Y(_02675_));
 sky130_fd_sc_hd__o22a_1 _09758_ (.A1(net47),
    .A2(net68),
    .B1(net66),
    .B2(net45),
    .X(_02676_));
 sky130_fd_sc_hd__xnor2_1 _09759_ (.A(net145),
    .B(_02676_),
    .Y(_02677_));
 sky130_fd_sc_hd__o32a_1 _09760_ (.A1(net131),
    .A2(_00513_),
    .A3(_00515_),
    .B1(net105),
    .B2(net44),
    .X(_02678_));
 sky130_fd_sc_hd__xnor2_1 _09761_ (.A(net174),
    .B(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__nand2_1 _09762_ (.A(_02677_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__xnor2_1 _09763_ (.A(_02677_),
    .B(_02679_),
    .Y(_02681_));
 sky130_fd_sc_hd__or2_1 _09764_ (.A(_02675_),
    .B(_02681_),
    .X(_02682_));
 sky130_fd_sc_hd__nand2_1 _09765_ (.A(_02675_),
    .B(_02681_),
    .Y(_02683_));
 sky130_fd_sc_hd__nand2_1 _09766_ (.A(_02682_),
    .B(_02683_),
    .Y(_02684_));
 sky130_fd_sc_hd__o22a_2 _09767_ (.A1(net42),
    .A2(net83),
    .B1(net79),
    .B2(net40),
    .X(_02685_));
 sky130_fd_sc_hd__xnor2_4 _09768_ (.A(net118),
    .B(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__o22a_1 _09769_ (.A1(net103),
    .A2(net24),
    .B1(net22),
    .B2(net100),
    .X(_02687_));
 sky130_fd_sc_hd__xnor2_1 _09770_ (.A(net86),
    .B(_02687_),
    .Y(_02688_));
 sky130_fd_sc_hd__o22a_1 _09771_ (.A1(net56),
    .A2(net75),
    .B1(net72),
    .B2(net53),
    .X(_02689_));
 sky130_fd_sc_hd__xnor2_1 _09772_ (.A(net108),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__and2_1 _09773_ (.A(_02688_),
    .B(_02690_),
    .X(_02691_));
 sky130_fd_sc_hd__or2_1 _09774_ (.A(_02688_),
    .B(_02690_),
    .X(_02692_));
 sky130_fd_sc_hd__nand2b_2 _09775_ (.A_N(_02691_),
    .B(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__xor2_4 _09776_ (.A(_02686_),
    .B(_02693_),
    .X(_02694_));
 sky130_fd_sc_hd__a22o_1 _09777_ (.A1(_06702_),
    .A2(_00812_),
    .B1(net11),
    .B2(_06726_),
    .X(_02695_));
 sky130_fd_sc_hd__xnor2_2 _09778_ (.A(net181),
    .B(_02695_),
    .Y(_02696_));
 sky130_fd_sc_hd__and2_1 _09779_ (.A(_06736_),
    .B(_02696_),
    .X(_02697_));
 sky130_fd_sc_hd__xnor2_4 _09780_ (.A(net198),
    .B(_02696_),
    .Y(_02698_));
 sky130_fd_sc_hd__a21oi_1 _09781_ (.A1(_00154_),
    .A2(net6),
    .B1(net202),
    .Y(_02699_));
 sky130_fd_sc_hd__a31o_2 _09782_ (.A1(net202),
    .A2(_00155_),
    .A3(net6),
    .B1(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__xnor2_4 _09783_ (.A(_02698_),
    .B(_02700_),
    .Y(_02701_));
 sky130_fd_sc_hd__nor2_1 _09784_ (.A(_02694_),
    .B(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__xor2_4 _09785_ (.A(_02694_),
    .B(_02701_),
    .X(_02703_));
 sky130_fd_sc_hd__xnor2_2 _09786_ (.A(_02684_),
    .B(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__nand2_1 _09787_ (.A(_02673_),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__xnor2_1 _09788_ (.A(_02673_),
    .B(_02704_),
    .Y(_02706_));
 sky130_fd_sc_hd__xor2_1 _09789_ (.A(_02665_),
    .B(_02706_),
    .X(_02707_));
 sky130_fd_sc_hd__a21bo_1 _09790_ (.A1(_02468_),
    .A2(_02475_),
    .B1_N(_02473_),
    .X(_02708_));
 sky130_fd_sc_hd__o22a_1 _09791_ (.A1(net21),
    .A2(_00442_),
    .B1(net77),
    .B2(net19),
    .X(_02709_));
 sky130_fd_sc_hd__xnor2_1 _09792_ (.A(net97),
    .B(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__o22a_1 _09793_ (.A1(net28),
    .A2(net74),
    .B1(net70),
    .B2(net26),
    .X(_02711_));
 sky130_fd_sc_hd__xnor2_1 _09794_ (.A(net88),
    .B(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__o22a_1 _09795_ (.A1(net39),
    .A2(_00391_),
    .B1(_00398_),
    .B2(net37),
    .X(_02713_));
 sky130_fd_sc_hd__xnor2_1 _09796_ (.A(net99),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__and2_1 _09797_ (.A(_02712_),
    .B(_02714_),
    .X(_02715_));
 sky130_fd_sc_hd__or2_1 _09798_ (.A(_02712_),
    .B(_02714_),
    .X(_02716_));
 sky130_fd_sc_hd__nand2b_1 _09799_ (.A_N(_02715_),
    .B(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__xnor2_1 _09800_ (.A(_02710_),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__a31o_1 _09801_ (.A1(net153),
    .A2(net63),
    .A3(_02528_),
    .B1(_02527_),
    .X(_02719_));
 sky130_fd_sc_hd__xnor2_1 _09802_ (.A(_02718_),
    .B(_02719_),
    .Y(_02720_));
 sky130_fd_sc_hd__and2b_1 _09803_ (.A_N(_02720_),
    .B(_02708_),
    .X(_02721_));
 sky130_fd_sc_hd__xnor2_1 _09804_ (.A(_02708_),
    .B(_02720_),
    .Y(_02722_));
 sky130_fd_sc_hd__and2_1 _09805_ (.A(_02707_),
    .B(_02722_),
    .X(_02723_));
 sky130_fd_sc_hd__nor2_1 _09806_ (.A(_02707_),
    .B(_02722_),
    .Y(_02724_));
 sky130_fd_sc_hd__nor2_2 _09807_ (.A(_02723_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__xor2_4 _09808_ (.A(_02658_),
    .B(_02725_),
    .X(_02726_));
 sky130_fd_sc_hd__a21o_2 _09809_ (.A1(_02481_),
    .A2(_02553_),
    .B1(_02551_),
    .X(_02727_));
 sky130_fd_sc_hd__a21o_1 _09810_ (.A1(_02556_),
    .A2(_02560_),
    .B1(_02559_),
    .X(_02728_));
 sky130_fd_sc_hd__or2_2 _09811_ (.A(_02477_),
    .B(_02480_),
    .X(_02729_));
 sky130_fd_sc_hd__or2_1 _09812_ (.A(_02530_),
    .B(_02532_),
    .X(_02730_));
 sky130_fd_sc_hd__o21a_1 _09813_ (.A1(_02536_),
    .A2(_02549_),
    .B1(_02548_),
    .X(_02731_));
 sky130_fd_sc_hd__o21ba_1 _09814_ (.A1(_02530_),
    .A2(_02532_),
    .B1_N(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__xnor2_2 _09815_ (.A(_02730_),
    .B(_02731_),
    .Y(_02733_));
 sky130_fd_sc_hd__xor2_2 _09816_ (.A(_02729_),
    .B(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__xnor2_2 _09817_ (.A(_02728_),
    .B(_02734_),
    .Y(_02735_));
 sky130_fd_sc_hd__nand2b_1 _09818_ (.A_N(_02735_),
    .B(_02727_),
    .Y(_02736_));
 sky130_fd_sc_hd__xnor2_4 _09819_ (.A(_02727_),
    .B(_02735_),
    .Y(_02737_));
 sky130_fd_sc_hd__and2_1 _09820_ (.A(_02726_),
    .B(_02737_),
    .X(_02738_));
 sky130_fd_sc_hd__xor2_4 _09821_ (.A(_02726_),
    .B(_02737_),
    .X(_02739_));
 sky130_fd_sc_hd__xnor2_4 _09822_ (.A(_02643_),
    .B(_02739_),
    .Y(_02740_));
 sky130_fd_sc_hd__or2_1 _09823_ (.A(_02642_),
    .B(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__xnor2_4 _09824_ (.A(_02642_),
    .B(_02740_),
    .Y(_02742_));
 sky130_fd_sc_hd__or4_1 _09825_ (.A(_02123_),
    .B(_02233_),
    .C(_02346_),
    .D(_02569_),
    .X(_02743_));
 sky130_fd_sc_hd__o22a_1 _09826_ (.A1(_02246_),
    .A2(_02344_),
    .B1(_02464_),
    .B2(_02568_),
    .X(_02744_));
 sky130_fd_sc_hd__a21o_1 _09827_ (.A1(_02464_),
    .A2(_02568_),
    .B1(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__or4_1 _09828_ (.A(_02232_),
    .B(_02243_),
    .C(_02346_),
    .D(_02569_),
    .X(_02746_));
 sky130_fd_sc_hd__o211a_2 _09829_ (.A1(_02127_),
    .A2(_02743_),
    .B1(_02745_),
    .C1(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__xor2_2 _09830_ (.A(_02742_),
    .B(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__a21o_1 _09831_ (.A1(_02641_),
    .A2(_02748_),
    .B1(net235),
    .X(_02749_));
 sky130_fd_sc_hd__o21ba_1 _09832_ (.A1(_02641_),
    .A2(_02748_),
    .B1_N(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__o21bai_1 _09833_ (.A1(net135),
    .A2(_01876_),
    .B1_N(_01925_),
    .Y(_02751_));
 sky130_fd_sc_hd__o311a_1 _09834_ (.A1(net135),
    .A2(_01874_),
    .A3(_01876_),
    .B1(net233),
    .C1(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__o21a_1 _09835_ (.A1(net215),
    .A2(_02605_),
    .B1(_02452_),
    .X(_02753_));
 sky130_fd_sc_hd__o21a_1 _09836_ (.A1(net218),
    .A2(_02753_),
    .B1(_02453_),
    .X(_02754_));
 sky130_fd_sc_hd__o21ai_2 _09837_ (.A1(net221),
    .A2(_02754_),
    .B1(_02456_),
    .Y(_02755_));
 sky130_fd_sc_hd__inv_2 _09838_ (.A(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__nor2_1 _09839_ (.A(net169),
    .B(_02755_),
    .Y(_02757_));
 sky130_fd_sc_hd__mux2_1 _09840_ (.A0(_02362_),
    .A1(_02368_),
    .S(_06569_),
    .X(_02758_));
 sky130_fd_sc_hd__mux2_1 _09841_ (.A0(_02365_),
    .A1(_02384_),
    .S(_06569_),
    .X(_02759_));
 sky130_fd_sc_hd__mux2_1 _09842_ (.A0(_02758_),
    .A1(_02759_),
    .S(net215),
    .X(_02760_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(_02374_),
    .A1(_02399_),
    .S(_06569_),
    .X(_02761_));
 sky130_fd_sc_hd__mux2_1 _09844_ (.A0(_02377_),
    .A1(_02381_),
    .S(net213),
    .X(_02762_));
 sky130_fd_sc_hd__mux2_1 _09845_ (.A0(_02761_),
    .A1(_02762_),
    .S(net217),
    .X(_02763_));
 sky130_fd_sc_hd__mux2_1 _09846_ (.A0(_02760_),
    .A1(_02763_),
    .S(net218),
    .X(_02764_));
 sky130_fd_sc_hd__mux2_1 _09847_ (.A0(_02389_),
    .A1(_02414_),
    .S(_06569_),
    .X(_02765_));
 sky130_fd_sc_hd__mux2_1 _09848_ (.A0(_02392_),
    .A1(_02396_),
    .S(net213),
    .X(_02766_));
 sky130_fd_sc_hd__mux2_1 _09849_ (.A0(_02765_),
    .A1(_02766_),
    .S(net217),
    .X(_02767_));
 sky130_fd_sc_hd__mux2_1 _09850_ (.A0(_02407_),
    .A1(_02411_),
    .S(net214),
    .X(_02768_));
 sky130_fd_sc_hd__mux2_1 _09851_ (.A0(_02631_),
    .A1(_02768_),
    .S(net217),
    .X(_02769_));
 sky130_fd_sc_hd__mux2_1 _09852_ (.A0(_02767_),
    .A1(_02769_),
    .S(net218),
    .X(_02770_));
 sky130_fd_sc_hd__mux2_1 _09853_ (.A0(_02764_),
    .A1(_02770_),
    .S(net221),
    .X(_02771_));
 sky130_fd_sc_hd__o21a_1 _09854_ (.A1(_02420_),
    .A2(_02614_),
    .B1(_02612_),
    .X(_02772_));
 sky130_fd_sc_hd__nor2_1 _09855_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02773_));
 sky130_fd_sc_hd__nand2_1 _09856_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02774_));
 sky130_fd_sc_hd__nand2b_1 _09857_ (.A_N(_02773_),
    .B(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__xnor2_2 _09858_ (.A(_02772_),
    .B(_02775_),
    .Y(_02776_));
 sky130_fd_sc_hd__a21o_1 _09859_ (.A1(net244),
    .A2(_02776_),
    .B1(_06667_),
    .X(_02777_));
 sky130_fd_sc_hd__nand2_1 _09860_ (.A(_02425_),
    .B(_02777_),
    .Y(_02778_));
 sky130_fd_sc_hd__o21ai_1 _09861_ (.A1(\div_res[1] ),
    .A2(\div_res[0] ),
    .B1(net140),
    .Y(_02779_));
 sky130_fd_sc_hd__xnor2_1 _09862_ (.A(\div_res[2] ),
    .B(_02779_),
    .Y(_02780_));
 sky130_fd_sc_hd__a21o_1 _09863_ (.A1(_06572_),
    .A2(_06637_),
    .B1(_06573_),
    .X(_02781_));
 sky130_fd_sc_hd__a21o_1 _09864_ (.A1(_06570_),
    .A2(_06579_),
    .B1(net283),
    .X(_02782_));
 sky130_fd_sc_hd__nand2_1 _09865_ (.A(net283),
    .B(_02781_),
    .Y(_02783_));
 sky130_fd_sc_hd__a21oi_1 _09866_ (.A1(_02782_),
    .A2(_02783_),
    .B1(_06565_),
    .Y(_02784_));
 sky130_fd_sc_hd__a31o_1 _09867_ (.A1(_06565_),
    .A2(_02782_),
    .A3(_02783_),
    .B1(_02427_),
    .X(_02785_));
 sky130_fd_sc_hd__a21oi_1 _09868_ (.A1(_06563_),
    .A2(net195),
    .B1(net193),
    .Y(_02786_));
 sky130_fd_sc_hd__o21a_1 _09869_ (.A1(\div_shifter[33] ),
    .A2(\div_shifter[32] ),
    .B1(net230),
    .X(_02787_));
 sky130_fd_sc_hd__xnor2_2 _09870_ (.A(\div_shifter[34] ),
    .B(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand3_2 _09871_ (.A(_06684_),
    .B(_00151_),
    .C(net256),
    .Y(_02789_));
 sky130_fd_sc_hd__o221a_1 _09872_ (.A1(reg1_val[2]),
    .A2(net232),
    .B1(_02788_),
    .B2(net192),
    .C1(_02789_),
    .X(_02790_));
 sky130_fd_sc_hd__o221a_1 _09873_ (.A1(_06560_),
    .A2(net203),
    .B1(net194),
    .B2(_06563_),
    .C1(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__o221a_1 _09874_ (.A1(net223),
    .A2(_02777_),
    .B1(_02786_),
    .B2(_06564_),
    .C1(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__o21ai_1 _09875_ (.A1(_02784_),
    .A2(_02785_),
    .B1(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__a221o_1 _09876_ (.A1(_02771_),
    .A2(_02778_),
    .B1(_02780_),
    .B2(_02443_),
    .C1(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__o41a_2 _09877_ (.A1(_02750_),
    .A2(_02752_),
    .A3(_02757_),
    .A4(_02794_),
    .B1(net241),
    .X(_02795_));
 sky130_fd_sc_hd__nand3_2 _09878_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .C(curr_PC[2]),
    .Y(_02796_));
 sky130_fd_sc_hd__a21o_1 _09879_ (.A1(curr_PC[0]),
    .A2(curr_PC[1]),
    .B1(curr_PC[2]),
    .X(_02797_));
 sky130_fd_sc_hd__a31o_4 _09880_ (.A1(net242),
    .A2(_02796_),
    .A3(_02797_),
    .B1(_02795_),
    .X(dest_val[2]));
 sky130_fd_sc_hd__or4b_2 _09881_ (.A(_02241_),
    .B(_02347_),
    .C(_02748_),
    .D_N(_02574_),
    .X(_02798_));
 sky130_fd_sc_hd__a21oi_4 _09882_ (.A1(_02643_),
    .A2(_02739_),
    .B1(_02738_),
    .Y(_02799_));
 sky130_fd_sc_hd__a21bo_2 _09883_ (.A1(_02728_),
    .A2(_02734_),
    .B1_N(_02736_),
    .X(_02800_));
 sky130_fd_sc_hd__a31oi_4 _09884_ (.A1(_02682_),
    .A2(_02683_),
    .A3(_02703_),
    .B1(_02702_),
    .Y(_02801_));
 sky130_fd_sc_hd__o22a_1 _09885_ (.A1(net33),
    .A2(_00371_),
    .B1(net110),
    .B2(net35),
    .X(_02802_));
 sky130_fd_sc_hd__xnor2_1 _09886_ (.A(net95),
    .B(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__inv_2 _09887_ (.A(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__a22o_1 _09888_ (.A1(net112),
    .A2(net17),
    .B1(net13),
    .B2(net107),
    .X(_02805_));
 sky130_fd_sc_hd__xnor2_1 _09889_ (.A(net65),
    .B(_02805_),
    .Y(_02806_));
 sky130_fd_sc_hd__a22o_1 _09890_ (.A1(net14),
    .A2(_00375_),
    .B1(_00392_),
    .B2(net30),
    .X(_02807_));
 sky130_fd_sc_hd__xnor2_1 _09891_ (.A(net91),
    .B(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _09892_ (.A(_02806_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__xnor2_1 _09893_ (.A(_02806_),
    .B(_02808_),
    .Y(_02810_));
 sky130_fd_sc_hd__xnor2_1 _09894_ (.A(_02804_),
    .B(_02810_),
    .Y(_02811_));
 sky130_fd_sc_hd__a21oi_1 _09895_ (.A1(_02662_),
    .A2(_02664_),
    .B1(_02811_),
    .Y(_02812_));
 sky130_fd_sc_hd__and3_1 _09896_ (.A(_02662_),
    .B(_02664_),
    .C(_02811_),
    .X(_02813_));
 sky130_fd_sc_hd__nor2_2 _09897_ (.A(_02812_),
    .B(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__xnor2_4 _09898_ (.A(_02801_),
    .B(_02814_),
    .Y(_02815_));
 sky130_fd_sc_hd__a21bo_1 _09899_ (.A1(_02646_),
    .A2(_02653_),
    .B1_N(_02651_),
    .X(_02816_));
 sky130_fd_sc_hd__o22a_1 _09900_ (.A1(net21),
    .A2(net77),
    .B1(net74),
    .B2(net18),
    .X(_02817_));
 sky130_fd_sc_hd__xnor2_1 _09901_ (.A(net96),
    .B(_02817_),
    .Y(_02818_));
 sky130_fd_sc_hd__o22a_1 _09902_ (.A1(net103),
    .A2(net27),
    .B1(net70),
    .B2(net29),
    .X(_02819_));
 sky130_fd_sc_hd__xnor2_1 _09903_ (.A(net90),
    .B(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__o22a_1 _09904_ (.A1(net38),
    .A2(_00398_),
    .B1(_00442_),
    .B2(net36),
    .X(_02821_));
 sky130_fd_sc_hd__xnor2_1 _09905_ (.A(net99),
    .B(_02821_),
    .Y(_02822_));
 sky130_fd_sc_hd__nand2_1 _09906_ (.A(_02820_),
    .B(_02822_),
    .Y(_02823_));
 sky130_fd_sc_hd__or2_1 _09907_ (.A(_02820_),
    .B(_02822_),
    .X(_02824_));
 sky130_fd_sc_hd__nand2_1 _09908_ (.A(_02823_),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__xnor2_1 _09909_ (.A(_02818_),
    .B(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__a31o_1 _09910_ (.A1(net150),
    .A2(net63),
    .A3(_02671_),
    .B1(_02670_),
    .X(_02827_));
 sky130_fd_sc_hd__nand2_1 _09911_ (.A(_02826_),
    .B(_02827_),
    .Y(_02828_));
 sky130_fd_sc_hd__xnor2_1 _09912_ (.A(_02826_),
    .B(_02827_),
    .Y(_02829_));
 sky130_fd_sc_hd__nand2b_1 _09913_ (.A_N(_02829_),
    .B(_02816_),
    .Y(_02830_));
 sky130_fd_sc_hd__xnor2_1 _09914_ (.A(_02816_),
    .B(_02829_),
    .Y(_02831_));
 sky130_fd_sc_hd__a21o_1 _09915_ (.A1(_02686_),
    .A2(_02692_),
    .B1(_02691_),
    .X(_02832_));
 sky130_fd_sc_hd__o21ai_1 _09916_ (.A1(_02675_),
    .A2(_02681_),
    .B1(_02680_),
    .Y(_02833_));
 sky130_fd_sc_hd__a21o_1 _09917_ (.A1(_02710_),
    .A2(_02716_),
    .B1(_02715_),
    .X(_02834_));
 sky130_fd_sc_hd__nand2_1 _09918_ (.A(_02833_),
    .B(_02834_),
    .Y(_02835_));
 sky130_fd_sc_hd__xor2_1 _09919_ (.A(_02833_),
    .B(_02834_),
    .X(_02836_));
 sky130_fd_sc_hd__and2_1 _09920_ (.A(_02832_),
    .B(_02836_),
    .X(_02837_));
 sky130_fd_sc_hd__nand2_1 _09921_ (.A(_02832_),
    .B(_02836_),
    .Y(_02838_));
 sky130_fd_sc_hd__nor2_1 _09922_ (.A(_02832_),
    .B(_02836_),
    .Y(_02839_));
 sky130_fd_sc_hd__nor2_1 _09923_ (.A(_02837_),
    .B(_02839_),
    .Y(_02840_));
 sky130_fd_sc_hd__a22o_1 _09924_ (.A1(_00136_),
    .A2(net129),
    .B1(net127),
    .B2(_00177_),
    .X(_02841_));
 sky130_fd_sc_hd__xnor2_2 _09925_ (.A(net155),
    .B(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__o22a_1 _09926_ (.A1(net45),
    .A2(net68),
    .B1(net66),
    .B2(net49),
    .X(_02843_));
 sky130_fd_sc_hd__xnor2_1 _09927_ (.A(net145),
    .B(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__nand2_1 _09928_ (.A(_00197_),
    .B(_00516_),
    .Y(_02845_));
 sky130_fd_sc_hd__nand2_1 _09929_ (.A(_00204_),
    .B(_00812_),
    .Y(_02846_));
 sky130_fd_sc_hd__a21o_1 _09930_ (.A1(_02845_),
    .A2(_02846_),
    .B1(_00188_),
    .X(_02847_));
 sky130_fd_sc_hd__nand3_1 _09931_ (.A(_00188_),
    .B(_02845_),
    .C(_02846_),
    .Y(_02848_));
 sky130_fd_sc_hd__and3_1 _09932_ (.A(_02844_),
    .B(_02847_),
    .C(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__a21oi_1 _09933_ (.A1(_02847_),
    .A2(_02848_),
    .B1(_02844_),
    .Y(_02850_));
 sky130_fd_sc_hd__or2_1 _09934_ (.A(_02849_),
    .B(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__xnor2_2 _09935_ (.A(_02842_),
    .B(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__o22a_1 _09936_ (.A1(net40),
    .A2(net83),
    .B1(net79),
    .B2(net56),
    .X(_02853_));
 sky130_fd_sc_hd__xnor2_1 _09937_ (.A(net117),
    .B(_02853_),
    .Y(_02854_));
 sky130_fd_sc_hd__inv_2 _09938_ (.A(_02854_),
    .Y(_02855_));
 sky130_fd_sc_hd__o22a_1 _09939_ (.A1(net100),
    .A2(net25),
    .B1(net23),
    .B2(net42),
    .X(_02856_));
 sky130_fd_sc_hd__xnor2_1 _09940_ (.A(net86),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__o22a_1 _09941_ (.A1(net53),
    .A2(net75),
    .B1(net72),
    .B2(net47),
    .X(_02858_));
 sky130_fd_sc_hd__xnor2_1 _09942_ (.A(net109),
    .B(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__nand2_1 _09943_ (.A(_02857_),
    .B(_02859_),
    .Y(_02860_));
 sky130_fd_sc_hd__or2_1 _09944_ (.A(_02857_),
    .B(_02859_),
    .X(_02861_));
 sky130_fd_sc_hd__nand2_1 _09945_ (.A(_02860_),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__xnor2_1 _09946_ (.A(_02855_),
    .B(_02862_),
    .Y(_02863_));
 sky130_fd_sc_hd__a22o_1 _09947_ (.A1(_06702_),
    .A2(net11),
    .B1(net6),
    .B2(_06726_),
    .X(_02864_));
 sky130_fd_sc_hd__xnor2_2 _09948_ (.A(net181),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__nand2_1 _09949_ (.A(net198),
    .B(_02865_),
    .Y(_02866_));
 sky130_fd_sc_hd__xnor2_2 _09950_ (.A(net199),
    .B(_02865_),
    .Y(_02867_));
 sky130_fd_sc_hd__xnor2_2 _09951_ (.A(net202),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__or2_1 _09952_ (.A(_02863_),
    .B(_02868_),
    .X(_02869_));
 sky130_fd_sc_hd__xnor2_1 _09953_ (.A(_02863_),
    .B(_02868_),
    .Y(_02870_));
 sky130_fd_sc_hd__xor2_1 _09954_ (.A(_02852_),
    .B(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__nand2_1 _09955_ (.A(net148),
    .B(net63),
    .Y(_02872_));
 sky130_fd_sc_hd__a21oi_2 _09956_ (.A1(_02698_),
    .A2(_02700_),
    .B1(_02697_),
    .Y(_02873_));
 sky130_fd_sc_hd__a22o_1 _09957_ (.A1(_00287_),
    .A2(net9),
    .B1(net4),
    .B2(_00266_),
    .X(_02874_));
 sky130_fd_sc_hd__xnor2_1 _09958_ (.A(net60),
    .B(_02874_),
    .Y(_02875_));
 sky130_fd_sc_hd__and2b_1 _09959_ (.A_N(_02873_),
    .B(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__xnor2_1 _09960_ (.A(_02873_),
    .B(_02875_),
    .Y(_02877_));
 sky130_fd_sc_hd__xnor2_1 _09961_ (.A(_02872_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__nand2_1 _09962_ (.A(_02871_),
    .B(_02878_),
    .Y(_02879_));
 sky130_fd_sc_hd__xnor2_1 _09963_ (.A(_02871_),
    .B(_02878_),
    .Y(_02880_));
 sky130_fd_sc_hd__xnor2_1 _09964_ (.A(_02840_),
    .B(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__and2_1 _09965_ (.A(_02831_),
    .B(_02881_),
    .X(_02882_));
 sky130_fd_sc_hd__nor2_1 _09966_ (.A(_02831_),
    .B(_02881_),
    .Y(_02883_));
 sky130_fd_sc_hd__nor2_2 _09967_ (.A(_02882_),
    .B(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__xor2_4 _09968_ (.A(_02815_),
    .B(_02884_),
    .X(_02885_));
 sky130_fd_sc_hd__a21o_1 _09969_ (.A1(_02658_),
    .A2(_02725_),
    .B1(_02723_),
    .X(_02886_));
 sky130_fd_sc_hd__o21ai_4 _09970_ (.A1(_02654_),
    .A2(_02655_),
    .B1(_02657_),
    .Y(_02887_));
 sky130_fd_sc_hd__o21a_2 _09971_ (.A1(_02665_),
    .A2(_02706_),
    .B1(_02705_),
    .X(_02888_));
 sky130_fd_sc_hd__a21o_1 _09972_ (.A1(_02718_),
    .A2(_02719_),
    .B1(_02721_),
    .X(_02889_));
 sky130_fd_sc_hd__and2b_1 _09973_ (.A_N(_02888_),
    .B(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__xnor2_4 _09974_ (.A(_02888_),
    .B(_02889_),
    .Y(_02891_));
 sky130_fd_sc_hd__xnor2_4 _09975_ (.A(_02887_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__a21oi_4 _09976_ (.A1(_02729_),
    .A2(_02733_),
    .B1(_02732_),
    .Y(_02893_));
 sky130_fd_sc_hd__xnor2_2 _09977_ (.A(_02892_),
    .B(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__nand2b_1 _09978_ (.A_N(_02894_),
    .B(_02886_),
    .Y(_02895_));
 sky130_fd_sc_hd__xnor2_2 _09979_ (.A(_02886_),
    .B(_02894_),
    .Y(_02896_));
 sky130_fd_sc_hd__and2_1 _09980_ (.A(_02885_),
    .B(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__xor2_4 _09981_ (.A(_02885_),
    .B(_02896_),
    .X(_02898_));
 sky130_fd_sc_hd__xnor2_4 _09982_ (.A(_02800_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__or2_2 _09983_ (.A(_02799_),
    .B(_02899_),
    .X(_02900_));
 sky130_fd_sc_hd__and2_1 _09984_ (.A(_02799_),
    .B(_02899_),
    .X(_02901_));
 sky130_fd_sc_hd__xnor2_4 _09985_ (.A(_02799_),
    .B(_02899_),
    .Y(_02902_));
 sky130_fd_sc_hd__or4_1 _09986_ (.A(_02233_),
    .B(_02346_),
    .C(_02569_),
    .D(_02742_),
    .X(_02903_));
 sky130_fd_sc_hd__o22ai_1 _09987_ (.A1(_02464_),
    .A2(_02568_),
    .B1(_02642_),
    .B2(_02740_),
    .Y(_02904_));
 sky130_fd_sc_hd__a21bo_1 _09988_ (.A1(_02642_),
    .A2(_02740_),
    .B1_N(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__or4_1 _09989_ (.A(_02345_),
    .B(_02569_),
    .C(_02571_),
    .D(_02742_),
    .X(_02906_));
 sky130_fd_sc_hd__o211a_2 _09990_ (.A1(_02239_),
    .A2(_02903_),
    .B1(_02905_),
    .C1(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__xor2_4 _09991_ (.A(_02902_),
    .B(_02907_),
    .X(_02908_));
 sky130_fd_sc_hd__a21oi_1 _09992_ (.A1(net137),
    .A2(_02798_),
    .B1(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__a31o_1 _09993_ (.A1(net137),
    .A2(_02798_),
    .A3(_02908_),
    .B1(net235),
    .X(_02910_));
 sky130_fd_sc_hd__and3_1 _09994_ (.A(net137),
    .B(_01926_),
    .C(_01928_),
    .X(_02911_));
 sky130_fd_sc_hd__a21oi_1 _09995_ (.A1(net137),
    .A2(_01926_),
    .B1(_01928_),
    .Y(_02912_));
 sky130_fd_sc_hd__nor2_1 _09996_ (.A(_02911_),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__mux2_1 _09997_ (.A0(_02583_),
    .A1(_02586_),
    .S(_06569_),
    .X(_02914_));
 sky130_fd_sc_hd__mux2_1 _09998_ (.A0(_02585_),
    .A1(_02593_),
    .S(_06569_),
    .X(_02915_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(_02914_),
    .A1(_02915_),
    .S(net215),
    .X(_02916_));
 sky130_fd_sc_hd__mux2_1 _10000_ (.A0(_02589_),
    .A1(_02601_),
    .S(_06569_),
    .X(_02917_));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(_02590_),
    .A1(_02592_),
    .S(net213),
    .X(_02918_));
 sky130_fd_sc_hd__mux2_1 _10002_ (.A0(_02917_),
    .A1(_02918_),
    .S(net217),
    .X(_02919_));
 sky130_fd_sc_hd__mux2_1 _10003_ (.A0(_02916_),
    .A1(_02919_),
    .S(net218),
    .X(_02920_));
 sky130_fd_sc_hd__mux2_1 _10004_ (.A0(_02597_),
    .A1(_02607_),
    .S(_06569_),
    .X(_02921_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(_02598_),
    .A1(_02600_),
    .S(net213),
    .X(_02922_));
 sky130_fd_sc_hd__mux2_1 _10006_ (.A0(_02921_),
    .A1(_02922_),
    .S(net217),
    .X(_02923_));
 sky130_fd_sc_hd__mux2_1 _10007_ (.A0(_02604_),
    .A1(_02606_),
    .S(net214),
    .X(_02924_));
 sky130_fd_sc_hd__mux2_1 _10008_ (.A0(_02451_),
    .A1(_02924_),
    .S(net217),
    .X(_02925_));
 sky130_fd_sc_hd__mux2_1 _10009_ (.A0(_02923_),
    .A1(_02925_),
    .S(net219),
    .X(_02926_));
 sky130_fd_sc_hd__mux2_2 _10010_ (.A0(_02920_),
    .A1(_02926_),
    .S(net221),
    .X(_02927_));
 sky130_fd_sc_hd__o21a_1 _10011_ (.A1(_02772_),
    .A2(_02773_),
    .B1(_02774_),
    .X(_02928_));
 sky130_fd_sc_hd__nor2_1 _10012_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02929_));
 sky130_fd_sc_hd__or2_1 _10013_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .X(_02930_));
 sky130_fd_sc_hd__nand2_1 _10014_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02931_));
 sky130_fd_sc_hd__a21oi_1 _10015_ (.A1(_02930_),
    .A2(_02931_),
    .B1(_02928_),
    .Y(_02932_));
 sky130_fd_sc_hd__and3_1 _10016_ (.A(_02928_),
    .B(_02930_),
    .C(_02931_),
    .X(_02933_));
 sky130_fd_sc_hd__or3_1 _10017_ (.A(net223),
    .B(_02932_),
    .C(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__o211a_1 _10018_ (.A1(net244),
    .A2(_02927_),
    .B1(_02934_),
    .C1(net205),
    .X(_02935_));
 sky130_fd_sc_hd__o21a_1 _10019_ (.A1(net216),
    .A2(_02408_),
    .B1(_02452_),
    .X(_02936_));
 sky130_fd_sc_hd__o21a_1 _10020_ (.A1(net219),
    .A2(_02936_),
    .B1(_02453_),
    .X(_02937_));
 sky130_fd_sc_hd__o21ai_2 _10021_ (.A1(net221),
    .A2(_02937_),
    .B1(_02456_),
    .Y(_02938_));
 sky130_fd_sc_hd__inv_2 _10022_ (.A(_02938_),
    .Y(_02939_));
 sky130_fd_sc_hd__a22o_1 _10023_ (.A1(net167),
    .A2(_02927_),
    .B1(_02939_),
    .B2(net172),
    .X(_02940_));
 sky130_fd_sc_hd__a211oi_1 _10024_ (.A1(_06563_),
    .A2(_02781_),
    .B1(_06564_),
    .C1(net295),
    .Y(_02941_));
 sky130_fd_sc_hd__a31oi_1 _10025_ (.A1(net295),
    .A2(_06562_),
    .A3(_06580_),
    .B1(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__xnor2_1 _10026_ (.A(_06558_),
    .B(_02942_),
    .Y(_02943_));
 sky130_fd_sc_hd__or3_1 _10027_ (.A(\div_res[2] ),
    .B(\div_res[1] ),
    .C(\div_res[0] ),
    .X(_02944_));
 sky130_fd_sc_hd__a21oi_1 _10028_ (.A1(net140),
    .A2(_02944_),
    .B1(\div_res[3] ),
    .Y(_02945_));
 sky130_fd_sc_hd__a31o_1 _10029_ (.A1(\div_res[3] ),
    .A2(net139),
    .A3(_02944_),
    .B1(net189),
    .X(_02946_));
 sky130_fd_sc_hd__a21oi_1 _10030_ (.A1(_06557_),
    .A2(net195),
    .B1(net193),
    .Y(_02947_));
 sky130_fd_sc_hd__or3_1 _10031_ (.A(\div_shifter[34] ),
    .B(\div_shifter[33] ),
    .C(\div_shifter[32] ),
    .X(_02948_));
 sky130_fd_sc_hd__a21oi_1 _10032_ (.A1(net230),
    .A2(_02948_),
    .B1(\div_shifter[35] ),
    .Y(_02949_));
 sky130_fd_sc_hd__a31o_1 _10033_ (.A1(\div_shifter[35] ),
    .A2(net230),
    .A3(_02948_),
    .B1(net192),
    .X(_02950_));
 sky130_fd_sc_hd__o2bb2a_1 _10034_ (.A1_N(_06691_),
    .A2_N(net256),
    .B1(net231),
    .B2(reg1_val[3]),
    .X(_02951_));
 sky130_fd_sc_hd__o221a_1 _10035_ (.A1(_06553_),
    .A2(net203),
    .B1(_02949_),
    .B2(_02950_),
    .C1(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__o221a_1 _10036_ (.A1(_06557_),
    .A2(net194),
    .B1(_02947_),
    .B2(_06556_),
    .C1(_02952_),
    .X(_02953_));
 sky130_fd_sc_hd__o21ai_1 _10037_ (.A1(_02945_),
    .A2(_02946_),
    .B1(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__a211o_1 _10038_ (.A1(net234),
    .A2(_02943_),
    .B1(_02954_),
    .C1(_02935_),
    .X(_02955_));
 sky130_fd_sc_hd__a211o_1 _10039_ (.A1(net233),
    .A2(_02913_),
    .B1(_02940_),
    .C1(_02955_),
    .X(_02956_));
 sky130_fd_sc_hd__o21bai_2 _10040_ (.A1(_02909_),
    .A2(_02910_),
    .B1_N(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__nor2_2 _10041_ (.A(_04620_),
    .B(_02796_),
    .Y(_02958_));
 sky130_fd_sc_hd__a21o_1 _10042_ (.A1(_04620_),
    .A2(_02796_),
    .B1(net237),
    .X(_02959_));
 sky130_fd_sc_hd__a2bb2o_4 _10043_ (.A1_N(_02958_),
    .A2_N(_02959_),
    .B1(net237),
    .B2(_02957_),
    .X(dest_val[3]));
 sky130_fd_sc_hd__nor2_1 _10044_ (.A(_02798_),
    .B(_02908_),
    .Y(_02960_));
 sky130_fd_sc_hd__or2_1 _10045_ (.A(net135),
    .B(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__a21oi_4 _10046_ (.A1(_02800_),
    .A2(_02898_),
    .B1(_02897_),
    .Y(_02962_));
 sky130_fd_sc_hd__o21ai_4 _10047_ (.A1(_02892_),
    .A2(_02893_),
    .B1(_02895_),
    .Y(_02963_));
 sky130_fd_sc_hd__o21a_2 _10048_ (.A1(_02852_),
    .A2(_02870_),
    .B1(_02869_),
    .X(_02964_));
 sky130_fd_sc_hd__o22a_1 _10049_ (.A1(net35),
    .A2(net123),
    .B1(net120),
    .B2(net33),
    .X(_02965_));
 sky130_fd_sc_hd__xnor2_1 _10050_ (.A(net95),
    .B(_02965_),
    .Y(_02966_));
 sky130_fd_sc_hd__inv_2 _10051_ (.A(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__a22o_1 _10052_ (.A1(net111),
    .A2(net17),
    .B1(net13),
    .B2(net112),
    .X(_02968_));
 sky130_fd_sc_hd__xnor2_1 _10053_ (.A(net65),
    .B(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__a22o_1 _10054_ (.A1(net14),
    .A2(_00392_),
    .B1(_00397_),
    .B2(net30),
    .X(_02970_));
 sky130_fd_sc_hd__xnor2_1 _10055_ (.A(net91),
    .B(_02970_),
    .Y(_02971_));
 sky130_fd_sc_hd__nand2_1 _10056_ (.A(_02969_),
    .B(_02971_),
    .Y(_02972_));
 sky130_fd_sc_hd__xnor2_1 _10057_ (.A(_02969_),
    .B(_02971_),
    .Y(_02973_));
 sky130_fd_sc_hd__xnor2_1 _10058_ (.A(_02967_),
    .B(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__a21oi_1 _10059_ (.A1(_02835_),
    .A2(_02838_),
    .B1(_02974_),
    .Y(_02975_));
 sky130_fd_sc_hd__and3_1 _10060_ (.A(_02835_),
    .B(_02838_),
    .C(_02974_),
    .X(_02976_));
 sky130_fd_sc_hd__nor2_2 _10061_ (.A(_02975_),
    .B(_02976_),
    .Y(_02977_));
 sky130_fd_sc_hd__and2b_1 _10062_ (.A_N(_02964_),
    .B(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__xnor2_4 _10063_ (.A(_02964_),
    .B(_02977_),
    .Y(_02979_));
 sky130_fd_sc_hd__o21ai_1 _10064_ (.A1(_02855_),
    .A2(_02862_),
    .B1(_02860_),
    .Y(_02980_));
 sky130_fd_sc_hd__a21bo_1 _10065_ (.A1(_02818_),
    .A2(_02824_),
    .B1_N(_02823_),
    .X(_02981_));
 sky130_fd_sc_hd__o21bai_2 _10066_ (.A1(_02842_),
    .A2(_02850_),
    .B1_N(_02849_),
    .Y(_02982_));
 sky130_fd_sc_hd__nand2_1 _10067_ (.A(_02981_),
    .B(_02982_),
    .Y(_02983_));
 sky130_fd_sc_hd__xor2_1 _10068_ (.A(_02981_),
    .B(_02982_),
    .X(_02984_));
 sky130_fd_sc_hd__nand2_2 _10069_ (.A(_02980_),
    .B(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__or2_1 _10070_ (.A(_02980_),
    .B(_02984_),
    .X(_02986_));
 sky130_fd_sc_hd__nand2_4 _10071_ (.A(_02985_),
    .B(_02986_),
    .Y(_02987_));
 sky130_fd_sc_hd__o22a_1 _10072_ (.A1(net49),
    .A2(net68),
    .B1(net66),
    .B2(net51),
    .X(_02988_));
 sky130_fd_sc_hd__xnor2_1 _10073_ (.A(net145),
    .B(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__inv_2 _10074_ (.A(_02989_),
    .Y(_02990_));
 sky130_fd_sc_hd__o22a_1 _10075_ (.A1(net47),
    .A2(net75),
    .B1(net72),
    .B2(net45),
    .X(_02991_));
 sky130_fd_sc_hd__xnor2_1 _10076_ (.A(net108),
    .B(_02991_),
    .Y(_02992_));
 sky130_fd_sc_hd__o32a_1 _10077_ (.A1(_00232_),
    .A2(_00513_),
    .A3(_00515_),
    .B1(_00227_),
    .B2(net44),
    .X(_02993_));
 sky130_fd_sc_hd__xnor2_1 _10078_ (.A(net154),
    .B(_02993_),
    .Y(_02994_));
 sky130_fd_sc_hd__nand2_1 _10079_ (.A(_02992_),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__or2_1 _10080_ (.A(_02992_),
    .B(_02994_),
    .X(_02996_));
 sky130_fd_sc_hd__nand2_1 _10081_ (.A(_02995_),
    .B(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__xnor2_1 _10082_ (.A(_02990_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__o22a_1 _10083_ (.A1(net42),
    .A2(net25),
    .B1(net23),
    .B2(net40),
    .X(_02999_));
 sky130_fd_sc_hd__xnor2_1 _10084_ (.A(net87),
    .B(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__inv_2 _10085_ (.A(_03000_),
    .Y(_03001_));
 sky130_fd_sc_hd__o22a_1 _10086_ (.A1(net103),
    .A2(net29),
    .B1(net27),
    .B2(_00230_),
    .X(_03002_));
 sky130_fd_sc_hd__xnor2_2 _10087_ (.A(net89),
    .B(_03002_),
    .Y(_03003_));
 sky130_fd_sc_hd__o22a_1 _10088_ (.A1(net56),
    .A2(net83),
    .B1(net79),
    .B2(net53),
    .X(_03004_));
 sky130_fd_sc_hd__xnor2_2 _10089_ (.A(net117),
    .B(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__and2_1 _10090_ (.A(_03003_),
    .B(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__xnor2_2 _10091_ (.A(_03003_),
    .B(_03005_),
    .Y(_03007_));
 sky130_fd_sc_hd__nor2_1 _10092_ (.A(_03001_),
    .B(_03007_),
    .Y(_03008_));
 sky130_fd_sc_hd__xnor2_2 _10093_ (.A(_03001_),
    .B(_03007_),
    .Y(_03009_));
 sky130_fd_sc_hd__o22a_1 _10094_ (.A1(net105),
    .A2(_00811_),
    .B1(net10),
    .B2(net131),
    .X(_03010_));
 sky130_fd_sc_hd__xnor2_2 _10095_ (.A(net174),
    .B(_03010_),
    .Y(_03011_));
 sky130_fd_sc_hd__nand2_1 _10096_ (.A(_06697_),
    .B(net6),
    .Y(_03012_));
 sky130_fd_sc_hd__a22o_1 _10097_ (.A1(_06700_),
    .A2(net6),
    .B1(_03012_),
    .B2(net179),
    .X(_03013_));
 sky130_fd_sc_hd__nor2_1 _10098_ (.A(_03011_),
    .B(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__xor2_2 _10099_ (.A(_03011_),
    .B(_03013_),
    .X(_03015_));
 sky130_fd_sc_hd__xnor2_1 _10100_ (.A(_03009_),
    .B(_03015_),
    .Y(_03016_));
 sky130_fd_sc_hd__or2_1 _10101_ (.A(_02998_),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__nand2_1 _10102_ (.A(_02998_),
    .B(_03016_),
    .Y(_03018_));
 sky130_fd_sc_hd__and2_2 _10103_ (.A(_03017_),
    .B(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__nand2_2 _10104_ (.A(_00266_),
    .B(net63),
    .Y(_03020_));
 sky130_fd_sc_hd__a21bo_2 _10105_ (.A1(net202),
    .A2(_02867_),
    .B1_N(_02866_),
    .X(_03021_));
 sky130_fd_sc_hd__a22o_1 _10106_ (.A1(net107),
    .A2(net9),
    .B1(net4),
    .B2(_00287_),
    .X(_03022_));
 sky130_fd_sc_hd__xnor2_2 _10107_ (.A(net60),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__and2_1 _10108_ (.A(_03021_),
    .B(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__xor2_4 _10109_ (.A(_03021_),
    .B(_03023_),
    .X(_03025_));
 sky130_fd_sc_hd__xnor2_4 _10110_ (.A(_03020_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__nand2_1 _10111_ (.A(_03019_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__xnor2_4 _10112_ (.A(_03019_),
    .B(_03026_),
    .Y(_03028_));
 sky130_fd_sc_hd__xor2_4 _10113_ (.A(_02987_),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__o21ai_1 _10114_ (.A1(_02804_),
    .A2(_02810_),
    .B1(_02809_),
    .Y(_03030_));
 sky130_fd_sc_hd__inv_2 _10115_ (.A(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__o22a_1 _10116_ (.A1(net20),
    .A2(net74),
    .B1(net70),
    .B2(net18),
    .X(_03032_));
 sky130_fd_sc_hd__xnor2_1 _10117_ (.A(net96),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__o22a_1 _10118_ (.A1(net39),
    .A2(net82),
    .B1(net77),
    .B2(net37),
    .X(_03034_));
 sky130_fd_sc_hd__xnor2_1 _10119_ (.A(net99),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__nand2_2 _10120_ (.A(_03033_),
    .B(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__or2_1 _10121_ (.A(_03033_),
    .B(_03035_),
    .X(_03037_));
 sky130_fd_sc_hd__and2_1 _10122_ (.A(_03036_),
    .B(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__a31o_1 _10123_ (.A1(net148),
    .A2(net63),
    .A3(_02877_),
    .B1(_02876_),
    .X(_03039_));
 sky130_fd_sc_hd__and2_1 _10124_ (.A(_03038_),
    .B(_03039_),
    .X(_03040_));
 sky130_fd_sc_hd__xnor2_1 _10125_ (.A(_03038_),
    .B(_03039_),
    .Y(_03041_));
 sky130_fd_sc_hd__nor2_1 _10126_ (.A(_03031_),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__and2_1 _10127_ (.A(_03031_),
    .B(_03041_),
    .X(_03043_));
 sky130_fd_sc_hd__nor2_2 _10128_ (.A(_03042_),
    .B(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__and2_1 _10129_ (.A(_03029_),
    .B(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__xor2_4 _10130_ (.A(_03029_),
    .B(_03044_),
    .X(_03046_));
 sky130_fd_sc_hd__xor2_4 _10131_ (.A(_02979_),
    .B(_03046_),
    .X(_03047_));
 sky130_fd_sc_hd__a21o_1 _10132_ (.A1(_02815_),
    .A2(_02884_),
    .B1(_02882_),
    .X(_03048_));
 sky130_fd_sc_hd__o21bai_2 _10133_ (.A1(_02801_),
    .A2(_02813_),
    .B1_N(_02812_),
    .Y(_03049_));
 sky130_fd_sc_hd__nand2_1 _10134_ (.A(_02828_),
    .B(_02830_),
    .Y(_03050_));
 sky130_fd_sc_hd__o31a_1 _10135_ (.A1(_02837_),
    .A2(_02839_),
    .A3(_02880_),
    .B1(_02879_),
    .X(_03051_));
 sky130_fd_sc_hd__a21o_1 _10136_ (.A1(_02828_),
    .A2(_02830_),
    .B1(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__xnor2_2 _10137_ (.A(_03050_),
    .B(_03051_),
    .Y(_03053_));
 sky130_fd_sc_hd__xnor2_2 _10138_ (.A(_03049_),
    .B(_03053_),
    .Y(_03054_));
 sky130_fd_sc_hd__a21oi_2 _10139_ (.A1(_02887_),
    .A2(_02891_),
    .B1(_02890_),
    .Y(_03055_));
 sky130_fd_sc_hd__xnor2_1 _10140_ (.A(_03054_),
    .B(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__nand2b_1 _10141_ (.A_N(_03056_),
    .B(_03048_),
    .Y(_03057_));
 sky130_fd_sc_hd__xnor2_2 _10142_ (.A(_03048_),
    .B(_03056_),
    .Y(_03058_));
 sky130_fd_sc_hd__and2_1 _10143_ (.A(_03047_),
    .B(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__xor2_4 _10144_ (.A(_03047_),
    .B(_03058_),
    .X(_03060_));
 sky130_fd_sc_hd__xnor2_4 _10145_ (.A(_02963_),
    .B(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__or2_1 _10146_ (.A(_02962_),
    .B(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__and2_1 _10147_ (.A(_02962_),
    .B(_03061_),
    .X(_03063_));
 sky130_fd_sc_hd__xnor2_4 _10148_ (.A(_02962_),
    .B(_03061_),
    .Y(_03064_));
 sky130_fd_sc_hd__inv_2 _10149_ (.A(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__or4_1 _10150_ (.A(_02346_),
    .B(_02569_),
    .C(_02742_),
    .D(_02902_),
    .X(_03066_));
 sky130_fd_sc_hd__a21o_1 _10151_ (.A1(_02242_),
    .A2(_02244_),
    .B1(_03066_),
    .X(_03067_));
 sky130_fd_sc_hd__a21o_1 _10152_ (.A1(_02741_),
    .A2(_02900_),
    .B1(_02901_),
    .X(_03068_));
 sky130_fd_sc_hd__o31a_1 _10153_ (.A1(_02742_),
    .A2(_02745_),
    .A3(_02902_),
    .B1(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__a21oi_1 _10154_ (.A1(_03067_),
    .A2(_03069_),
    .B1(_03065_),
    .Y(_03070_));
 sky130_fd_sc_hd__and3_1 _10155_ (.A(_03065_),
    .B(_03067_),
    .C(_03069_),
    .X(_03071_));
 sky130_fd_sc_hd__nor2_1 _10156_ (.A(_03070_),
    .B(_03071_),
    .Y(_03072_));
 sky130_fd_sc_hd__o21ai_1 _10157_ (.A1(_02961_),
    .A2(_03072_),
    .B1(_02348_),
    .Y(_03073_));
 sky130_fd_sc_hd__a21oi_1 _10158_ (.A1(_02961_),
    .A2(_03072_),
    .B1(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__o21ai_1 _10159_ (.A1(net134),
    .A2(_01929_),
    .B1(_01930_),
    .Y(_03075_));
 sky130_fd_sc_hd__or3_1 _10160_ (.A(net134),
    .B(_01929_),
    .C(_01930_),
    .X(_03076_));
 sky130_fd_sc_hd__a211o_1 _10161_ (.A1(_06563_),
    .A2(_02781_),
    .B1(_06564_),
    .C1(_06556_),
    .X(_03077_));
 sky130_fd_sc_hd__a21oi_1 _10162_ (.A1(_06557_),
    .A2(_03077_),
    .B1(net295),
    .Y(_03078_));
 sky130_fd_sc_hd__a31o_1 _10163_ (.A1(net295),
    .A2(_06555_),
    .A3(_06581_),
    .B1(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__nand2_1 _10164_ (.A(_06551_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__or2_1 _10165_ (.A(_06551_),
    .B(_03079_),
    .X(_03081_));
 sky130_fd_sc_hd__o21a_1 _10166_ (.A1(_02928_),
    .A2(_02929_),
    .B1(_02931_),
    .X(_03082_));
 sky130_fd_sc_hd__nor2_1 _10167_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_03083_));
 sky130_fd_sc_hd__nand2_1 _10168_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_03084_));
 sky130_fd_sc_hd__nand2b_1 _10169_ (.A_N(_03083_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__xnor2_1 _10170_ (.A(_03082_),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__mux2_1 _10171_ (.A0(_02369_),
    .A1(_02385_),
    .S(net215),
    .X(_03087_));
 sky130_fd_sc_hd__or2_1 _10172_ (.A(net217),
    .B(_02400_),
    .X(_03088_));
 sky130_fd_sc_hd__o21ai_1 _10173_ (.A1(net215),
    .A2(_02378_),
    .B1(_03088_),
    .Y(_03089_));
 sky130_fd_sc_hd__nand2_1 _10174_ (.A(net218),
    .B(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__o211a_1 _10175_ (.A1(net218),
    .A2(_03087_),
    .B1(_03090_),
    .C1(net220),
    .X(_03091_));
 sky130_fd_sc_hd__or2_1 _10176_ (.A(net217),
    .B(_02415_),
    .X(_03092_));
 sky130_fd_sc_hd__o21ai_1 _10177_ (.A1(net215),
    .A2(_02393_),
    .B1(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__inv_2 _10178_ (.A(_03093_),
    .Y(_03094_));
 sky130_fd_sc_hd__mux2_1 _10179_ (.A0(_02936_),
    .A1(_03094_),
    .S(_06553_),
    .X(_03095_));
 sky130_fd_sc_hd__a21oi_2 _10180_ (.A1(net221),
    .A2(_03095_),
    .B1(_03091_),
    .Y(_03096_));
 sky130_fd_sc_hd__mux2_1 _10181_ (.A0(_03086_),
    .A1(_03096_),
    .S(net223),
    .X(_03097_));
 sky130_fd_sc_hd__or4_2 _10182_ (.A(\div_res[3] ),
    .B(\div_res[2] ),
    .C(\div_res[1] ),
    .D(\div_res[0] ),
    .X(_03098_));
 sky130_fd_sc_hd__a21oi_1 _10183_ (.A1(net140),
    .A2(_03098_),
    .B1(\div_res[4] ),
    .Y(_03099_));
 sky130_fd_sc_hd__a311o_1 _10184_ (.A1(\div_res[4] ),
    .A2(net140),
    .A3(_03098_),
    .B1(_03099_),
    .C1(net189),
    .X(_03100_));
 sky130_fd_sc_hd__a21oi_1 _10185_ (.A1(_06550_),
    .A2(net195),
    .B1(net193),
    .Y(_03101_));
 sky130_fd_sc_hd__or4_2 _10186_ (.A(\div_shifter[35] ),
    .B(\div_shifter[34] ),
    .C(\div_shifter[33] ),
    .D(\div_shifter[32] ),
    .X(_03102_));
 sky130_fd_sc_hd__a21oi_1 _10187_ (.A1(net230),
    .A2(_03102_),
    .B1(\div_shifter[36] ),
    .Y(_03103_));
 sky130_fd_sc_hd__a31o_1 _10188_ (.A1(\div_shifter[36] ),
    .A2(net230),
    .A3(_03102_),
    .B1(net191),
    .X(_03104_));
 sky130_fd_sc_hd__o2bb2a_1 _10189_ (.A1_N(_06695_),
    .A2_N(net256),
    .B1(net231),
    .B2(reg1_val[4]),
    .X(_03105_));
 sky130_fd_sc_hd__o221a_1 _10190_ (.A1(_06547_),
    .A2(net203),
    .B1(_03103_),
    .B2(_03104_),
    .C1(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__o221a_1 _10191_ (.A1(_06550_),
    .A2(net194),
    .B1(_03101_),
    .B2(_06549_),
    .C1(_03106_),
    .X(_03107_));
 sky130_fd_sc_hd__o21a_1 _10192_ (.A1(net219),
    .A2(_02925_),
    .B1(_02453_),
    .X(_03108_));
 sky130_fd_sc_hd__o21ai_2 _10193_ (.A1(net221),
    .A2(_03108_),
    .B1(_02456_),
    .Y(_03109_));
 sky130_fd_sc_hd__o211a_1 _10194_ (.A1(net169),
    .A2(_03109_),
    .B1(_03107_),
    .C1(_03100_),
    .X(_03110_));
 sky130_fd_sc_hd__o221ai_2 _10195_ (.A1(_02425_),
    .A2(_03096_),
    .B1(_03097_),
    .B2(_06667_),
    .C1(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__a31o_1 _10196_ (.A1(net234),
    .A2(_03080_),
    .A3(_03081_),
    .B1(_03111_),
    .X(_03112_));
 sky130_fd_sc_hd__a311o_1 _10197_ (.A1(net233),
    .A2(_03075_),
    .A3(_03076_),
    .B1(_03112_),
    .C1(_03074_),
    .X(_03113_));
 sky130_fd_sc_hd__xor2_1 _10198_ (.A(curr_PC[4]),
    .B(_02958_),
    .X(_03114_));
 sky130_fd_sc_hd__mux2_8 _10199_ (.A0(_03113_),
    .A1(_03114_),
    .S(net242),
    .X(dest_val[4]));
 sky130_fd_sc_hd__nand2_1 _10200_ (.A(_02960_),
    .B(_03072_),
    .Y(_03115_));
 sky130_fd_sc_hd__and2_1 _10201_ (.A(net137),
    .B(_03115_),
    .X(_03116_));
 sky130_fd_sc_hd__a21oi_4 _10202_ (.A1(_02963_),
    .A2(_03060_),
    .B1(_03059_),
    .Y(_03117_));
 sky130_fd_sc_hd__o21ai_4 _10203_ (.A1(_03054_),
    .A2(_03055_),
    .B1(_03057_),
    .Y(_03118_));
 sky130_fd_sc_hd__o21ai_4 _10204_ (.A1(_03009_),
    .A2(_03015_),
    .B1(_03017_),
    .Y(_03119_));
 sky130_fd_sc_hd__a22o_1 _10205_ (.A1(net14),
    .A2(_00397_),
    .B1(_00443_),
    .B2(net30),
    .X(_03120_));
 sky130_fd_sc_hd__xnor2_1 _10206_ (.A(net91),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__o22a_1 _10207_ (.A1(net34),
    .A2(net120),
    .B1(_00391_),
    .B2(net32),
    .X(_03122_));
 sky130_fd_sc_hd__xnor2_1 _10208_ (.A(net94),
    .B(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__o22a_1 _10209_ (.A1(net39),
    .A2(net77),
    .B1(net74),
    .B2(net36),
    .X(_03124_));
 sky130_fd_sc_hd__xnor2_1 _10210_ (.A(net98),
    .B(_03124_),
    .Y(_03125_));
 sky130_fd_sc_hd__and2_1 _10211_ (.A(_03123_),
    .B(_03125_),
    .X(_03126_));
 sky130_fd_sc_hd__nor2_1 _10212_ (.A(_03123_),
    .B(_03125_),
    .Y(_03127_));
 sky130_fd_sc_hd__or2_1 _10213_ (.A(_03126_),
    .B(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__inv_2 _10214_ (.A(_03128_),
    .Y(_03129_));
 sky130_fd_sc_hd__xor2_1 _10215_ (.A(_03121_),
    .B(_03128_),
    .X(_03130_));
 sky130_fd_sc_hd__a21oi_1 _10216_ (.A1(_02983_),
    .A2(_02985_),
    .B1(_03130_),
    .Y(_03131_));
 sky130_fd_sc_hd__and3_1 _10217_ (.A(_02983_),
    .B(_02985_),
    .C(_03130_),
    .X(_03132_));
 sky130_fd_sc_hd__nor2_2 _10218_ (.A(_03131_),
    .B(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__xor2_4 _10219_ (.A(_03119_),
    .B(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__o21ai_4 _10220_ (.A1(_02990_),
    .A2(_02997_),
    .B1(_02995_),
    .Y(_03135_));
 sky130_fd_sc_hd__o21ba_1 _10221_ (.A1(_03006_),
    .A2(_03008_),
    .B1_N(_03014_),
    .X(_03136_));
 sky130_fd_sc_hd__or3b_2 _10222_ (.A(_03006_),
    .B(_03008_),
    .C_N(_03014_),
    .X(_03137_));
 sky130_fd_sc_hd__nand2b_1 _10223_ (.A_N(_03136_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__xnor2_2 _10224_ (.A(_03135_),
    .B(_03138_),
    .Y(_03139_));
 sky130_fd_sc_hd__nand2_1 _10225_ (.A(_00287_),
    .B(net63),
    .Y(_03140_));
 sky130_fd_sc_hd__o2bb2a_1 _10226_ (.A1_N(net122),
    .A2_N(net16),
    .B1(_00797_),
    .B2(_00415_),
    .X(_03141_));
 sky130_fd_sc_hd__xnor2_1 _10227_ (.A(_00787_),
    .B(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__nand2b_1 _10228_ (.A_N(_03140_),
    .B(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__xnor2_1 _10229_ (.A(_03140_),
    .B(_03142_),
    .Y(_03144_));
 sky130_fd_sc_hd__a22o_1 _10230_ (.A1(net112),
    .A2(net9),
    .B1(net4),
    .B2(net107),
    .X(_03145_));
 sky130_fd_sc_hd__xnor2_1 _10231_ (.A(net59),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__nand2_1 _10232_ (.A(_03144_),
    .B(_03146_),
    .Y(_03147_));
 sky130_fd_sc_hd__or2_1 _10233_ (.A(_03144_),
    .B(_03146_),
    .X(_03148_));
 sky130_fd_sc_hd__nand2_1 _10234_ (.A(_03147_),
    .B(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__o22a_1 _10235_ (.A1(net105),
    .A2(net10),
    .B1(net5),
    .B2(net131),
    .X(_03150_));
 sky130_fd_sc_hd__xnor2_1 _10236_ (.A(net175),
    .B(_03150_),
    .Y(_03151_));
 sky130_fd_sc_hd__a22o_1 _10237_ (.A1(net129),
    .A2(_00516_),
    .B1(_00812_),
    .B2(net127),
    .X(_03152_));
 sky130_fd_sc_hd__xnor2_1 _10238_ (.A(net155),
    .B(_03152_),
    .Y(_03153_));
 sky130_fd_sc_hd__nor2_1 _10239_ (.A(net179),
    .B(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__xnor2_1 _10240_ (.A(_06689_),
    .B(_03153_),
    .Y(_03155_));
 sky130_fd_sc_hd__xnor2_1 _10241_ (.A(_03151_),
    .B(_03155_),
    .Y(_03156_));
 sky130_fd_sc_hd__o22a_1 _10242_ (.A1(net45),
    .A2(net75),
    .B1(net72),
    .B2(net49),
    .X(_03157_));
 sky130_fd_sc_hd__xnor2_1 _10243_ (.A(net108),
    .B(_03157_),
    .Y(_03158_));
 sky130_fd_sc_hd__inv_2 _10244_ (.A(_03158_),
    .Y(_03159_));
 sky130_fd_sc_hd__o22a_1 _10245_ (.A1(net53),
    .A2(net83),
    .B1(net79),
    .B2(net47),
    .X(_03160_));
 sky130_fd_sc_hd__xnor2_2 _10246_ (.A(net117),
    .B(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__o22a_1 _10247_ (.A1(net51),
    .A2(net68),
    .B1(net66),
    .B2(net44),
    .X(_03162_));
 sky130_fd_sc_hd__xnor2_2 _10248_ (.A(net145),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__and2_1 _10249_ (.A(_03161_),
    .B(_03163_),
    .X(_03164_));
 sky130_fd_sc_hd__xnor2_2 _10250_ (.A(_03161_),
    .B(_03163_),
    .Y(_03165_));
 sky130_fd_sc_hd__nor2_1 _10251_ (.A(_03159_),
    .B(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__xnor2_2 _10252_ (.A(_03159_),
    .B(_03165_),
    .Y(_03167_));
 sky130_fd_sc_hd__xor2_1 _10253_ (.A(_03036_),
    .B(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__nand2b_1 _10254_ (.A_N(_03156_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__xor2_1 _10255_ (.A(_03156_),
    .B(_03168_),
    .X(_03170_));
 sky130_fd_sc_hd__nor2_1 _10256_ (.A(_03149_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__nand2_1 _10257_ (.A(_03149_),
    .B(_03170_),
    .Y(_03172_));
 sky130_fd_sc_hd__and2b_1 _10258_ (.A_N(_03171_),
    .B(_03172_),
    .X(_03173_));
 sky130_fd_sc_hd__xor2_1 _10259_ (.A(_03139_),
    .B(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__o21ai_2 _10260_ (.A1(_02967_),
    .A2(_02973_),
    .B1(_02972_),
    .Y(_03175_));
 sky130_fd_sc_hd__inv_2 _10261_ (.A(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__o22a_1 _10262_ (.A1(net100),
    .A2(net29),
    .B1(_00373_),
    .B2(net42),
    .X(_03177_));
 sky130_fd_sc_hd__xnor2_2 _10263_ (.A(net88),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__inv_2 _10264_ (.A(_03178_),
    .Y(_03179_));
 sky130_fd_sc_hd__o22a_1 _10265_ (.A1(net103),
    .A2(net18),
    .B1(net70),
    .B2(net20),
    .X(_03180_));
 sky130_fd_sc_hd__xnor2_1 _10266_ (.A(net96),
    .B(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__o22a_1 _10267_ (.A1(net40),
    .A2(net25),
    .B1(net23),
    .B2(net56),
    .X(_03182_));
 sky130_fd_sc_hd__xnor2_1 _10268_ (.A(net87),
    .B(_03182_),
    .Y(_03183_));
 sky130_fd_sc_hd__nand2_1 _10269_ (.A(_03181_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__xnor2_1 _10270_ (.A(_03181_),
    .B(_03183_),
    .Y(_03185_));
 sky130_fd_sc_hd__xnor2_1 _10271_ (.A(_03178_),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__a31o_1 _10272_ (.A1(_00266_),
    .A2(net63),
    .A3(_03025_),
    .B1(_03024_),
    .X(_03187_));
 sky130_fd_sc_hd__nand2_1 _10273_ (.A(_03186_),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__xnor2_1 _10274_ (.A(_03186_),
    .B(_03187_),
    .Y(_03189_));
 sky130_fd_sc_hd__xnor2_1 _10275_ (.A(_03175_),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__and2_1 _10276_ (.A(_03174_),
    .B(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__nor2_1 _10277_ (.A(_03174_),
    .B(_03190_),
    .Y(_03192_));
 sky130_fd_sc_hd__nor2_2 _10278_ (.A(_03191_),
    .B(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__xor2_4 _10279_ (.A(_03134_),
    .B(_03193_),
    .X(_03194_));
 sky130_fd_sc_hd__a21o_1 _10280_ (.A1(_02979_),
    .A2(_03046_),
    .B1(_03045_),
    .X(_03195_));
 sky130_fd_sc_hd__a21bo_1 _10281_ (.A1(_03049_),
    .A2(_03053_),
    .B1_N(_03052_),
    .X(_03196_));
 sky130_fd_sc_hd__or2_2 _10282_ (.A(_02975_),
    .B(_02978_),
    .X(_03197_));
 sky130_fd_sc_hd__o21ai_4 _10283_ (.A1(_02987_),
    .A2(_03028_),
    .B1(_03027_),
    .Y(_03198_));
 sky130_fd_sc_hd__o21ba_1 _10284_ (.A1(_03031_),
    .A2(_03041_),
    .B1_N(_03040_),
    .X(_03199_));
 sky130_fd_sc_hd__o21ai_1 _10285_ (.A1(_03040_),
    .A2(_03042_),
    .B1(_03198_),
    .Y(_03200_));
 sky130_fd_sc_hd__xnor2_4 _10286_ (.A(_03198_),
    .B(_03199_),
    .Y(_03201_));
 sky130_fd_sc_hd__xor2_2 _10287_ (.A(_03197_),
    .B(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__xnor2_2 _10288_ (.A(_03196_),
    .B(_03202_),
    .Y(_03203_));
 sky130_fd_sc_hd__nand2b_1 _10289_ (.A_N(_03203_),
    .B(_03195_),
    .Y(_03204_));
 sky130_fd_sc_hd__xnor2_2 _10290_ (.A(_03195_),
    .B(_03203_),
    .Y(_03205_));
 sky130_fd_sc_hd__and2_1 _10291_ (.A(_03194_),
    .B(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__xor2_4 _10292_ (.A(_03194_),
    .B(_03205_),
    .X(_03207_));
 sky130_fd_sc_hd__xnor2_4 _10293_ (.A(_03118_),
    .B(_03207_),
    .Y(_03208_));
 sky130_fd_sc_hd__or2_1 _10294_ (.A(_03117_),
    .B(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__and2_1 _10295_ (.A(_03117_),
    .B(_03208_),
    .X(_03210_));
 sky130_fd_sc_hd__xnor2_4 _10296_ (.A(_03117_),
    .B(_03208_),
    .Y(_03211_));
 sky130_fd_sc_hd__or2_1 _10297_ (.A(_02902_),
    .B(_03064_),
    .X(_03212_));
 sky130_fd_sc_hd__or4_1 _10298_ (.A(_02569_),
    .B(_02742_),
    .C(_02902_),
    .D(_03064_),
    .X(_03213_));
 sky130_fd_sc_hd__a21o_1 _10299_ (.A1(_02570_),
    .A2(_02572_),
    .B1(_03213_),
    .X(_03214_));
 sky130_fd_sc_hd__a21oi_2 _10300_ (.A1(_02900_),
    .A2(_03062_),
    .B1(_03063_),
    .Y(_03215_));
 sky130_fd_sc_hd__o21ba_1 _10301_ (.A1(_02905_),
    .A2(_03212_),
    .B1_N(_03215_),
    .X(_03216_));
 sky130_fd_sc_hd__nand2_1 _10302_ (.A(_03214_),
    .B(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__xnor2_2 _10303_ (.A(_03211_),
    .B(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__o21ai_1 _10304_ (.A1(_03116_),
    .A2(_03218_),
    .B1(_02348_),
    .Y(_03219_));
 sky130_fd_sc_hd__a21oi_1 _10305_ (.A1(_03116_),
    .A2(_03218_),
    .B1(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__nand3_1 _10306_ (.A(net136),
    .B(_01931_),
    .C(_01932_),
    .Y(_03221_));
 sky130_fd_sc_hd__a21o_1 _10307_ (.A1(net136),
    .A2(_01931_),
    .B1(_01932_),
    .X(_03222_));
 sky130_fd_sc_hd__a21o_1 _10308_ (.A1(_06557_),
    .A2(_03077_),
    .B1(_06549_),
    .X(_03223_));
 sky130_fd_sc_hd__a21oi_1 _10309_ (.A1(_06550_),
    .A2(_03223_),
    .B1(net295),
    .Y(_03224_));
 sky130_fd_sc_hd__a31o_1 _10310_ (.A1(net295),
    .A2(_06548_),
    .A3(_06582_),
    .B1(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__xor2_1 _10311_ (.A(_06544_),
    .B(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__o21ai_2 _10312_ (.A1(net219),
    .A2(_02769_),
    .B1(_02453_),
    .Y(_03227_));
 sky130_fd_sc_hd__inv_2 _10313_ (.A(_03227_),
    .Y(_03228_));
 sky130_fd_sc_hd__a21oi_2 _10314_ (.A1(net220),
    .A2(_03227_),
    .B1(_02455_),
    .Y(_03229_));
 sky130_fd_sc_hd__mux2_1 _10315_ (.A0(_02587_),
    .A1(_02594_),
    .S(net215),
    .X(_03230_));
 sky130_fd_sc_hd__mux2_1 _10316_ (.A0(_02591_),
    .A1(_02602_),
    .S(net215),
    .X(_03231_));
 sky130_fd_sc_hd__mux2_1 _10317_ (.A0(_03230_),
    .A1(_03231_),
    .S(net218),
    .X(_03232_));
 sky130_fd_sc_hd__mux2_1 _10318_ (.A0(_02599_),
    .A1(_02608_),
    .S(net215),
    .X(_03233_));
 sky130_fd_sc_hd__mux2_1 _10319_ (.A0(_02753_),
    .A1(_03233_),
    .S(_06553_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_2 _10320_ (.A0(_03232_),
    .A1(_03234_),
    .S(net221),
    .X(_03235_));
 sky130_fd_sc_hd__a21o_1 _10321_ (.A1(net223),
    .A2(net205),
    .B1(net167),
    .X(_03236_));
 sky130_fd_sc_hd__o21ai_1 _10322_ (.A1(\div_res[4] ),
    .A2(_03098_),
    .B1(net140),
    .Y(_03237_));
 sky130_fd_sc_hd__xnor2_1 _10323_ (.A(\div_res[5] ),
    .B(_03237_),
    .Y(_03238_));
 sky130_fd_sc_hd__a21oi_1 _10324_ (.A1(_06541_),
    .A2(net195),
    .B1(net193),
    .Y(_03239_));
 sky130_fd_sc_hd__or2_1 _10325_ (.A(\div_shifter[36] ),
    .B(_03102_),
    .X(_03240_));
 sky130_fd_sc_hd__a21oi_4 _10326_ (.A1(net230),
    .A2(_03240_),
    .B1(\div_shifter[37] ),
    .Y(_03241_));
 sky130_fd_sc_hd__a31o_1 _10327_ (.A1(\div_shifter[37] ),
    .A2(net230),
    .A3(_03240_),
    .B1(net192),
    .X(_03242_));
 sky130_fd_sc_hd__o2bb2a_1 _10328_ (.A1_N(_06687_),
    .A2_N(net256),
    .B1(net231),
    .B2(reg1_val[5]),
    .X(_03243_));
 sky130_fd_sc_hd__o221a_1 _10329_ (.A1(_06538_),
    .A2(net203),
    .B1(_03241_),
    .B2(_03242_),
    .C1(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__o221ai_2 _10330_ (.A1(_06541_),
    .A2(net194),
    .B1(_03239_),
    .B2(_06543_),
    .C1(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__o21a_1 _10331_ (.A1(_03082_),
    .A2(_03083_),
    .B1(_03084_),
    .X(_03246_));
 sky130_fd_sc_hd__nor2_1 _10332_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03247_));
 sky130_fd_sc_hd__nand2_1 _10333_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03248_));
 sky130_fd_sc_hd__and2b_1 _10334_ (.A_N(_03247_),
    .B(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__xnor2_1 _10335_ (.A(_03246_),
    .B(_03249_),
    .Y(_03250_));
 sky130_fd_sc_hd__a31o_1 _10336_ (.A1(net244),
    .A2(net205),
    .A3(_03250_),
    .B1(_03245_),
    .X(_03251_));
 sky130_fd_sc_hd__a221o_1 _10337_ (.A1(_03235_),
    .A2(_03236_),
    .B1(_03238_),
    .B2(_02443_),
    .C1(_03251_),
    .X(_03252_));
 sky130_fd_sc_hd__a221o_1 _10338_ (.A1(net234),
    .A2(_03226_),
    .B1(_03229_),
    .B2(net172),
    .C1(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__a311o_1 _10339_ (.A1(net233),
    .A2(_03221_),
    .A3(_03222_),
    .B1(_03253_),
    .C1(_03220_),
    .X(_03254_));
 sky130_fd_sc_hd__and3_1 _10340_ (.A(curr_PC[4]),
    .B(curr_PC[5]),
    .C(_02958_),
    .X(_03255_));
 sky130_fd_sc_hd__a21o_1 _10341_ (.A1(curr_PC[4]),
    .A2(_02958_),
    .B1(curr_PC[5]),
    .X(_03256_));
 sky130_fd_sc_hd__nand2_1 _10342_ (.A(net242),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__a2bb2o_4 _10343_ (.A1_N(_03255_),
    .A2_N(_03257_),
    .B1(net237),
    .B2(_03254_),
    .X(dest_val[5]));
 sky130_fd_sc_hd__or2_1 _10344_ (.A(_03115_),
    .B(_03218_),
    .X(_03258_));
 sky130_fd_sc_hd__a21oi_4 _10345_ (.A1(_03118_),
    .A2(_03207_),
    .B1(_03206_),
    .Y(_03259_));
 sky130_fd_sc_hd__a21bo_2 _10346_ (.A1(_03196_),
    .A2(_03202_),
    .B1_N(_03204_),
    .X(_03260_));
 sky130_fd_sc_hd__a21o_1 _10347_ (.A1(_03151_),
    .A2(_03155_),
    .B1(_03154_),
    .X(_03261_));
 sky130_fd_sc_hd__o211a_1 _10348_ (.A1(_03164_),
    .A2(_03166_),
    .B1(net107),
    .C1(net63),
    .X(_03262_));
 sky130_fd_sc_hd__a211o_1 _10349_ (.A1(net107),
    .A2(net63),
    .B1(_03164_),
    .C1(_03166_),
    .X(_03263_));
 sky130_fd_sc_hd__and2b_1 _10350_ (.A_N(_03262_),
    .B(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__xor2_1 _10351_ (.A(_03261_),
    .B(_03264_),
    .X(_03265_));
 sky130_fd_sc_hd__o22a_2 _10352_ (.A1(net49),
    .A2(net75),
    .B1(_00466_),
    .B2(net51),
    .X(_03266_));
 sky130_fd_sc_hd__xnor2_4 _10353_ (.A(net108),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__o32a_2 _10354_ (.A1(_00497_),
    .A2(_00513_),
    .A3(_00515_),
    .B1(net69),
    .B2(net44),
    .X(_03268_));
 sky130_fd_sc_hd__xnor2_4 _10355_ (.A(net145),
    .B(_03268_),
    .Y(_03269_));
 sky130_fd_sc_hd__o22a_1 _10356_ (.A1(net47),
    .A2(net83),
    .B1(net79),
    .B2(net45),
    .X(_03270_));
 sky130_fd_sc_hd__xnor2_2 _10357_ (.A(net117),
    .B(_03270_),
    .Y(_03271_));
 sky130_fd_sc_hd__and2_1 _10358_ (.A(_03269_),
    .B(_03271_),
    .X(_03272_));
 sky130_fd_sc_hd__xor2_4 _10359_ (.A(_03269_),
    .B(_03271_),
    .X(_03273_));
 sky130_fd_sc_hd__xnor2_4 _10360_ (.A(_03267_),
    .B(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__o21a_2 _10361_ (.A1(_03179_),
    .A2(_03185_),
    .B1(_03184_),
    .X(_03275_));
 sky130_fd_sc_hd__or2_1 _10362_ (.A(_03274_),
    .B(_03275_),
    .X(_03276_));
 sky130_fd_sc_hd__xnor2_4 _10363_ (.A(_03274_),
    .B(_03275_),
    .Y(_03277_));
 sky130_fd_sc_hd__a22o_1 _10364_ (.A1(net129),
    .A2(_00812_),
    .B1(net11),
    .B2(net127),
    .X(_03278_));
 sky130_fd_sc_hd__xor2_1 _10365_ (.A(net155),
    .B(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__or2_1 _10366_ (.A(_00193_),
    .B(net5),
    .X(_03280_));
 sky130_fd_sc_hd__a22o_1 _10367_ (.A1(_00195_),
    .A2(net6),
    .B1(_03280_),
    .B2(net175),
    .X(_03281_));
 sky130_fd_sc_hd__nor2_2 _10368_ (.A(_03279_),
    .B(_03281_),
    .Y(_03282_));
 sky130_fd_sc_hd__and2_1 _10369_ (.A(_03279_),
    .B(_03281_),
    .X(_03283_));
 sky130_fd_sc_hd__nor2_2 _10370_ (.A(_03282_),
    .B(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__xnor2_2 _10371_ (.A(_03277_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__a22o_1 _10372_ (.A1(_00375_),
    .A2(net17),
    .B1(net13),
    .B2(net122),
    .X(_03286_));
 sky130_fd_sc_hd__xnor2_2 _10373_ (.A(net65),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__a22o_1 _10374_ (.A1(net111),
    .A2(net9),
    .B1(net4),
    .B2(net112),
    .X(_03288_));
 sky130_fd_sc_hd__xnor2_2 _10375_ (.A(net60),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__o22a_1 _10376_ (.A1(net34),
    .A2(net115),
    .B1(_00398_),
    .B2(net32),
    .X(_03290_));
 sky130_fd_sc_hd__xnor2_2 _10377_ (.A(net94),
    .B(_03290_),
    .Y(_03291_));
 sky130_fd_sc_hd__and2_1 _10378_ (.A(_03289_),
    .B(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__xor2_2 _10379_ (.A(_03289_),
    .B(_03291_),
    .X(_03293_));
 sky130_fd_sc_hd__xnor2_2 _10380_ (.A(_03287_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__nor2_1 _10381_ (.A(_03285_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__xor2_2 _10382_ (.A(_03285_),
    .B(_03294_),
    .X(_03296_));
 sky130_fd_sc_hd__xor2_1 _10383_ (.A(_03265_),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__a21o_1 _10384_ (.A1(_03121_),
    .A2(_03129_),
    .B1(_03126_),
    .X(_03298_));
 sky130_fd_sc_hd__o22a_1 _10385_ (.A1(net56),
    .A2(net25),
    .B1(net23),
    .B2(net53),
    .X(_03299_));
 sky130_fd_sc_hd__xnor2_1 _10386_ (.A(net87),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__o22a_1 _10387_ (.A1(_00202_),
    .A2(net29),
    .B1(net27),
    .B2(net40),
    .X(_03301_));
 sky130_fd_sc_hd__xnor2_1 _10388_ (.A(net89),
    .B(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__nand2_1 _10389_ (.A(_03300_),
    .B(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__or2_1 _10390_ (.A(_03300_),
    .B(_03302_),
    .X(_03304_));
 sky130_fd_sc_hd__nand2_1 _10391_ (.A(_03303_),
    .B(_03304_),
    .Y(_03305_));
 sky130_fd_sc_hd__nand2_1 _10392_ (.A(_03143_),
    .B(_03147_),
    .Y(_03306_));
 sky130_fd_sc_hd__xor2_1 _10393_ (.A(_03305_),
    .B(_03306_),
    .X(_03307_));
 sky130_fd_sc_hd__and2b_1 _10394_ (.A_N(_03307_),
    .B(_03298_),
    .X(_03308_));
 sky130_fd_sc_hd__xnor2_1 _10395_ (.A(_03298_),
    .B(_03307_),
    .Y(_03309_));
 sky130_fd_sc_hd__and2_1 _10396_ (.A(_03297_),
    .B(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__nor2_1 _10397_ (.A(_03297_),
    .B(_03309_),
    .Y(_03311_));
 sky130_fd_sc_hd__nor2_2 _10398_ (.A(_03310_),
    .B(_03311_),
    .Y(_03312_));
 sky130_fd_sc_hd__o21ai_4 _10399_ (.A1(_03036_),
    .A2(_03167_),
    .B1(_03169_),
    .Y(_03313_));
 sky130_fd_sc_hd__o22a_2 _10400_ (.A1(net38),
    .A2(_00463_),
    .B1(net70),
    .B2(net36),
    .X(_03314_));
 sky130_fd_sc_hd__xnor2_4 _10401_ (.A(net98),
    .B(_03314_),
    .Y(_03315_));
 sky130_fd_sc_hd__o22a_2 _10402_ (.A1(_00219_),
    .A2(net20),
    .B1(net18),
    .B2(net100),
    .X(_03316_));
 sky130_fd_sc_hd__xnor2_4 _10403_ (.A(net97),
    .B(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__a22o_1 _10404_ (.A1(net14),
    .A2(_00443_),
    .B1(_00446_),
    .B2(net30),
    .X(_03318_));
 sky130_fd_sc_hd__xnor2_4 _10405_ (.A(net91),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__nand2_1 _10406_ (.A(_03317_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__xnor2_4 _10407_ (.A(_03317_),
    .B(_03319_),
    .Y(_03321_));
 sky130_fd_sc_hd__inv_2 _10408_ (.A(_03321_),
    .Y(_03322_));
 sky130_fd_sc_hd__nand2_1 _10409_ (.A(_03315_),
    .B(_03322_),
    .Y(_03323_));
 sky130_fd_sc_hd__xor2_4 _10410_ (.A(_03315_),
    .B(_03321_),
    .X(_03324_));
 sky130_fd_sc_hd__a21oi_4 _10411_ (.A1(_03135_),
    .A2(_03137_),
    .B1(_03136_),
    .Y(_03325_));
 sky130_fd_sc_hd__xnor2_4 _10412_ (.A(_03324_),
    .B(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__and2b_1 _10413_ (.A_N(_03326_),
    .B(_03313_),
    .X(_03327_));
 sky130_fd_sc_hd__xnor2_4 _10414_ (.A(_03313_),
    .B(_03326_),
    .Y(_03328_));
 sky130_fd_sc_hd__xor2_4 _10415_ (.A(_03312_),
    .B(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__a21o_1 _10416_ (.A1(_03134_),
    .A2(_03193_),
    .B1(_03191_),
    .X(_03330_));
 sky130_fd_sc_hd__a21o_1 _10417_ (.A1(_03119_),
    .A2(_03133_),
    .B1(_03131_),
    .X(_03331_));
 sky130_fd_sc_hd__a21oi_2 _10418_ (.A1(_03139_),
    .A2(_03172_),
    .B1(_03171_),
    .Y(_03332_));
 sky130_fd_sc_hd__o21ai_2 _10419_ (.A1(_03176_),
    .A2(_03189_),
    .B1(_03188_),
    .Y(_03333_));
 sky130_fd_sc_hd__and2b_1 _10420_ (.A_N(_03332_),
    .B(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__xnor2_2 _10421_ (.A(_03332_),
    .B(_03333_),
    .Y(_03335_));
 sky130_fd_sc_hd__xnor2_2 _10422_ (.A(_03331_),
    .B(_03335_),
    .Y(_03336_));
 sky130_fd_sc_hd__a21boi_4 _10423_ (.A1(_03197_),
    .A2(_03201_),
    .B1_N(_03200_),
    .Y(_03337_));
 sky130_fd_sc_hd__xnor2_2 _10424_ (.A(_03336_),
    .B(_03337_),
    .Y(_03338_));
 sky130_fd_sc_hd__and2b_1 _10425_ (.A_N(_03338_),
    .B(_03330_),
    .X(_03339_));
 sky130_fd_sc_hd__xnor2_2 _10426_ (.A(_03330_),
    .B(_03338_),
    .Y(_03340_));
 sky130_fd_sc_hd__and2_1 _10427_ (.A(_03329_),
    .B(_03340_),
    .X(_03341_));
 sky130_fd_sc_hd__xor2_4 _10428_ (.A(_03329_),
    .B(_03340_),
    .X(_03342_));
 sky130_fd_sc_hd__xnor2_4 _10429_ (.A(_03260_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__or2_1 _10430_ (.A(_03259_),
    .B(_03343_),
    .X(_03344_));
 sky130_fd_sc_hd__and2_1 _10431_ (.A(_03259_),
    .B(_03343_),
    .X(_03345_));
 sky130_fd_sc_hd__xnor2_4 _10432_ (.A(_03259_),
    .B(_03343_),
    .Y(_03346_));
 sky130_fd_sc_hd__or4_2 _10433_ (.A(_02742_),
    .B(_02902_),
    .C(_03064_),
    .D(_03211_),
    .X(_03347_));
 sky130_fd_sc_hd__a21o_1 _10434_ (.A1(_02745_),
    .A2(_02746_),
    .B1(_03347_),
    .X(_03348_));
 sky130_fd_sc_hd__or3_1 _10435_ (.A(_02127_),
    .B(_02743_),
    .C(_03347_),
    .X(_03349_));
 sky130_fd_sc_hd__a21oi_2 _10436_ (.A1(_03062_),
    .A2(_03209_),
    .B1(_03210_),
    .Y(_03350_));
 sky130_fd_sc_hd__a2111oi_1 _10437_ (.A1(_02741_),
    .A2(_02900_),
    .B1(_02901_),
    .C1(_03064_),
    .D1(_03211_),
    .Y(_03351_));
 sky130_fd_sc_hd__nor2_1 _10438_ (.A(_03350_),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__a31o_1 _10439_ (.A1(_03348_),
    .A2(_03349_),
    .A3(_03352_),
    .B1(_03346_),
    .X(_03353_));
 sky130_fd_sc_hd__o211ai_2 _10440_ (.A1(_02747_),
    .A2(_03347_),
    .B1(_03352_),
    .C1(_03346_),
    .Y(_03354_));
 sky130_fd_sc_hd__and2_1 _10441_ (.A(_03353_),
    .B(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__a21o_1 _10442_ (.A1(net137),
    .A2(_03258_),
    .B1(_03355_),
    .X(_03356_));
 sky130_fd_sc_hd__a31oi_1 _10443_ (.A1(net137),
    .A2(_03258_),
    .A3(_03355_),
    .B1(net235),
    .Y(_03357_));
 sky130_fd_sc_hd__o21a_1 _10444_ (.A1(_01931_),
    .A2(_01932_),
    .B1(net136),
    .X(_03358_));
 sky130_fd_sc_hd__xnor2_1 _10445_ (.A(_01933_),
    .B(_03358_),
    .Y(_03359_));
 sky130_fd_sc_hd__a31oi_1 _10446_ (.A1(_06541_),
    .A2(_06550_),
    .A3(_03223_),
    .B1(_06543_),
    .Y(_03360_));
 sky130_fd_sc_hd__and3_1 _10447_ (.A(net295),
    .B(_06540_),
    .C(_06583_),
    .X(_03361_));
 sky130_fd_sc_hd__a21o_1 _10448_ (.A1(net283),
    .A2(_03360_),
    .B1(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__xor2_1 _10449_ (.A(_06535_),
    .B(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__o21ai_2 _10450_ (.A1(net219),
    .A2(_02609_),
    .B1(_02453_),
    .Y(_03364_));
 sky130_fd_sc_hd__inv_2 _10451_ (.A(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__a21oi_2 _10452_ (.A1(net220),
    .A2(_03364_),
    .B1(_02455_),
    .Y(_03366_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(_02759_),
    .A1(_02762_),
    .S(net215),
    .X(_03367_));
 sky130_fd_sc_hd__mux2_1 _10454_ (.A0(_02761_),
    .A1(_02766_),
    .S(net215),
    .X(_03368_));
 sky130_fd_sc_hd__mux2_1 _10455_ (.A0(_03367_),
    .A1(_03368_),
    .S(net218),
    .X(_03369_));
 sky130_fd_sc_hd__mux2_1 _10456_ (.A0(_02765_),
    .A1(_02768_),
    .S(net216),
    .X(_03370_));
 sky130_fd_sc_hd__mux2_1 _10457_ (.A0(_02632_),
    .A1(_03370_),
    .S(_06553_),
    .X(_03371_));
 sky130_fd_sc_hd__mux2_1 _10458_ (.A0(_03369_),
    .A1(_03371_),
    .S(net221),
    .X(_03372_));
 sky130_fd_sc_hd__or3_1 _10459_ (.A(\div_res[5] ),
    .B(\div_res[4] ),
    .C(_03098_),
    .X(_03373_));
 sky130_fd_sc_hd__a21oi_1 _10460_ (.A1(net140),
    .A2(_03373_),
    .B1(\div_res[6] ),
    .Y(_03374_));
 sky130_fd_sc_hd__a31o_1 _10461_ (.A1(\div_res[6] ),
    .A2(net140),
    .A3(_03373_),
    .B1(net189),
    .X(_03375_));
 sky130_fd_sc_hd__a21oi_1 _10462_ (.A1(_06534_),
    .A2(net195),
    .B1(net193),
    .Y(_03376_));
 sky130_fd_sc_hd__or3_2 _10463_ (.A(\div_shifter[37] ),
    .B(\div_shifter[36] ),
    .C(_03102_),
    .X(_03377_));
 sky130_fd_sc_hd__a21oi_4 _10464_ (.A1(net230),
    .A2(_03377_),
    .B1(\div_shifter[38] ),
    .Y(_03378_));
 sky130_fd_sc_hd__a31o_2 _10465_ (.A1(\div_shifter[38] ),
    .A2(net230),
    .A3(_03377_),
    .B1(net192),
    .X(_03379_));
 sky130_fd_sc_hd__o2bb2a_1 _10466_ (.A1_N(_00190_),
    .A2_N(net256),
    .B1(net231),
    .B2(reg1_val[6]),
    .X(_03380_));
 sky130_fd_sc_hd__o221a_1 _10467_ (.A1(_06530_),
    .A2(net203),
    .B1(_03378_),
    .B2(_03379_),
    .C1(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__o221a_1 _10468_ (.A1(_06534_),
    .A2(net194),
    .B1(_03376_),
    .B2(_06532_),
    .C1(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__o21a_1 _10469_ (.A1(_03246_),
    .A2(_03247_),
    .B1(_03248_),
    .X(_03383_));
 sky130_fd_sc_hd__nor2_1 _10470_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03384_));
 sky130_fd_sc_hd__nand2_1 _10471_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03385_));
 sky130_fd_sc_hd__nand2b_1 _10472_ (.A_N(_03384_),
    .B(_03385_),
    .Y(_03386_));
 sky130_fd_sc_hd__xnor2_1 _10473_ (.A(_03383_),
    .B(_03386_),
    .Y(_03387_));
 sky130_fd_sc_hd__o31a_1 _10474_ (.A1(net223),
    .A2(_06667_),
    .A3(_03387_),
    .B1(_03382_),
    .X(_03388_));
 sky130_fd_sc_hd__o21ai_1 _10475_ (.A1(_03374_),
    .A2(_03375_),
    .B1(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__a221o_1 _10476_ (.A1(net172),
    .A2(_03366_),
    .B1(_03372_),
    .B2(_03236_),
    .C1(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__a21o_1 _10477_ (.A1(net234),
    .A2(_03363_),
    .B1(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__a221o_1 _10478_ (.A1(_03356_),
    .A2(_03357_),
    .B1(_03359_),
    .B2(net233),
    .C1(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__or2_1 _10479_ (.A(curr_PC[6]),
    .B(_03255_),
    .X(_03393_));
 sky130_fd_sc_hd__and2_1 _10480_ (.A(curr_PC[6]),
    .B(_03255_),
    .X(_03394_));
 sky130_fd_sc_hd__nor2_1 _10481_ (.A(net237),
    .B(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__a22o_4 _10482_ (.A1(net237),
    .A2(_03392_),
    .B1(_03393_),
    .B2(_03395_),
    .X(dest_val[6]));
 sky130_fd_sc_hd__o21a_1 _10483_ (.A1(_03258_),
    .A2(_03355_),
    .B1(net137),
    .X(_03396_));
 sky130_fd_sc_hd__a21oi_4 _10484_ (.A1(_03260_),
    .A2(_03342_),
    .B1(_03341_),
    .Y(_03397_));
 sky130_fd_sc_hd__o21bai_4 _10485_ (.A1(_03336_),
    .A2(_03337_),
    .B1_N(_03339_),
    .Y(_03398_));
 sky130_fd_sc_hd__o21ai_4 _10486_ (.A1(_03277_),
    .A2(_03284_),
    .B1(_03276_),
    .Y(_03399_));
 sky130_fd_sc_hd__a21o_2 _10487_ (.A1(_03261_),
    .A2(_03263_),
    .B1(_03262_),
    .X(_03400_));
 sky130_fd_sc_hd__o22a_2 _10488_ (.A1(_00230_),
    .A2(net20),
    .B1(net18),
    .B2(net42),
    .X(_03401_));
 sky130_fd_sc_hd__xnor2_4 _10489_ (.A(_00274_),
    .B(_03401_),
    .Y(_03402_));
 sky130_fd_sc_hd__o22a_1 _10490_ (.A1(_00219_),
    .A2(net36),
    .B1(net70),
    .B2(net38),
    .X(_03403_));
 sky130_fd_sc_hd__xnor2_1 _10491_ (.A(_00262_),
    .B(_03403_),
    .Y(_03404_));
 sky130_fd_sc_hd__o22a_1 _10492_ (.A1(net41),
    .A2(net29),
    .B1(net27),
    .B2(net57),
    .X(_03405_));
 sky130_fd_sc_hd__xnor2_1 _10493_ (.A(net89),
    .B(_03405_),
    .Y(_03406_));
 sky130_fd_sc_hd__nand2_1 _10494_ (.A(_03404_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__or2_1 _10495_ (.A(_03404_),
    .B(_03406_),
    .X(_03408_));
 sky130_fd_sc_hd__nand2_2 _10496_ (.A(_03407_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__xor2_4 _10497_ (.A(_03402_),
    .B(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__nand2_1 _10498_ (.A(_03400_),
    .B(_03410_),
    .Y(_03411_));
 sky130_fd_sc_hd__xor2_4 _10499_ (.A(_03400_),
    .B(_03410_),
    .X(_03412_));
 sky130_fd_sc_hd__xnor2_4 _10500_ (.A(_03399_),
    .B(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__o22a_1 _10501_ (.A1(net46),
    .A2(net84),
    .B1(net80),
    .B2(net49),
    .X(_03414_));
 sky130_fd_sc_hd__xnor2_1 _10502_ (.A(net117),
    .B(_03414_),
    .Y(_03415_));
 sky130_fd_sc_hd__inv_2 _10503_ (.A(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__o22a_1 _10504_ (.A1(net54),
    .A2(net25),
    .B1(net23),
    .B2(net48),
    .X(_03417_));
 sky130_fd_sc_hd__xnor2_1 _10505_ (.A(net87),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__o22a_1 _10506_ (.A1(net51),
    .A2(_00460_),
    .B1(_00466_),
    .B2(net43),
    .X(_03419_));
 sky130_fd_sc_hd__xnor2_1 _10507_ (.A(net108),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__xnor2_1 _10508_ (.A(_03418_),
    .B(_03420_),
    .Y(_03421_));
 sky130_fd_sc_hd__or2_1 _10509_ (.A(_03416_),
    .B(_03421_),
    .X(_03422_));
 sky130_fd_sc_hd__nand2_1 _10510_ (.A(_03416_),
    .B(_03421_),
    .Y(_03423_));
 sky130_fd_sc_hd__nand2_1 _10511_ (.A(_03422_),
    .B(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__a21o_1 _10512_ (.A1(_03287_),
    .A2(_03293_),
    .B1(_03292_),
    .X(_03425_));
 sky130_fd_sc_hd__xor2_1 _10513_ (.A(_03424_),
    .B(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__a21oi_1 _10514_ (.A1(_03320_),
    .A2(_03323_),
    .B1(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__and3_1 _10515_ (.A(_03320_),
    .B(_03323_),
    .C(_03426_),
    .X(_03428_));
 sky130_fd_sc_hd__nor2_1 _10516_ (.A(_03427_),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__a22o_1 _10517_ (.A1(net122),
    .A2(net9),
    .B1(net4),
    .B2(net111),
    .X(_03430_));
 sky130_fd_sc_hd__xnor2_1 _10518_ (.A(net63),
    .B(_03430_),
    .Y(_03431_));
 sky130_fd_sc_hd__nor2_1 _10519_ (.A(_03282_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__and2_1 _10520_ (.A(_03282_),
    .B(_03431_),
    .X(_03433_));
 sky130_fd_sc_hd__nor2_1 _10521_ (.A(_03432_),
    .B(_03433_),
    .Y(_03434_));
 sky130_fd_sc_hd__nor2_1 _10522_ (.A(net113),
    .B(net60),
    .Y(_03435_));
 sky130_fd_sc_hd__xnor2_1 _10523_ (.A(_03434_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__o22a_1 _10524_ (.A1(net34),
    .A2(_00398_),
    .B1(_00442_),
    .B2(net32),
    .X(_03437_));
 sky130_fd_sc_hd__xnor2_1 _10525_ (.A(_00302_),
    .B(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__o22a_1 _10526_ (.A1(_00336_),
    .A2(net77),
    .B1(_00463_),
    .B2(_00342_),
    .X(_03439_));
 sky130_fd_sc_hd__xnor2_1 _10527_ (.A(net92),
    .B(_03439_),
    .Y(_03440_));
 sky130_fd_sc_hd__o2bb2a_1 _10528_ (.A1_N(_00392_),
    .A2_N(net16),
    .B1(_00797_),
    .B2(net120),
    .X(_03441_));
 sky130_fd_sc_hd__xnor2_1 _10529_ (.A(_00787_),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__nand2_1 _10530_ (.A(_03440_),
    .B(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__xnor2_1 _10531_ (.A(_03440_),
    .B(_03442_),
    .Y(_03444_));
 sky130_fd_sc_hd__or2_1 _10532_ (.A(_03438_),
    .B(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__nand2_1 _10533_ (.A(_03438_),
    .B(_03444_),
    .Y(_03446_));
 sky130_fd_sc_hd__and2_1 _10534_ (.A(_03445_),
    .B(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__a21o_1 _10535_ (.A1(_03267_),
    .A2(_03273_),
    .B1(_03272_),
    .X(_03448_));
 sky130_fd_sc_hd__a22o_1 _10536_ (.A1(net129),
    .A2(net11),
    .B1(net6),
    .B2(net127),
    .X(_03449_));
 sky130_fd_sc_hd__xor2_2 _10537_ (.A(net155),
    .B(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__or3_1 _10538_ (.A(net69),
    .B(_00513_),
    .C(_00515_),
    .X(_03451_));
 sky130_fd_sc_hd__a21o_1 _10539_ (.A1(_00809_),
    .A2(_00810_),
    .B1(_00497_),
    .X(_03452_));
 sky130_fd_sc_hd__a21bo_1 _10540_ (.A1(_03451_),
    .A2(_03452_),
    .B1_N(net146),
    .X(_03453_));
 sky130_fd_sc_hd__nand3b_1 _10541_ (.A_N(net146),
    .B(_03451_),
    .C(_03452_),
    .Y(_03454_));
 sky130_fd_sc_hd__nand3_2 _10542_ (.A(_00188_),
    .B(_03453_),
    .C(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__a21o_1 _10543_ (.A1(_03453_),
    .A2(_03454_),
    .B1(_00188_),
    .X(_03456_));
 sky130_fd_sc_hd__nand3_2 _10544_ (.A(_03450_),
    .B(_03455_),
    .C(_03456_),
    .Y(_03457_));
 sky130_fd_sc_hd__a21o_1 _10545_ (.A1(_03455_),
    .A2(_03456_),
    .B1(_03450_),
    .X(_03458_));
 sky130_fd_sc_hd__nand3_2 _10546_ (.A(_03448_),
    .B(_03457_),
    .C(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__a21o_1 _10547_ (.A1(_03457_),
    .A2(_03458_),
    .B1(_03448_),
    .X(_03460_));
 sky130_fd_sc_hd__nand3b_1 _10548_ (.A_N(_03303_),
    .B(_03459_),
    .C(_03460_),
    .Y(_03461_));
 sky130_fd_sc_hd__a21bo_1 _10549_ (.A1(_03459_),
    .A2(_03460_),
    .B1_N(_03303_),
    .X(_03462_));
 sky130_fd_sc_hd__and3_1 _10550_ (.A(_03447_),
    .B(_03461_),
    .C(_03462_),
    .X(_03463_));
 sky130_fd_sc_hd__a21oi_1 _10551_ (.A1(_03461_),
    .A2(_03462_),
    .B1(_03447_),
    .Y(_03464_));
 sky130_fd_sc_hd__or3_1 _10552_ (.A(_03436_),
    .B(_03463_),
    .C(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__o21ai_1 _10553_ (.A1(_03463_),
    .A2(_03464_),
    .B1(_03436_),
    .Y(_03466_));
 sky130_fd_sc_hd__and3_1 _10554_ (.A(_03429_),
    .B(_03465_),
    .C(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__a21oi_1 _10555_ (.A1(_03465_),
    .A2(_03466_),
    .B1(_03429_),
    .Y(_03468_));
 sky130_fd_sc_hd__nor2_2 _10556_ (.A(_03467_),
    .B(_03468_),
    .Y(_03469_));
 sky130_fd_sc_hd__xnor2_4 _10557_ (.A(_03413_),
    .B(_03469_),
    .Y(_03470_));
 sky130_fd_sc_hd__a21o_1 _10558_ (.A1(_03312_),
    .A2(_03328_),
    .B1(_03310_),
    .X(_03471_));
 sky130_fd_sc_hd__a21oi_1 _10559_ (.A1(_03331_),
    .A2(_03335_),
    .B1(_03334_),
    .Y(_03472_));
 sky130_fd_sc_hd__o21bai_1 _10560_ (.A1(_03324_),
    .A2(_03325_),
    .B1_N(_03327_),
    .Y(_03473_));
 sky130_fd_sc_hd__a21oi_2 _10561_ (.A1(_03265_),
    .A2(_03296_),
    .B1(_03295_),
    .Y(_03474_));
 sky130_fd_sc_hd__a31oi_2 _10562_ (.A1(_03303_),
    .A2(_03304_),
    .A3(_03306_),
    .B1(_03308_),
    .Y(_03475_));
 sky130_fd_sc_hd__nor2_1 _10563_ (.A(_03474_),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__xor2_1 _10564_ (.A(_03474_),
    .B(_03475_),
    .X(_03477_));
 sky130_fd_sc_hd__xnor2_1 _10565_ (.A(_03473_),
    .B(_03477_),
    .Y(_03478_));
 sky130_fd_sc_hd__or2_1 _10566_ (.A(_03472_),
    .B(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__xnor2_1 _10567_ (.A(_03472_),
    .B(_03478_),
    .Y(_03480_));
 sky130_fd_sc_hd__nand2b_1 _10568_ (.A_N(_03480_),
    .B(_03471_),
    .Y(_03481_));
 sky130_fd_sc_hd__xnor2_2 _10569_ (.A(_03471_),
    .B(_03480_),
    .Y(_03482_));
 sky130_fd_sc_hd__and2_1 _10570_ (.A(_03470_),
    .B(_03482_),
    .X(_03483_));
 sky130_fd_sc_hd__xor2_4 _10571_ (.A(_03470_),
    .B(_03482_),
    .X(_03484_));
 sky130_fd_sc_hd__xnor2_4 _10572_ (.A(_03398_),
    .B(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__or2_1 _10573_ (.A(_03397_),
    .B(_03485_),
    .X(_03486_));
 sky130_fd_sc_hd__and2_1 _10574_ (.A(_03397_),
    .B(_03485_),
    .X(_03487_));
 sky130_fd_sc_hd__xnor2_4 _10575_ (.A(_03397_),
    .B(_03485_),
    .Y(_03488_));
 sky130_fd_sc_hd__nor2_1 _10576_ (.A(_03211_),
    .B(_03346_),
    .Y(_03489_));
 sky130_fd_sc_hd__or4_1 _10577_ (.A(_02902_),
    .B(_03064_),
    .C(_03211_),
    .D(_03346_),
    .X(_03490_));
 sky130_fd_sc_hd__a21o_1 _10578_ (.A1(_02905_),
    .A2(_02906_),
    .B1(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__or3_1 _10579_ (.A(_02239_),
    .B(_02903_),
    .C(_03490_),
    .X(_03492_));
 sky130_fd_sc_hd__a21oi_2 _10580_ (.A1(_03209_),
    .A2(_03344_),
    .B1(_03345_),
    .Y(_03493_));
 sky130_fd_sc_hd__a21oi_1 _10581_ (.A1(_03215_),
    .A2(_03489_),
    .B1(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__o21ai_1 _10582_ (.A1(_02907_),
    .A2(_03490_),
    .B1(_03494_),
    .Y(_03495_));
 sky130_fd_sc_hd__xnor2_2 _10583_ (.A(_03488_),
    .B(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__o21ai_1 _10584_ (.A1(_03396_),
    .A2(_03496_),
    .B1(_02348_),
    .Y(_03497_));
 sky130_fd_sc_hd__a21oi_1 _10585_ (.A1(_03396_),
    .A2(_03496_),
    .B1(_03497_),
    .Y(_03498_));
 sky130_fd_sc_hd__o21ai_1 _10586_ (.A1(net134),
    .A2(_01934_),
    .B1(_01937_),
    .Y(_03499_));
 sky130_fd_sc_hd__o31a_1 _10587_ (.A1(net134),
    .A2(_01934_),
    .A3(_01937_),
    .B1(net233),
    .X(_03500_));
 sky130_fd_sc_hd__and3_1 _10588_ (.A(net295),
    .B(_06531_),
    .C(_06584_),
    .X(_03501_));
 sky130_fd_sc_hd__nor2_1 _10589_ (.A(_06533_),
    .B(_03360_),
    .Y(_03502_));
 sky130_fd_sc_hd__nor2_1 _10590_ (.A(_06532_),
    .B(_03502_),
    .Y(_03503_));
 sky130_fd_sc_hd__a21o_1 _10591_ (.A1(net283),
    .A2(_03503_),
    .B1(_03501_),
    .X(_03504_));
 sky130_fd_sc_hd__nand2_1 _10592_ (.A(_06527_),
    .B(_03504_),
    .Y(_03505_));
 sky130_fd_sc_hd__o211a_1 _10593_ (.A1(_06527_),
    .A2(_03504_),
    .B1(_03505_),
    .C1(net234),
    .X(_03506_));
 sky130_fd_sc_hd__o21ai_2 _10594_ (.A1(net219),
    .A2(_02416_),
    .B1(_02453_),
    .Y(_03507_));
 sky130_fd_sc_hd__inv_2 _10595_ (.A(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__a21oi_2 _10596_ (.A1(net220),
    .A2(_03507_),
    .B1(_02455_),
    .Y(_03509_));
 sky130_fd_sc_hd__mux2_1 _10597_ (.A0(_02915_),
    .A1(_02918_),
    .S(net215),
    .X(_03510_));
 sky130_fd_sc_hd__mux2_1 _10598_ (.A0(_02917_),
    .A1(_02922_),
    .S(net215),
    .X(_03511_));
 sky130_fd_sc_hd__mux2_1 _10599_ (.A0(_03510_),
    .A1(_03511_),
    .S(net218),
    .X(_03512_));
 sky130_fd_sc_hd__mux2_1 _10600_ (.A0(_02921_),
    .A1(_02924_),
    .S(net215),
    .X(_03513_));
 sky130_fd_sc_hd__and3_1 _10601_ (.A(net218),
    .B(_02451_),
    .C(_02452_),
    .X(_03514_));
 sky130_fd_sc_hd__a21o_1 _10602_ (.A1(_06553_),
    .A2(_03513_),
    .B1(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__mux2_1 _10603_ (.A0(_03512_),
    .A1(_03515_),
    .S(net222),
    .X(_03516_));
 sky130_fd_sc_hd__or2_1 _10604_ (.A(\div_res[6] ),
    .B(_03373_),
    .X(_03517_));
 sky130_fd_sc_hd__a21oi_1 _10605_ (.A1(net140),
    .A2(_03517_),
    .B1(\div_res[7] ),
    .Y(_03518_));
 sky130_fd_sc_hd__a31o_1 _10606_ (.A1(\div_res[7] ),
    .A2(net140),
    .A3(_03517_),
    .B1(net189),
    .X(_03519_));
 sky130_fd_sc_hd__a21oi_1 _10607_ (.A1(_06526_),
    .A2(net195),
    .B1(net193),
    .Y(_03520_));
 sky130_fd_sc_hd__nor2_1 _10608_ (.A(reg1_val[7]),
    .B(net232),
    .Y(_03521_));
 sky130_fd_sc_hd__a221o_2 _10609_ (.A1(_06523_),
    .A2(_06677_),
    .B1(_00186_),
    .B2(net257),
    .C1(_03521_),
    .X(_03522_));
 sky130_fd_sc_hd__or2_1 _10610_ (.A(\div_shifter[38] ),
    .B(_03377_),
    .X(_03523_));
 sky130_fd_sc_hd__a21oi_1 _10611_ (.A1(net229),
    .A2(_03523_),
    .B1(\div_shifter[39] ),
    .Y(_03524_));
 sky130_fd_sc_hd__a31o_1 _10612_ (.A1(\div_shifter[39] ),
    .A2(net229),
    .A3(_03523_),
    .B1(net191),
    .X(_03525_));
 sky130_fd_sc_hd__o21ba_1 _10613_ (.A1(_03524_),
    .A2(_03525_),
    .B1_N(_03522_),
    .X(_03526_));
 sky130_fd_sc_hd__o221a_1 _10614_ (.A1(_06526_),
    .A2(net194),
    .B1(_03520_),
    .B2(_06525_),
    .C1(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__o21ai_1 _10615_ (.A1(_03518_),
    .A2(_03519_),
    .B1(_03527_),
    .Y(_03528_));
 sky130_fd_sc_hd__o21a_1 _10616_ (.A1(_03383_),
    .A2(_03384_),
    .B1(_03385_),
    .X(_03529_));
 sky130_fd_sc_hd__nor2_1 _10617_ (.A(net287),
    .B(curr_PC[7]),
    .Y(_03530_));
 sky130_fd_sc_hd__nand2_1 _10618_ (.A(net287),
    .B(curr_PC[7]),
    .Y(_03531_));
 sky130_fd_sc_hd__and2b_1 _10619_ (.A_N(_03530_),
    .B(_03531_),
    .X(_03532_));
 sky130_fd_sc_hd__xnor2_1 _10620_ (.A(_03529_),
    .B(_03532_),
    .Y(_03533_));
 sky130_fd_sc_hd__a31o_1 _10621_ (.A1(net244),
    .A2(net205),
    .A3(_03533_),
    .B1(_03528_),
    .X(_03534_));
 sky130_fd_sc_hd__a221o_1 _10622_ (.A1(net172),
    .A2(_03509_),
    .B1(_03516_),
    .B2(_03236_),
    .C1(_03534_),
    .X(_03535_));
 sky130_fd_sc_hd__a211o_1 _10623_ (.A1(_03499_),
    .A2(_03500_),
    .B1(_03506_),
    .C1(_03535_),
    .X(_03536_));
 sky130_fd_sc_hd__o21a_1 _10624_ (.A1(_03498_),
    .A2(_03536_),
    .B1(net238),
    .X(_03537_));
 sky130_fd_sc_hd__nand2_1 _10625_ (.A(curr_PC[7]),
    .B(_03394_),
    .Y(_03538_));
 sky130_fd_sc_hd__or2_1 _10626_ (.A(curr_PC[7]),
    .B(_03394_),
    .X(_03539_));
 sky130_fd_sc_hd__a31o_4 _10627_ (.A1(net242),
    .A2(_03538_),
    .A3(_03539_),
    .B1(_03537_),
    .X(dest_val[7]));
 sky130_fd_sc_hd__a21oi_2 _10628_ (.A1(_03344_),
    .A2(_03486_),
    .B1(_03487_),
    .Y(_03540_));
 sky130_fd_sc_hd__nor2_1 _10629_ (.A(_03346_),
    .B(_03488_),
    .Y(_03541_));
 sky130_fd_sc_hd__a21oi_1 _10630_ (.A1(_03350_),
    .A2(_03541_),
    .B1(_03540_),
    .Y(_03542_));
 sky130_fd_sc_hd__or4_2 _10631_ (.A(_03064_),
    .B(_03211_),
    .C(_03346_),
    .D(_03488_),
    .X(_03543_));
 sky130_fd_sc_hd__a211o_1 _10632_ (.A1(_02242_),
    .A2(_02244_),
    .B1(_03066_),
    .C1(_03543_),
    .X(_03544_));
 sky130_fd_sc_hd__o211a_4 _10633_ (.A1(_03069_),
    .A2(_03543_),
    .B1(_03544_),
    .C1(_03542_),
    .X(_03545_));
 sky130_fd_sc_hd__a21o_2 _10634_ (.A1(_03398_),
    .A2(_03484_),
    .B1(_03483_),
    .X(_03546_));
 sky130_fd_sc_hd__a22o_1 _10635_ (.A1(_00375_),
    .A2(net8),
    .B1(net3),
    .B2(net122),
    .X(_03547_));
 sky130_fd_sc_hd__xnor2_1 _10636_ (.A(net59),
    .B(_03547_),
    .Y(_03548_));
 sky130_fd_sc_hd__nand2_1 _10637_ (.A(net111),
    .B(net61),
    .Y(_03549_));
 sky130_fd_sc_hd__a22o_1 _10638_ (.A1(_00397_),
    .A2(net16),
    .B1(net12),
    .B2(_00392_),
    .X(_03550_));
 sky130_fd_sc_hd__xnor2_1 _10639_ (.A(net64),
    .B(_03550_),
    .Y(_03551_));
 sky130_fd_sc_hd__nand2b_1 _10640_ (.A_N(_03549_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__xnor2_1 _10641_ (.A(_03549_),
    .B(_03551_),
    .Y(_03553_));
 sky130_fd_sc_hd__nand2_1 _10642_ (.A(_03548_),
    .B(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__or2_1 _10643_ (.A(_03548_),
    .B(_03553_),
    .X(_03555_));
 sky130_fd_sc_hd__nand2_1 _10644_ (.A(_03554_),
    .B(_03555_),
    .Y(_03556_));
 sky130_fd_sc_hd__a21bo_1 _10645_ (.A1(_03418_),
    .A2(_03420_),
    .B1_N(_03422_),
    .X(_03557_));
 sky130_fd_sc_hd__a21bo_1 _10646_ (.A1(_03450_),
    .A2(_03456_),
    .B1_N(_03455_),
    .X(_03558_));
 sky130_fd_sc_hd__o22a_1 _10647_ (.A1(net69),
    .A2(_00811_),
    .B1(net10),
    .B2(_00497_),
    .X(_03559_));
 sky130_fd_sc_hd__xnor2_1 _10648_ (.A(net145),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__nand2_1 _10649_ (.A(_00224_),
    .B(net6),
    .Y(_03561_));
 sky130_fd_sc_hd__a22o_1 _10650_ (.A1(_00226_),
    .A2(net6),
    .B1(_03561_),
    .B2(net155),
    .X(_03562_));
 sky130_fd_sc_hd__nor2_1 _10651_ (.A(_03560_),
    .B(_03562_),
    .Y(_03563_));
 sky130_fd_sc_hd__xor2_1 _10652_ (.A(_03560_),
    .B(_03562_),
    .X(_03564_));
 sky130_fd_sc_hd__a21oi_1 _10653_ (.A1(_03455_),
    .A2(_03457_),
    .B1(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__xnor2_1 _10654_ (.A(_03558_),
    .B(_03564_),
    .Y(_03566_));
 sky130_fd_sc_hd__and2_1 _10655_ (.A(_03557_),
    .B(_03566_),
    .X(_03567_));
 sky130_fd_sc_hd__xnor2_1 _10656_ (.A(_03557_),
    .B(_03566_),
    .Y(_03568_));
 sky130_fd_sc_hd__a22o_1 _10657_ (.A1(net15),
    .A2(net73),
    .B1(net71),
    .B2(net31),
    .X(_03569_));
 sky130_fd_sc_hd__xnor2_1 _10658_ (.A(net92),
    .B(_03569_),
    .Y(_03570_));
 sky130_fd_sc_hd__o22a_1 _10659_ (.A1(_00219_),
    .A2(net39),
    .B1(net36),
    .B2(net100),
    .X(_03571_));
 sky130_fd_sc_hd__xnor2_1 _10660_ (.A(_00262_),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__o22a_1 _10661_ (.A1(net34),
    .A2(net82),
    .B1(net77),
    .B2(net32),
    .X(_03573_));
 sky130_fd_sc_hd__xnor2_1 _10662_ (.A(net94),
    .B(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__nand2_1 _10663_ (.A(_03572_),
    .B(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__or2_1 _10664_ (.A(_03572_),
    .B(_03574_),
    .X(_03576_));
 sky130_fd_sc_hd__nand2_1 _10665_ (.A(_03575_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__xnor2_1 _10666_ (.A(_03570_),
    .B(_03577_),
    .Y(_03578_));
 sky130_fd_sc_hd__or2_1 _10667_ (.A(_03568_),
    .B(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__xnor2_1 _10668_ (.A(_03568_),
    .B(_03578_),
    .Y(_03580_));
 sky130_fd_sc_hd__xor2_1 _10669_ (.A(_03556_),
    .B(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__o21ai_2 _10670_ (.A1(_03402_),
    .A2(_03409_),
    .B1(_03407_),
    .Y(_03582_));
 sky130_fd_sc_hd__o22a_1 _10671_ (.A1(net50),
    .A2(net84),
    .B1(net80),
    .B2(net51),
    .X(_03583_));
 sky130_fd_sc_hd__xnor2_1 _10672_ (.A(net117),
    .B(_03583_),
    .Y(_03584_));
 sky130_fd_sc_hd__o32a_1 _10673_ (.A1(_00466_),
    .A2(_00513_),
    .A3(_00515_),
    .B1(_00460_),
    .B2(net43),
    .X(_03585_));
 sky130_fd_sc_hd__xnor2_1 _10674_ (.A(net109),
    .B(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__nand2_1 _10675_ (.A(_03584_),
    .B(_03586_),
    .Y(_03587_));
 sky130_fd_sc_hd__or2_1 _10676_ (.A(_03584_),
    .B(_03586_),
    .X(_03588_));
 sky130_fd_sc_hd__nand2_1 _10677_ (.A(_03587_),
    .B(_03588_),
    .Y(_03589_));
 sky130_fd_sc_hd__a21oi_2 _10678_ (.A1(_03443_),
    .A2(_03445_),
    .B1(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__and3_1 _10679_ (.A(_03443_),
    .B(_03445_),
    .C(_03589_),
    .X(_03591_));
 sky130_fd_sc_hd__or2_1 _10680_ (.A(_03590_),
    .B(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__and2b_1 _10681_ (.A_N(_03592_),
    .B(_03582_),
    .X(_03593_));
 sky130_fd_sc_hd__xnor2_1 _10682_ (.A(_03582_),
    .B(_03592_),
    .Y(_03594_));
 sky130_fd_sc_hd__nand2_1 _10683_ (.A(_03581_),
    .B(_03594_),
    .Y(_03595_));
 sky130_fd_sc_hd__or2_1 _10684_ (.A(_03581_),
    .B(_03594_),
    .X(_03596_));
 sky130_fd_sc_hd__nand2_1 _10685_ (.A(_03595_),
    .B(_03596_),
    .Y(_03597_));
 sky130_fd_sc_hd__nand2_1 _10686_ (.A(_03459_),
    .B(_03461_),
    .Y(_03598_));
 sky130_fd_sc_hd__a21o_1 _10687_ (.A1(_03434_),
    .A2(_03435_),
    .B1(_03432_),
    .X(_03599_));
 sky130_fd_sc_hd__o22a_1 _10688_ (.A1(net57),
    .A2(net29),
    .B1(net27),
    .B2(net54),
    .X(_03600_));
 sky130_fd_sc_hd__xnor2_1 _10689_ (.A(net89),
    .B(_03600_),
    .Y(_03601_));
 sky130_fd_sc_hd__inv_2 _10690_ (.A(_03601_),
    .Y(_03602_));
 sky130_fd_sc_hd__o22a_1 _10691_ (.A1(net48),
    .A2(net25),
    .B1(net23),
    .B2(net46),
    .X(_03603_));
 sky130_fd_sc_hd__xnor2_1 _10692_ (.A(net87),
    .B(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__o22a_1 _10693_ (.A1(net42),
    .A2(net20),
    .B1(net18),
    .B2(net41),
    .X(_03605_));
 sky130_fd_sc_hd__xnor2_1 _10694_ (.A(net97),
    .B(_03605_),
    .Y(_03606_));
 sky130_fd_sc_hd__nand2_1 _10695_ (.A(_03604_),
    .B(_03606_),
    .Y(_03607_));
 sky130_fd_sc_hd__or2_1 _10696_ (.A(_03604_),
    .B(_03606_),
    .X(_03608_));
 sky130_fd_sc_hd__nand2_1 _10697_ (.A(_03607_),
    .B(_03608_),
    .Y(_03609_));
 sky130_fd_sc_hd__or2_1 _10698_ (.A(_03602_),
    .B(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__nand2_1 _10699_ (.A(_03602_),
    .B(_03609_),
    .Y(_03611_));
 sky130_fd_sc_hd__nand2_1 _10700_ (.A(_03610_),
    .B(_03611_),
    .Y(_03612_));
 sky130_fd_sc_hd__and3_1 _10701_ (.A(_03599_),
    .B(_03610_),
    .C(_03611_),
    .X(_03613_));
 sky130_fd_sc_hd__xnor2_1 _10702_ (.A(_03599_),
    .B(_03612_),
    .Y(_03614_));
 sky130_fd_sc_hd__xnor2_1 _10703_ (.A(_03598_),
    .B(_03614_),
    .Y(_03615_));
 sky130_fd_sc_hd__xor2_1 _10704_ (.A(_03597_),
    .B(_03615_),
    .X(_03616_));
 sky130_fd_sc_hd__o21ba_1 _10705_ (.A1(_03413_),
    .A2(_03468_),
    .B1_N(_03467_),
    .X(_03617_));
 sky130_fd_sc_hd__a21bo_1 _10706_ (.A1(_03399_),
    .A2(_03412_),
    .B1_N(_03411_),
    .X(_03618_));
 sky130_fd_sc_hd__a31oi_2 _10707_ (.A1(_03422_),
    .A2(_03423_),
    .A3(_03425_),
    .B1(_03427_),
    .Y(_03619_));
 sky130_fd_sc_hd__o21ba_1 _10708_ (.A1(_03436_),
    .A2(_03464_),
    .B1_N(_03463_),
    .X(_03620_));
 sky130_fd_sc_hd__nor2_1 _10709_ (.A(_03619_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__xor2_1 _10710_ (.A(_03619_),
    .B(_03620_),
    .X(_03622_));
 sky130_fd_sc_hd__xnor2_1 _10711_ (.A(_03618_),
    .B(_03622_),
    .Y(_03623_));
 sky130_fd_sc_hd__a21oi_1 _10712_ (.A1(_03473_),
    .A2(_03477_),
    .B1(_03476_),
    .Y(_03624_));
 sky130_fd_sc_hd__xor2_1 _10713_ (.A(_03623_),
    .B(_03624_),
    .X(_03625_));
 sky130_fd_sc_hd__nand2b_1 _10714_ (.A_N(_03617_),
    .B(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__xnor2_1 _10715_ (.A(_03617_),
    .B(_03625_),
    .Y(_03627_));
 sky130_fd_sc_hd__nand2_1 _10716_ (.A(_03616_),
    .B(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__xnor2_1 _10717_ (.A(_03616_),
    .B(_03627_),
    .Y(_03629_));
 sky130_fd_sc_hd__a21o_1 _10718_ (.A1(_03479_),
    .A2(_03481_),
    .B1(_03629_),
    .X(_03630_));
 sky130_fd_sc_hd__nand3_1 _10719_ (.A(_03479_),
    .B(_03481_),
    .C(_03629_),
    .Y(_03631_));
 sky130_fd_sc_hd__and2_2 _10720_ (.A(_03630_),
    .B(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__nand2_1 _10721_ (.A(_03546_),
    .B(_03632_),
    .Y(_03633_));
 sky130_fd_sc_hd__nor2_1 _10722_ (.A(_03546_),
    .B(_03632_),
    .Y(_03634_));
 sky130_fd_sc_hd__xnor2_4 _10723_ (.A(_03546_),
    .B(_03632_),
    .Y(_03635_));
 sky130_fd_sc_hd__xor2_4 _10724_ (.A(_03545_),
    .B(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__a2111o_1 _10725_ (.A1(_03353_),
    .A2(_03354_),
    .B1(_02241_),
    .C1(_03070_),
    .D1(_03071_),
    .X(_03637_));
 sky130_fd_sc_hd__or4b_1 _10726_ (.A(_02347_),
    .B(_02748_),
    .C(_02908_),
    .D_N(_02574_),
    .X(_03638_));
 sky130_fd_sc_hd__or4_2 _10727_ (.A(_03218_),
    .B(_03496_),
    .C(_03637_),
    .D(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__a21o_1 _10728_ (.A1(net137),
    .A2(_03639_),
    .B1(_03636_),
    .X(_03640_));
 sky130_fd_sc_hd__and3_1 _10729_ (.A(net137),
    .B(_03636_),
    .C(_03639_),
    .X(_03641_));
 sky130_fd_sc_hd__and3b_1 _10730_ (.A_N(_03641_),
    .B(_02348_),
    .C(_03640_),
    .X(_03642_));
 sky130_fd_sc_hd__or3_1 _10731_ (.A(net134),
    .B(_01938_),
    .C(_01939_),
    .X(_03643_));
 sky130_fd_sc_hd__o21ai_1 _10732_ (.A1(net134),
    .A2(_01938_),
    .B1(_01939_),
    .Y(_03644_));
 sky130_fd_sc_hd__o31a_1 _10733_ (.A1(_06525_),
    .A2(_06532_),
    .A3(_03502_),
    .B1(_06526_),
    .X(_03645_));
 sky130_fd_sc_hd__nor2_1 _10734_ (.A(net295),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__a31o_1 _10735_ (.A1(net295),
    .A2(_06524_),
    .A3(_06585_),
    .B1(_03646_),
    .X(_03647_));
 sky130_fd_sc_hd__nand2_1 _10736_ (.A(_06521_),
    .B(_03647_),
    .Y(_03648_));
 sky130_fd_sc_hd__o211a_1 _10737_ (.A1(_06521_),
    .A2(_03647_),
    .B1(_03648_),
    .C1(net234),
    .X(_03649_));
 sky130_fd_sc_hd__o21a_1 _10738_ (.A1(_03529_),
    .A2(_03530_),
    .B1(_03531_),
    .X(_03650_));
 sky130_fd_sc_hd__nor2_1 _10739_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03651_));
 sky130_fd_sc_hd__nand2_1 _10740_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03652_));
 sky130_fd_sc_hd__nand2b_1 _10741_ (.A_N(_03651_),
    .B(_03652_),
    .Y(_03653_));
 sky130_fd_sc_hd__xor2_1 _10742_ (.A(_03650_),
    .B(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__mux2_1 _10743_ (.A0(_02386_),
    .A1(_02401_),
    .S(net219),
    .X(_03655_));
 sky130_fd_sc_hd__mux2_2 _10744_ (.A0(_03508_),
    .A1(_03655_),
    .S(net220),
    .X(_03656_));
 sky130_fd_sc_hd__mux2_1 _10745_ (.A0(_03654_),
    .A1(_03656_),
    .S(net223),
    .X(_03657_));
 sky130_fd_sc_hd__nor2_1 _10746_ (.A(\div_res[7] ),
    .B(_03517_),
    .Y(_03658_));
 sky130_fd_sc_hd__o21bai_1 _10747_ (.A1(_06681_),
    .A2(_03658_),
    .B1_N(\div_res[8] ),
    .Y(_03659_));
 sky130_fd_sc_hd__or3b_1 _10748_ (.A(_03658_),
    .B(_06681_),
    .C_N(\div_res[8] ),
    .X(_03660_));
 sky130_fd_sc_hd__a21oi_1 _10749_ (.A1(_06520_),
    .A2(net195),
    .B1(net193),
    .Y(_03661_));
 sky130_fd_sc_hd__nand3_1 _10750_ (.A(_00212_),
    .B(_00222_),
    .C(net256),
    .Y(_03662_));
 sky130_fd_sc_hd__o221a_1 _10751_ (.A1(_06517_),
    .A2(net203),
    .B1(net231),
    .B2(reg1_val[8]),
    .C1(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__or2_1 _10752_ (.A(\div_shifter[39] ),
    .B(_03523_),
    .X(_03664_));
 sky130_fd_sc_hd__a21oi_2 _10753_ (.A1(net227),
    .A2(_03664_),
    .B1(\div_shifter[40] ),
    .Y(_03665_));
 sky130_fd_sc_hd__a31o_1 _10754_ (.A1(\div_shifter[40] ),
    .A2(net227),
    .A3(_03664_),
    .B1(net191),
    .X(_03666_));
 sky130_fd_sc_hd__o22a_1 _10755_ (.A1(_06520_),
    .A2(net194),
    .B1(_03665_),
    .B2(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__o211ai_1 _10756_ (.A1(_06519_),
    .A2(_03661_),
    .B1(_03663_),
    .C1(_03667_),
    .Y(_03668_));
 sky130_fd_sc_hd__a31o_1 _10757_ (.A1(_02443_),
    .A2(_03659_),
    .A3(_03660_),
    .B1(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__o21a_1 _10758_ (.A1(net222),
    .A2(_03515_),
    .B1(_02456_),
    .X(_03670_));
 sky130_fd_sc_hd__a221o_1 _10759_ (.A1(net167),
    .A2(_03656_),
    .B1(_03670_),
    .B2(net171),
    .C1(_03669_),
    .X(_03671_));
 sky130_fd_sc_hd__a211o_1 _10760_ (.A1(net205),
    .A2(_03657_),
    .B1(_03671_),
    .C1(_03649_),
    .X(_03672_));
 sky130_fd_sc_hd__a311o_1 _10761_ (.A1(net233),
    .A2(_03643_),
    .A3(_03644_),
    .B1(_03672_),
    .C1(_03642_),
    .X(_03673_));
 sky130_fd_sc_hd__a31o_1 _10762_ (.A1(curr_PC[6]),
    .A2(curr_PC[7]),
    .A3(_03255_),
    .B1(curr_PC[8]),
    .X(_03674_));
 sky130_fd_sc_hd__and3_2 _10763_ (.A(curr_PC[7]),
    .B(curr_PC[8]),
    .C(_03394_),
    .X(_03675_));
 sky130_fd_sc_hd__nor2_1 _10764_ (.A(net237),
    .B(_03675_),
    .Y(_03676_));
 sky130_fd_sc_hd__a22o_4 _10765_ (.A1(net237),
    .A2(_03673_),
    .B1(_03674_),
    .B2(_03676_),
    .X(dest_val[8]));
 sky130_fd_sc_hd__xnor2_2 _10766_ (.A(curr_PC[9]),
    .B(_03675_),
    .Y(_03677_));
 sky130_fd_sc_hd__nor2_1 _10767_ (.A(_03636_),
    .B(_03639_),
    .Y(_03678_));
 sky130_fd_sc_hd__o21ai_1 _10768_ (.A1(_03623_),
    .A2(_03624_),
    .B1(_03626_),
    .Y(_03679_));
 sky130_fd_sc_hd__o22a_1 _10769_ (.A1(net46),
    .A2(net25),
    .B1(net23),
    .B2(net50),
    .X(_03680_));
 sky130_fd_sc_hd__xnor2_2 _10770_ (.A(_00359_),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__o22a_1 _10771_ (.A1(net51),
    .A2(net84),
    .B1(net79),
    .B2(net43),
    .X(_03682_));
 sky130_fd_sc_hd__xnor2_1 _10772_ (.A(net117),
    .B(_03682_),
    .Y(_03683_));
 sky130_fd_sc_hd__o22a_1 _10773_ (.A1(net54),
    .A2(net29),
    .B1(net27),
    .B2(net48),
    .X(_03684_));
 sky130_fd_sc_hd__xnor2_1 _10774_ (.A(net89),
    .B(_03684_),
    .Y(_03685_));
 sky130_fd_sc_hd__nand2_1 _10775_ (.A(_03683_),
    .B(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__or2_1 _10776_ (.A(_03683_),
    .B(_03685_),
    .X(_03687_));
 sky130_fd_sc_hd__nand2_1 _10777_ (.A(_03686_),
    .B(_03687_),
    .Y(_03688_));
 sky130_fd_sc_hd__xnor2_1 _10778_ (.A(_03681_),
    .B(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__a21oi_1 _10779_ (.A1(_03552_),
    .A2(_03554_),
    .B1(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__and3_1 _10780_ (.A(_03552_),
    .B(_03554_),
    .C(_03689_),
    .X(_03691_));
 sky130_fd_sc_hd__or2_1 _10781_ (.A(_03690_),
    .B(_03691_),
    .X(_03692_));
 sky130_fd_sc_hd__o21ba_1 _10782_ (.A1(_03565_),
    .A2(_03567_),
    .B1_N(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__or3b_1 _10783_ (.A(_03565_),
    .B(_03567_),
    .C_N(_03692_),
    .X(_03694_));
 sky130_fd_sc_hd__and2b_1 _10784_ (.A_N(_03693_),
    .B(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__o22a_1 _10785_ (.A1(net69),
    .A2(net10),
    .B1(net5),
    .B2(net67),
    .X(_03696_));
 sky130_fd_sc_hd__xnor2_2 _10786_ (.A(net145),
    .B(_03696_),
    .Y(_03697_));
 sky130_fd_sc_hd__or3_1 _10787_ (.A(_00460_),
    .B(_00513_),
    .C(_00515_),
    .X(_03698_));
 sky130_fd_sc_hd__a21o_1 _10788_ (.A1(_00809_),
    .A2(_00810_),
    .B1(_00466_),
    .X(_03699_));
 sky130_fd_sc_hd__a21o_1 _10789_ (.A1(_03698_),
    .A2(_03699_),
    .B1(_00431_),
    .X(_03700_));
 sky130_fd_sc_hd__nand3_1 _10790_ (.A(_00431_),
    .B(_03698_),
    .C(_03699_),
    .Y(_03701_));
 sky130_fd_sc_hd__and3b_1 _10791_ (.A_N(net155),
    .B(_03700_),
    .C(_03701_),
    .X(_03702_));
 sky130_fd_sc_hd__a21bo_1 _10792_ (.A1(_03700_),
    .A2(_03701_),
    .B1_N(net155),
    .X(_03703_));
 sky130_fd_sc_hd__and2b_1 _10793_ (.A_N(_03702_),
    .B(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__xnor2_2 _10794_ (.A(_03697_),
    .B(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__o21a_1 _10795_ (.A1(_03570_),
    .A2(_03577_),
    .B1(_03575_),
    .X(_03706_));
 sky130_fd_sc_hd__xnor2_1 _10796_ (.A(_03705_),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__a21oi_1 _10797_ (.A1(_03607_),
    .A2(_03610_),
    .B1(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__and3_1 _10798_ (.A(_03607_),
    .B(_03610_),
    .C(_03707_),
    .X(_03709_));
 sky130_fd_sc_hd__a22o_1 _10799_ (.A1(_00443_),
    .A2(net16),
    .B1(net12),
    .B2(_00397_),
    .X(_03710_));
 sky130_fd_sc_hd__xnor2_1 _10800_ (.A(net64),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__inv_2 _10801_ (.A(_03711_),
    .Y(_03712_));
 sky130_fd_sc_hd__a22o_1 _10802_ (.A1(_00392_),
    .A2(net8),
    .B1(net4),
    .B2(_00375_),
    .X(_03713_));
 sky130_fd_sc_hd__xnor2_1 _10803_ (.A(net59),
    .B(_03713_),
    .Y(_03714_));
 sky130_fd_sc_hd__o22a_1 _10804_ (.A1(net34),
    .A2(net77),
    .B1(_00463_),
    .B2(net32),
    .X(_03715_));
 sky130_fd_sc_hd__xnor2_1 _10805_ (.A(net94),
    .B(_03715_),
    .Y(_03716_));
 sky130_fd_sc_hd__xnor2_1 _10806_ (.A(_03714_),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__or2_1 _10807_ (.A(_03712_),
    .B(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__nand2_1 _10808_ (.A(_03712_),
    .B(_03717_),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_1 _10809_ (.A(_03718_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__nand2_1 _10810_ (.A(net122),
    .B(net62),
    .Y(_03721_));
 sky130_fd_sc_hd__xor2_1 _10811_ (.A(_03587_),
    .B(_03721_),
    .X(_03722_));
 sky130_fd_sc_hd__nand2b_1 _10812_ (.A_N(_03563_),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__xnor2_1 _10813_ (.A(_03563_),
    .B(_03722_),
    .Y(_03724_));
 sky130_fd_sc_hd__o22a_1 _10814_ (.A1(net100),
    .A2(net38),
    .B1(net36),
    .B2(net42),
    .X(_03725_));
 sky130_fd_sc_hd__xnor2_1 _10815_ (.A(_00263_),
    .B(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__o22a_1 _10816_ (.A1(_00219_),
    .A2(_00342_),
    .B1(net70),
    .B2(_00336_),
    .X(_03727_));
 sky130_fd_sc_hd__xnor2_1 _10817_ (.A(net92),
    .B(_03727_),
    .Y(_03728_));
 sky130_fd_sc_hd__o22a_1 _10818_ (.A1(net41),
    .A2(net20),
    .B1(net18),
    .B2(net57),
    .X(_03729_));
 sky130_fd_sc_hd__xnor2_1 _10819_ (.A(_00273_),
    .B(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__nand2_1 _10820_ (.A(_03728_),
    .B(_03730_),
    .Y(_03731_));
 sky130_fd_sc_hd__xnor2_1 _10821_ (.A(_03728_),
    .B(_03730_),
    .Y(_03732_));
 sky130_fd_sc_hd__or2_1 _10822_ (.A(_03726_),
    .B(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__nand2_1 _10823_ (.A(_03726_),
    .B(_03732_),
    .Y(_03734_));
 sky130_fd_sc_hd__and2_1 _10824_ (.A(_03733_),
    .B(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__and2_1 _10825_ (.A(_03724_),
    .B(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__inv_2 _10826_ (.A(_03736_),
    .Y(_03737_));
 sky130_fd_sc_hd__nor2_1 _10827_ (.A(_03724_),
    .B(_03735_),
    .Y(_03738_));
 sky130_fd_sc_hd__or3_1 _10828_ (.A(_03720_),
    .B(_03736_),
    .C(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__o21ai_1 _10829_ (.A1(_03736_),
    .A2(_03738_),
    .B1(_03720_),
    .Y(_03740_));
 sky130_fd_sc_hd__or4bb_1 _10830_ (.A(_03708_),
    .B(_03709_),
    .C_N(_03739_),
    .D_N(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__a2bb2o_1 _10831_ (.A1_N(_03708_),
    .A2_N(_03709_),
    .B1(_03739_),
    .B2(_03740_),
    .X(_03742_));
 sky130_fd_sc_hd__and3_1 _10832_ (.A(_03695_),
    .B(_03741_),
    .C(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__a21oi_1 _10833_ (.A1(_03741_),
    .A2(_03742_),
    .B1(_03695_),
    .Y(_03744_));
 sky130_fd_sc_hd__nor2_1 _10834_ (.A(_03743_),
    .B(_03744_),
    .Y(_03745_));
 sky130_fd_sc_hd__o21ai_1 _10835_ (.A1(_03597_),
    .A2(_03615_),
    .B1(_03595_),
    .Y(_03746_));
 sky130_fd_sc_hd__a21o_1 _10836_ (.A1(_03598_),
    .A2(_03614_),
    .B1(_03613_),
    .X(_03747_));
 sky130_fd_sc_hd__o21ai_1 _10837_ (.A1(_03556_),
    .A2(_03580_),
    .B1(_03579_),
    .Y(_03748_));
 sky130_fd_sc_hd__nor2_1 _10838_ (.A(_03590_),
    .B(_03593_),
    .Y(_03749_));
 sky130_fd_sc_hd__o21a_1 _10839_ (.A1(_03590_),
    .A2(_03593_),
    .B1(_03748_),
    .X(_03750_));
 sky130_fd_sc_hd__xnor2_1 _10840_ (.A(_03748_),
    .B(_03749_),
    .Y(_03751_));
 sky130_fd_sc_hd__xnor2_1 _10841_ (.A(_03747_),
    .B(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__a21oi_1 _10842_ (.A1(_03618_),
    .A2(_03622_),
    .B1(_03621_),
    .Y(_03753_));
 sky130_fd_sc_hd__xnor2_1 _10843_ (.A(_03752_),
    .B(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__nand2b_1 _10844_ (.A_N(_03754_),
    .B(_03746_),
    .Y(_03755_));
 sky130_fd_sc_hd__xnor2_1 _10845_ (.A(_03746_),
    .B(_03754_),
    .Y(_03756_));
 sky130_fd_sc_hd__nand2_1 _10846_ (.A(_03745_),
    .B(_03756_),
    .Y(_03757_));
 sky130_fd_sc_hd__xnor2_1 _10847_ (.A(_03745_),
    .B(_03756_),
    .Y(_03758_));
 sky130_fd_sc_hd__nand2b_1 _10848_ (.A_N(_03758_),
    .B(_03679_),
    .Y(_03759_));
 sky130_fd_sc_hd__xor2_1 _10849_ (.A(_03679_),
    .B(_03758_),
    .X(_03760_));
 sky130_fd_sc_hd__a21oi_1 _10850_ (.A1(_03628_),
    .A2(_03630_),
    .B1(_03760_),
    .Y(_03761_));
 sky130_fd_sc_hd__a21o_1 _10851_ (.A1(_03628_),
    .A2(_03630_),
    .B1(_03760_),
    .X(_03762_));
 sky130_fd_sc_hd__and3_1 _10852_ (.A(_03628_),
    .B(_03630_),
    .C(_03760_),
    .X(_03763_));
 sky130_fd_sc_hd__or2_4 _10853_ (.A(_03761_),
    .B(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__a21oi_2 _10854_ (.A1(_03486_),
    .A2(_03633_),
    .B1(_03634_),
    .Y(_03765_));
 sky130_fd_sc_hd__nor2_1 _10855_ (.A(_03488_),
    .B(_03635_),
    .Y(_03766_));
 sky130_fd_sc_hd__a21oi_1 _10856_ (.A1(_03493_),
    .A2(_03766_),
    .B1(_03765_),
    .Y(_03767_));
 sky130_fd_sc_hd__or4_1 _10857_ (.A(_03211_),
    .B(_03346_),
    .C(_03488_),
    .D(_03635_),
    .X(_03768_));
 sky130_fd_sc_hd__a211o_1 _10858_ (.A1(_02570_),
    .A2(_02572_),
    .B1(_03213_),
    .C1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__o211a_4 _10859_ (.A1(_03216_),
    .A2(_03768_),
    .B1(_03769_),
    .C1(_03767_),
    .X(_03770_));
 sky130_fd_sc_hd__xnor2_4 _10860_ (.A(_03764_),
    .B(_03770_),
    .Y(_03771_));
 sky130_fd_sc_hd__o21ai_1 _10861_ (.A1(net134),
    .A2(_03678_),
    .B1(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__or3_1 _10862_ (.A(net135),
    .B(_03678_),
    .C(_03771_),
    .X(_03773_));
 sky130_fd_sc_hd__nand2_1 _10863_ (.A(_03772_),
    .B(_03773_),
    .Y(_03774_));
 sky130_fd_sc_hd__or3_1 _10864_ (.A(net134),
    .B(_01940_),
    .C(_01941_),
    .X(_03775_));
 sky130_fd_sc_hd__o21a_1 _10865_ (.A1(net134),
    .A2(_01940_),
    .B1(_01941_),
    .X(_03776_));
 sky130_fd_sc_hd__or3b_1 _10866_ (.A(_03776_),
    .B(_02434_),
    .C_N(_03775_),
    .X(_03777_));
 sky130_fd_sc_hd__or3_1 _10867_ (.A(net283),
    .B(_06518_),
    .C(_06586_),
    .X(_03778_));
 sky130_fd_sc_hd__o21a_1 _10868_ (.A1(_06519_),
    .A2(_03645_),
    .B1(_06520_),
    .X(_03779_));
 sky130_fd_sc_hd__o21a_1 _10869_ (.A1(net295),
    .A2(_03779_),
    .B1(_03778_),
    .X(_03780_));
 sky130_fd_sc_hd__nor2_1 _10870_ (.A(_06514_),
    .B(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__a211o_1 _10871_ (.A1(_06514_),
    .A2(_03780_),
    .B1(_03781_),
    .C1(_02427_),
    .X(_03782_));
 sky130_fd_sc_hd__o21a_1 _10872_ (.A1(_03650_),
    .A2(_03651_),
    .B1(_03652_),
    .X(_03783_));
 sky130_fd_sc_hd__nor2_1 _10873_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03784_));
 sky130_fd_sc_hd__nand2_1 _10874_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03785_));
 sky130_fd_sc_hd__nand2b_1 _10875_ (.A_N(_03784_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__xor2_1 _10876_ (.A(_03783_),
    .B(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(_02595_),
    .A1(_02603_),
    .S(net219),
    .X(_03788_));
 sky130_fd_sc_hd__mux2_2 _10878_ (.A0(_03365_),
    .A1(_03788_),
    .S(net220),
    .X(_03789_));
 sky130_fd_sc_hd__inv_2 _10879_ (.A(_03789_),
    .Y(_03790_));
 sky130_fd_sc_hd__nor2_1 _10880_ (.A(net223),
    .B(_03787_),
    .Y(_03791_));
 sky130_fd_sc_hd__a211o_1 _10881_ (.A1(net223),
    .A2(_03790_),
    .B1(_03791_),
    .C1(_06667_),
    .X(_03792_));
 sky130_fd_sc_hd__or3_1 _10882_ (.A(\div_res[8] ),
    .B(\div_res[7] ),
    .C(_03517_),
    .X(_03793_));
 sky130_fd_sc_hd__a21oi_1 _10883_ (.A1(net139),
    .A2(_03793_),
    .B1(\div_res[9] ),
    .Y(_03794_));
 sky130_fd_sc_hd__a311o_1 _10884_ (.A1(\div_res[9] ),
    .A2(net139),
    .A3(_03793_),
    .B1(_03794_),
    .C1(net189),
    .X(_03795_));
 sky130_fd_sc_hd__or2_1 _10885_ (.A(\div_shifter[40] ),
    .B(_03664_),
    .X(_03796_));
 sky130_fd_sc_hd__a21oi_1 _10886_ (.A1(net228),
    .A2(_03796_),
    .B1(\div_shifter[41] ),
    .Y(_03797_));
 sky130_fd_sc_hd__a31o_1 _10887_ (.A1(\div_shifter[41] ),
    .A2(net227),
    .A3(_03796_),
    .B1(net191),
    .X(_03798_));
 sky130_fd_sc_hd__or2_1 _10888_ (.A(_03797_),
    .B(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__nand2_1 _10889_ (.A(_06509_),
    .B(_06677_),
    .Y(_03800_));
 sky130_fd_sc_hd__o211a_1 _10890_ (.A1(reg1_val[9]),
    .A2(net232),
    .B1(_03800_),
    .C1(net241),
    .X(_03801_));
 sky130_fd_sc_hd__a22o_1 _10891_ (.A1(_06513_),
    .A2(net195),
    .B1(net257),
    .B2(_00214_),
    .X(_03802_));
 sky130_fd_sc_hd__o221a_1 _10892_ (.A1(_06512_),
    .A2(net194),
    .B1(_02440_),
    .B2(_06511_),
    .C1(_03801_),
    .X(_03803_));
 sky130_fd_sc_hd__and4b_1 _10893_ (.A_N(_03802_),
    .B(_03803_),
    .C(_03795_),
    .D(_03799_),
    .X(_03804_));
 sky130_fd_sc_hd__o21ai_2 _10894_ (.A1(net221),
    .A2(_03371_),
    .B1(_02456_),
    .Y(_03805_));
 sky130_fd_sc_hd__inv_2 _10895_ (.A(_03805_),
    .Y(_03806_));
 sky130_fd_sc_hd__o221a_1 _10896_ (.A1(_02425_),
    .A2(_03790_),
    .B1(_03805_),
    .B2(net169),
    .C1(_03804_),
    .X(_03807_));
 sky130_fd_sc_hd__and3_1 _10897_ (.A(_03782_),
    .B(_03792_),
    .C(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__o211a_1 _10898_ (.A1(net235),
    .A2(_03774_),
    .B1(_03777_),
    .C1(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__a21oi_4 _10899_ (.A1(net242),
    .A2(_03677_),
    .B1(_03809_),
    .Y(dest_val[9]));
 sky130_fd_sc_hd__nand2_1 _10900_ (.A(_03678_),
    .B(_03771_),
    .Y(_03810_));
 sky130_fd_sc_hd__o21ai_1 _10901_ (.A1(_03752_),
    .A2(_03753_),
    .B1(_03755_),
    .Y(_03811_));
 sky130_fd_sc_hd__o22a_1 _10902_ (.A1(net34),
    .A2(_00463_),
    .B1(_00468_),
    .B2(net32),
    .X(_03812_));
 sky130_fd_sc_hd__xnor2_1 _10903_ (.A(_00302_),
    .B(_03812_),
    .Y(_03813_));
 sky130_fd_sc_hd__a22o_1 _10904_ (.A1(net102),
    .A2(net15),
    .B1(net31),
    .B2(net101),
    .X(_03814_));
 sky130_fd_sc_hd__xnor2_1 _10905_ (.A(_00309_),
    .B(_03814_),
    .Y(_03815_));
 sky130_fd_sc_hd__a22o_1 _10906_ (.A1(_00446_),
    .A2(net16),
    .B1(net12),
    .B2(_00443_),
    .X(_03816_));
 sky130_fd_sc_hd__xnor2_1 _10907_ (.A(net64),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__nand2_1 _10908_ (.A(_03815_),
    .B(_03817_),
    .Y(_03818_));
 sky130_fd_sc_hd__xnor2_1 _10909_ (.A(_03815_),
    .B(_03817_),
    .Y(_03819_));
 sky130_fd_sc_hd__xnor2_1 _10910_ (.A(_03813_),
    .B(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21o_1 _10911_ (.A1(_03697_),
    .A2(_03703_),
    .B1(_03702_),
    .X(_03821_));
 sky130_fd_sc_hd__a22o_1 _10912_ (.A1(_00397_),
    .A2(net9),
    .B1(net4),
    .B2(_00392_),
    .X(_03822_));
 sky130_fd_sc_hd__xnor2_1 _10913_ (.A(net59),
    .B(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__xor2_1 _10914_ (.A(_03821_),
    .B(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__nor2_1 _10915_ (.A(net120),
    .B(net59),
    .Y(_03825_));
 sky130_fd_sc_hd__and2_1 _10916_ (.A(_03824_),
    .B(_03825_),
    .X(_03826_));
 sky130_fd_sc_hd__xnor2_1 _10917_ (.A(_03824_),
    .B(_03825_),
    .Y(_03827_));
 sky130_fd_sc_hd__o22a_1 _10918_ (.A1(net56),
    .A2(net20),
    .B1(net19),
    .B2(net53),
    .X(_03828_));
 sky130_fd_sc_hd__xnor2_1 _10919_ (.A(_00273_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__o22a_1 _10920_ (.A1(_00202_),
    .A2(net38),
    .B1(net36),
    .B2(net41),
    .X(_03830_));
 sky130_fd_sc_hd__xnor2_1 _10921_ (.A(net98),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__o22a_1 _10922_ (.A1(net48),
    .A2(net29),
    .B1(net27),
    .B2(net45),
    .X(_03832_));
 sky130_fd_sc_hd__xnor2_1 _10923_ (.A(net89),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__and2_1 _10924_ (.A(_03831_),
    .B(_03833_),
    .X(_03834_));
 sky130_fd_sc_hd__or2_1 _10925_ (.A(_03831_),
    .B(_03833_),
    .X(_03835_));
 sky130_fd_sc_hd__nand2b_1 _10926_ (.A_N(_03834_),
    .B(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__xor2_1 _10927_ (.A(_03829_),
    .B(_03836_),
    .X(_03837_));
 sky130_fd_sc_hd__nor2_1 _10928_ (.A(_03827_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__xnor2_1 _10929_ (.A(_03827_),
    .B(_03837_),
    .Y(_03839_));
 sky130_fd_sc_hd__nor2_1 _10930_ (.A(_03820_),
    .B(_03839_),
    .Y(_03840_));
 sky130_fd_sc_hd__and2_1 _10931_ (.A(_03820_),
    .B(_03839_),
    .X(_03841_));
 sky130_fd_sc_hd__nor2_1 _10932_ (.A(_03840_),
    .B(_03841_),
    .Y(_03842_));
 sky130_fd_sc_hd__o21ai_2 _10933_ (.A1(_03681_),
    .A2(_03688_),
    .B1(_03686_),
    .Y(_03843_));
 sky130_fd_sc_hd__nand2_1 _10934_ (.A(_00493_),
    .B(net6),
    .Y(_03844_));
 sky130_fd_sc_hd__a22o_2 _10935_ (.A1(_00495_),
    .A2(net6),
    .B1(_03844_),
    .B2(net145),
    .X(_03845_));
 sky130_fd_sc_hd__a21oi_1 _10936_ (.A1(_03731_),
    .A2(_03733_),
    .B1(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__and3_1 _10937_ (.A(_03731_),
    .B(_03733_),
    .C(_03845_),
    .X(_03847_));
 sky130_fd_sc_hd__nor2_1 _10938_ (.A(_03846_),
    .B(_03847_),
    .Y(_03848_));
 sky130_fd_sc_hd__xor2_2 _10939_ (.A(_03843_),
    .B(_03848_),
    .X(_03849_));
 sky130_fd_sc_hd__nand2_1 _10940_ (.A(_03842_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__xnor2_1 _10941_ (.A(_03842_),
    .B(_03849_),
    .Y(_03851_));
 sky130_fd_sc_hd__o21ai_2 _10942_ (.A1(_03587_),
    .A2(_03721_),
    .B1(_03723_),
    .Y(_03852_));
 sky130_fd_sc_hd__o22a_1 _10943_ (.A1(net43),
    .A2(net83),
    .B1(net79),
    .B2(_00517_),
    .X(_03853_));
 sky130_fd_sc_hd__xnor2_1 _10944_ (.A(_00381_),
    .B(_03853_),
    .Y(_03854_));
 sky130_fd_sc_hd__o22a_1 _10945_ (.A1(_00460_),
    .A2(_00811_),
    .B1(net10),
    .B2(_00466_),
    .X(_03855_));
 sky130_fd_sc_hd__xnor2_1 _10946_ (.A(net109),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__o22a_1 _10947_ (.A1(net49),
    .A2(net25),
    .B1(net23),
    .B2(net52),
    .X(_03857_));
 sky130_fd_sc_hd__xnor2_1 _10948_ (.A(net87),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__and2_1 _10949_ (.A(_03856_),
    .B(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__xnor2_1 _10950_ (.A(_03856_),
    .B(_03858_),
    .Y(_03860_));
 sky130_fd_sc_hd__nor2_1 _10951_ (.A(_03854_),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__and2_1 _10952_ (.A(_03854_),
    .B(_03860_),
    .X(_03862_));
 sky130_fd_sc_hd__or2_1 _10953_ (.A(_03861_),
    .B(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__a21bo_1 _10954_ (.A1(_03714_),
    .A2(_03716_),
    .B1_N(_03718_),
    .X(_03864_));
 sky130_fd_sc_hd__nand2b_1 _10955_ (.A_N(_03863_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__xor2_1 _10956_ (.A(_03863_),
    .B(_03864_),
    .X(_03866_));
 sky130_fd_sc_hd__nand2b_1 _10957_ (.A_N(_03866_),
    .B(_03852_),
    .Y(_03867_));
 sky130_fd_sc_hd__xor2_1 _10958_ (.A(_03852_),
    .B(_03866_),
    .X(_03868_));
 sky130_fd_sc_hd__xor2_1 _10959_ (.A(_03851_),
    .B(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__a21bo_1 _10960_ (.A1(_03695_),
    .A2(_03742_),
    .B1_N(_03741_),
    .X(_03870_));
 sky130_fd_sc_hd__a21o_1 _10961_ (.A1(_03747_),
    .A2(_03751_),
    .B1(_03750_),
    .X(_03871_));
 sky130_fd_sc_hd__or2_1 _10962_ (.A(_03690_),
    .B(_03693_),
    .X(_03872_));
 sky130_fd_sc_hd__o21bai_1 _10963_ (.A1(_03705_),
    .A2(_03706_),
    .B1_N(_03708_),
    .Y(_03873_));
 sky130_fd_sc_hd__and2_1 _10964_ (.A(_03737_),
    .B(_03739_),
    .X(_03874_));
 sky130_fd_sc_hd__a21bo_1 _10965_ (.A1(_03737_),
    .A2(_03739_),
    .B1_N(_03873_),
    .X(_03875_));
 sky130_fd_sc_hd__xnor2_1 _10966_ (.A(_03873_),
    .B(_03874_),
    .Y(_03876_));
 sky130_fd_sc_hd__xor2_1 _10967_ (.A(_03872_),
    .B(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__xnor2_1 _10968_ (.A(_03871_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__nand2b_1 _10969_ (.A_N(_03878_),
    .B(_03870_),
    .Y(_03879_));
 sky130_fd_sc_hd__xnor2_1 _10970_ (.A(_03870_),
    .B(_03878_),
    .Y(_03880_));
 sky130_fd_sc_hd__nand2_1 _10971_ (.A(_03869_),
    .B(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__xnor2_1 _10972_ (.A(_03869_),
    .B(_03880_),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2b_1 _10973_ (.A_N(_03882_),
    .B(_03811_),
    .Y(_03883_));
 sky130_fd_sc_hd__xor2_1 _10974_ (.A(_03811_),
    .B(_03882_),
    .X(_03884_));
 sky130_fd_sc_hd__a21o_1 _10975_ (.A1(_03757_),
    .A2(_03759_),
    .B1(_03884_),
    .X(_03885_));
 sky130_fd_sc_hd__nand3_2 _10976_ (.A(_03757_),
    .B(_03759_),
    .C(_03884_),
    .Y(_03886_));
 sky130_fd_sc_hd__nand2_4 _10977_ (.A(_03885_),
    .B(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__a21oi_2 _10978_ (.A1(_03633_),
    .A2(_03762_),
    .B1(_03763_),
    .Y(_03888_));
 sky130_fd_sc_hd__nor2_1 _10979_ (.A(_03635_),
    .B(_03764_),
    .Y(_03889_));
 sky130_fd_sc_hd__a21oi_1 _10980_ (.A1(_03540_),
    .A2(_03889_),
    .B1(_03888_),
    .Y(_03890_));
 sky130_fd_sc_hd__or4_1 _10981_ (.A(_03346_),
    .B(_03488_),
    .C(_03635_),
    .D(_03764_),
    .X(_03891_));
 sky130_fd_sc_hd__o21bai_1 _10982_ (.A1(_03350_),
    .A2(_03351_),
    .B1_N(_03891_),
    .Y(_03892_));
 sky130_fd_sc_hd__o311a_4 _10983_ (.A1(_02747_),
    .A2(_03347_),
    .A3(_03891_),
    .B1(_03892_),
    .C1(_03890_),
    .X(_03893_));
 sky130_fd_sc_hd__xor2_4 _10984_ (.A(_03887_),
    .B(_03893_),
    .X(_03894_));
 sky130_fd_sc_hd__a21o_1 _10985_ (.A1(net136),
    .A2(_03810_),
    .B1(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__a31oi_1 _10986_ (.A1(net136),
    .A2(_03810_),
    .A3(_03894_),
    .B1(net235),
    .Y(_03896_));
 sky130_fd_sc_hd__a21oi_1 _10987_ (.A1(_01940_),
    .A2(_01941_),
    .B1(net134),
    .Y(_03897_));
 sky130_fd_sc_hd__xnor2_1 _10988_ (.A(_01945_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__o21a_1 _10989_ (.A1(_06511_),
    .A2(_03779_),
    .B1(_06512_),
    .X(_03899_));
 sky130_fd_sc_hd__nor2_1 _10990_ (.A(net293),
    .B(_03899_),
    .Y(_03900_));
 sky130_fd_sc_hd__a31o_1 _10991_ (.A1(net293),
    .A2(_06510_),
    .A3(_06587_),
    .B1(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__nand2_1 _10992_ (.A(_06507_),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__o21a_1 _10993_ (.A1(_06507_),
    .A2(_03901_),
    .B1(net234),
    .X(_03903_));
 sky130_fd_sc_hd__or2_1 _10994_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03904_));
 sky130_fd_sc_hd__and2_1 _10995_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03905_));
 sky130_fd_sc_hd__nand2_1 _10996_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .Y(_03906_));
 sky130_fd_sc_hd__o21ai_1 _10997_ (.A1(_03783_),
    .A2(_03784_),
    .B1(_03785_),
    .Y(_03907_));
 sky130_fd_sc_hd__a21oi_1 _10998_ (.A1(_03904_),
    .A2(_03906_),
    .B1(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__and3_1 _10999_ (.A(_03904_),
    .B(_03906_),
    .C(_03907_),
    .X(_03909_));
 sky130_fd_sc_hd__mux2_1 _11000_ (.A0(_02763_),
    .A1(_02767_),
    .S(net218),
    .X(_03910_));
 sky130_fd_sc_hd__mux2_1 _11001_ (.A0(_03228_),
    .A1(_03910_),
    .S(net220),
    .X(_03911_));
 sky130_fd_sc_hd__o21ai_1 _11002_ (.A1(_03908_),
    .A2(_03909_),
    .B1(net244),
    .Y(_03912_));
 sky130_fd_sc_hd__o211a_1 _11003_ (.A1(net244),
    .A2(_03911_),
    .B1(_03912_),
    .C1(net205),
    .X(_03913_));
 sky130_fd_sc_hd__or2_1 _11004_ (.A(\div_res[9] ),
    .B(_03793_),
    .X(_03914_));
 sky130_fd_sc_hd__a21oi_1 _11005_ (.A1(net139),
    .A2(_03914_),
    .B1(\div_res[10] ),
    .Y(_03915_));
 sky130_fd_sc_hd__a311o_1 _11006_ (.A1(\div_res[10] ),
    .A2(net139),
    .A3(_03914_),
    .B1(_03915_),
    .C1(net189),
    .X(_03916_));
 sky130_fd_sc_hd__or2_1 _11007_ (.A(\div_shifter[41] ),
    .B(_03796_),
    .X(_03917_));
 sky130_fd_sc_hd__a21oi_1 _11008_ (.A1(net228),
    .A2(_03917_),
    .B1(\div_shifter[42] ),
    .Y(_03918_));
 sky130_fd_sc_hd__a311o_1 _11009_ (.A1(\div_shifter[42] ),
    .A2(net228),
    .A3(_03917_),
    .B1(_03918_),
    .C1(net191),
    .X(_03919_));
 sky130_fd_sc_hd__nand2_1 _11010_ (.A(_00491_),
    .B(net256),
    .Y(_03920_));
 sky130_fd_sc_hd__o22a_1 _11011_ (.A1(_06502_),
    .A2(net203),
    .B1(net231),
    .B2(reg1_val[10]),
    .X(_03921_));
 sky130_fd_sc_hd__o221a_1 _11012_ (.A1(_06505_),
    .A2(net194),
    .B1(_02440_),
    .B2(_06504_),
    .C1(_03921_),
    .X(_03922_));
 sky130_fd_sc_hd__o211a_1 _11013_ (.A1(_06506_),
    .A2(_02429_),
    .B1(_03920_),
    .C1(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__nand3_1 _11014_ (.A(_03916_),
    .B(_03919_),
    .C(_03923_),
    .Y(_03924_));
 sky130_fd_sc_hd__o21a_1 _11015_ (.A1(net222),
    .A2(_03234_),
    .B1(_02456_),
    .X(_03925_));
 sky130_fd_sc_hd__a221o_1 _11016_ (.A1(net167),
    .A2(_03911_),
    .B1(_03925_),
    .B2(net171),
    .C1(_03924_),
    .X(_03926_));
 sky130_fd_sc_hd__a211o_1 _11017_ (.A1(_03902_),
    .A2(_03903_),
    .B1(_03913_),
    .C1(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__a221o_1 _11018_ (.A1(_03895_),
    .A2(_03896_),
    .B1(_03898_),
    .B2(net233),
    .C1(_03927_),
    .X(_03928_));
 sky130_fd_sc_hd__a21o_1 _11019_ (.A1(curr_PC[9]),
    .A2(_03675_),
    .B1(curr_PC[10]),
    .X(_03929_));
 sky130_fd_sc_hd__and3_1 _11020_ (.A(curr_PC[9]),
    .B(curr_PC[10]),
    .C(_03675_),
    .X(_03930_));
 sky130_fd_sc_hd__nor2_1 _11021_ (.A(net237),
    .B(_03930_),
    .Y(_03931_));
 sky130_fd_sc_hd__a22o_4 _11022_ (.A1(net237),
    .A2(_03928_),
    .B1(_03929_),
    .B2(_03931_),
    .X(dest_val[10]));
 sky130_fd_sc_hd__o21ai_1 _11023_ (.A1(_03810_),
    .A2(_03894_),
    .B1(net136),
    .Y(_03932_));
 sky130_fd_sc_hd__a21bo_1 _11024_ (.A1(_03871_),
    .A2(_03877_),
    .B1_N(_03879_),
    .X(_03933_));
 sky130_fd_sc_hd__a21o_1 _11025_ (.A1(_03829_),
    .A2(_03835_),
    .B1(_03834_),
    .X(_03934_));
 sky130_fd_sc_hd__nand2_1 _11026_ (.A(_03845_),
    .B(_03934_),
    .Y(_03935_));
 sky130_fd_sc_hd__xor2_1 _11027_ (.A(_03845_),
    .B(_03934_),
    .X(_03936_));
 sky130_fd_sc_hd__o21ai_1 _11028_ (.A1(_03859_),
    .A2(_03861_),
    .B1(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__or3_1 _11029_ (.A(_03859_),
    .B(_03861_),
    .C(_03936_),
    .X(_03938_));
 sky130_fd_sc_hd__and2_1 _11030_ (.A(_03937_),
    .B(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__a22o_1 _11031_ (.A1(net101),
    .A2(net14),
    .B1(net31),
    .B2(_00203_),
    .X(_03940_));
 sky130_fd_sc_hd__xnor2_1 _11032_ (.A(net92),
    .B(_03940_),
    .Y(_03941_));
 sky130_fd_sc_hd__o22a_1 _11033_ (.A1(net41),
    .A2(net38),
    .B1(net36),
    .B2(net57),
    .X(_03942_));
 sky130_fd_sc_hd__xnor2_1 _11034_ (.A(net98),
    .B(_03942_),
    .Y(_03943_));
 sky130_fd_sc_hd__o22a_1 _11035_ (.A1(_00219_),
    .A2(net32),
    .B1(net70),
    .B2(net34),
    .X(_03944_));
 sky130_fd_sc_hd__xnor2_1 _11036_ (.A(net94),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__nand2_1 _11037_ (.A(_03943_),
    .B(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__or2_1 _11038_ (.A(_03943_),
    .B(_03945_),
    .X(_03947_));
 sky130_fd_sc_hd__nand2_1 _11039_ (.A(_03946_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__or2_1 _11040_ (.A(_03941_),
    .B(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__nand2_1 _11041_ (.A(_03941_),
    .B(_03948_),
    .Y(_03950_));
 sky130_fd_sc_hd__nand2_1 _11042_ (.A(_03949_),
    .B(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__a22o_1 _11043_ (.A1(_00443_),
    .A2(net9),
    .B1(net4),
    .B2(_00397_),
    .X(_03952_));
 sky130_fd_sc_hd__xnor2_1 _11044_ (.A(net62),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__o2bb2a_1 _11045_ (.A1_N(net73),
    .A2_N(net16),
    .B1(_00797_),
    .B2(net77),
    .X(_03954_));
 sky130_fd_sc_hd__xnor2_1 _11046_ (.A(_00787_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__nor2_1 _11047_ (.A(net115),
    .B(net59),
    .Y(_03956_));
 sky130_fd_sc_hd__xnor2_1 _11048_ (.A(_03955_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__nor2_1 _11049_ (.A(_03953_),
    .B(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__and2_1 _11050_ (.A(_03953_),
    .B(_03957_),
    .X(_03959_));
 sky130_fd_sc_hd__or2_1 _11051_ (.A(_03958_),
    .B(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__o22a_1 _11052_ (.A1(net45),
    .A2(net29),
    .B1(net27),
    .B2(net49),
    .X(_03961_));
 sky130_fd_sc_hd__xor2_1 _11053_ (.A(net89),
    .B(_03961_),
    .X(_03962_));
 sky130_fd_sc_hd__o22a_1 _11054_ (.A1(net53),
    .A2(net20),
    .B1(net18),
    .B2(net47),
    .X(_03963_));
 sky130_fd_sc_hd__xnor2_1 _11055_ (.A(net97),
    .B(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__o22a_1 _11056_ (.A1(net51),
    .A2(net25),
    .B1(net23),
    .B2(net43),
    .X(_03965_));
 sky130_fd_sc_hd__xnor2_1 _11057_ (.A(net87),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__and2_1 _11058_ (.A(_03964_),
    .B(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__xnor2_1 _11059_ (.A(_03964_),
    .B(_03966_),
    .Y(_03968_));
 sky130_fd_sc_hd__nor2_1 _11060_ (.A(_03962_),
    .B(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__and2_1 _11061_ (.A(_03962_),
    .B(_03968_),
    .X(_03970_));
 sky130_fd_sc_hd__or2_1 _11062_ (.A(_03969_),
    .B(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__nor2_1 _11063_ (.A(_03960_),
    .B(_03971_),
    .Y(_03972_));
 sky130_fd_sc_hd__and2_1 _11064_ (.A(_03960_),
    .B(_03971_),
    .X(_03973_));
 sky130_fd_sc_hd__nor2_1 _11065_ (.A(_03972_),
    .B(_03973_),
    .Y(_03974_));
 sky130_fd_sc_hd__xnor2_1 _11066_ (.A(_03951_),
    .B(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__nand2_1 _11067_ (.A(_03939_),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__or2_1 _11068_ (.A(_03939_),
    .B(_03975_),
    .X(_03977_));
 sky130_fd_sc_hd__nand2_1 _11069_ (.A(_03976_),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__a21oi_1 _11070_ (.A1(_03821_),
    .A2(_03823_),
    .B1(_03826_),
    .Y(_03979_));
 sky130_fd_sc_hd__o22a_1 _11071_ (.A1(_00460_),
    .A2(net10),
    .B1(net5),
    .B2(_00466_),
    .X(_03980_));
 sky130_fd_sc_hd__xnor2_1 _11072_ (.A(net109),
    .B(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__o22a_1 _11073_ (.A1(net84),
    .A2(_00517_),
    .B1(_00811_),
    .B2(net80),
    .X(_03982_));
 sky130_fd_sc_hd__xnor2_1 _11074_ (.A(net117),
    .B(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__nand2b_1 _11075_ (.A_N(net145),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__xnor2_1 _11076_ (.A(net145),
    .B(_03983_),
    .Y(_03985_));
 sky130_fd_sc_hd__nand2_1 _11077_ (.A(_03981_),
    .B(_03985_),
    .Y(_03986_));
 sky130_fd_sc_hd__or2_1 _11078_ (.A(_03981_),
    .B(_03985_),
    .X(_03987_));
 sky130_fd_sc_hd__nand2_1 _11079_ (.A(_03986_),
    .B(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__o21a_1 _11080_ (.A1(_03813_),
    .A2(_03819_),
    .B1(_03818_),
    .X(_03989_));
 sky130_fd_sc_hd__or2_1 _11081_ (.A(_03988_),
    .B(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__nand2_1 _11082_ (.A(_03988_),
    .B(_03989_),
    .Y(_03991_));
 sky130_fd_sc_hd__nand2_1 _11083_ (.A(_03990_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__xnor2_1 _11084_ (.A(_03979_),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__xor2_1 _11085_ (.A(_03978_),
    .B(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__o21a_1 _11086_ (.A1(_03851_),
    .A2(_03868_),
    .B1(_03850_),
    .X(_03995_));
 sky130_fd_sc_hd__nand2_1 _11087_ (.A(_03865_),
    .B(_03867_),
    .Y(_03996_));
 sky130_fd_sc_hd__o21bai_1 _11088_ (.A1(_03820_),
    .A2(_03839_),
    .B1_N(_03838_),
    .Y(_03997_));
 sky130_fd_sc_hd__a21oi_1 _11089_ (.A1(_03843_),
    .A2(_03848_),
    .B1(_03846_),
    .Y(_03998_));
 sky130_fd_sc_hd__o21ba_1 _11090_ (.A1(_03838_),
    .A2(_03840_),
    .B1_N(_03998_),
    .X(_03999_));
 sky130_fd_sc_hd__xnor2_1 _11091_ (.A(_03997_),
    .B(_03998_),
    .Y(_04000_));
 sky130_fd_sc_hd__xnor2_1 _11092_ (.A(_03996_),
    .B(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__a21bo_1 _11093_ (.A1(_03872_),
    .A2(_03876_),
    .B1_N(_03875_),
    .X(_04002_));
 sky130_fd_sc_hd__nand2b_1 _11094_ (.A_N(_04001_),
    .B(_04002_),
    .Y(_04003_));
 sky130_fd_sc_hd__xnor2_1 _11095_ (.A(_04001_),
    .B(_04002_),
    .Y(_04004_));
 sky130_fd_sc_hd__nand2b_1 _11096_ (.A_N(_03995_),
    .B(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__xnor2_1 _11097_ (.A(_03995_),
    .B(_04004_),
    .Y(_04006_));
 sky130_fd_sc_hd__nand2_1 _11098_ (.A(_03994_),
    .B(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__xnor2_1 _11099_ (.A(_03994_),
    .B(_04006_),
    .Y(_04008_));
 sky130_fd_sc_hd__nand2b_1 _11100_ (.A_N(_04008_),
    .B(_03933_),
    .Y(_04009_));
 sky130_fd_sc_hd__xor2_1 _11101_ (.A(_03933_),
    .B(_04008_),
    .X(_04010_));
 sky130_fd_sc_hd__a21oi_1 _11102_ (.A1(_03881_),
    .A2(_03883_),
    .B1(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__a21o_1 _11103_ (.A1(_03881_),
    .A2(_03883_),
    .B1(_04010_),
    .X(_04012_));
 sky130_fd_sc_hd__and3_1 _11104_ (.A(_03881_),
    .B(_03883_),
    .C(_04010_),
    .X(_04013_));
 sky130_fd_sc_hd__or2_2 _11105_ (.A(_04011_),
    .B(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__nor2_1 _11106_ (.A(_03764_),
    .B(_03887_),
    .Y(_04015_));
 sky130_fd_sc_hd__nand2_1 _11107_ (.A(_03766_),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__a31o_1 _11108_ (.A1(_03491_),
    .A2(_03492_),
    .A3(_03494_),
    .B1(_04016_),
    .X(_04017_));
 sky130_fd_sc_hd__a21boi_2 _11109_ (.A1(_03762_),
    .A2(_03885_),
    .B1_N(_03886_),
    .Y(_04018_));
 sky130_fd_sc_hd__a21o_1 _11110_ (.A1(_03765_),
    .A2(_04015_),
    .B1(_04018_),
    .X(_04019_));
 sky130_fd_sc_hd__inv_2 _11111_ (.A(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__a21oi_1 _11112_ (.A1(_04017_),
    .A2(_04020_),
    .B1(_04014_),
    .Y(_04021_));
 sky130_fd_sc_hd__and3_1 _11113_ (.A(_04014_),
    .B(_04017_),
    .C(_04020_),
    .X(_04022_));
 sky130_fd_sc_hd__or2_2 _11114_ (.A(_04021_),
    .B(_04022_),
    .X(_04023_));
 sky130_fd_sc_hd__or2_1 _11115_ (.A(_03932_),
    .B(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__a21oi_1 _11116_ (.A1(_03932_),
    .A2(_04023_),
    .B1(net235),
    .Y(_04025_));
 sky130_fd_sc_hd__nor2_1 _11117_ (.A(net134),
    .B(_01946_),
    .Y(_04026_));
 sky130_fd_sc_hd__xnor2_1 _11118_ (.A(_01948_),
    .B(_04026_),
    .Y(_04027_));
 sky130_fd_sc_hd__o21a_1 _11119_ (.A1(_06506_),
    .A2(_03899_),
    .B1(_06505_),
    .X(_04028_));
 sky130_fd_sc_hd__nor2_1 _11120_ (.A(net293),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__a31o_1 _11121_ (.A1(net293),
    .A2(_06503_),
    .A3(_06588_),
    .B1(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__nand2_1 _11122_ (.A(_06478_),
    .B(_04030_),
    .Y(_04031_));
 sky130_fd_sc_hd__o211a_1 _11123_ (.A1(_06478_),
    .A2(_04030_),
    .B1(_04031_),
    .C1(net234),
    .X(_04032_));
 sky130_fd_sc_hd__or2_1 _11124_ (.A(net290),
    .B(curr_PC[11]),
    .X(_04033_));
 sky130_fd_sc_hd__and2_1 _11125_ (.A(net290),
    .B(curr_PC[11]),
    .X(_04034_));
 sky130_fd_sc_hd__nand2_1 _11126_ (.A(net290),
    .B(curr_PC[11]),
    .Y(_04035_));
 sky130_fd_sc_hd__a211o_1 _11127_ (.A1(_04033_),
    .A2(_04035_),
    .B1(_03905_),
    .C1(_03909_),
    .X(_04036_));
 sky130_fd_sc_hd__o211a_1 _11128_ (.A1(_03905_),
    .A2(_03909_),
    .B1(_04033_),
    .C1(_04035_),
    .X(_04037_));
 sky130_fd_sc_hd__nor2_1 _11129_ (.A(net223),
    .B(_04037_),
    .Y(_04038_));
 sky130_fd_sc_hd__mux2_1 _11130_ (.A0(_02919_),
    .A1(_02923_),
    .S(net218),
    .X(_04039_));
 sky130_fd_sc_hd__mux2_2 _11131_ (.A0(_03108_),
    .A1(_04039_),
    .S(net220),
    .X(_04040_));
 sky130_fd_sc_hd__a22o_1 _11132_ (.A1(_04036_),
    .A2(_04038_),
    .B1(_04040_),
    .B2(net223),
    .X(_04041_));
 sky130_fd_sc_hd__or2_1 _11133_ (.A(\div_res[10] ),
    .B(_03914_),
    .X(_04042_));
 sky130_fd_sc_hd__a21oi_1 _11134_ (.A1(net139),
    .A2(_04042_),
    .B1(\div_res[11] ),
    .Y(_04043_));
 sky130_fd_sc_hd__a31o_1 _11135_ (.A1(\div_res[11] ),
    .A2(net139),
    .A3(_04042_),
    .B1(net189),
    .X(_04044_));
 sky130_fd_sc_hd__o21a_1 _11136_ (.A1(\div_shifter[42] ),
    .A2(_03917_),
    .B1(net228),
    .X(_04045_));
 sky130_fd_sc_hd__xnor2_2 _11137_ (.A(\div_shifter[43] ),
    .B(_04045_),
    .Y(_04046_));
 sky130_fd_sc_hd__nand2_1 _11138_ (.A(_06452_),
    .B(net193),
    .Y(_04047_));
 sky130_fd_sc_hd__o221a_1 _11139_ (.A1(_06435_),
    .A2(net203),
    .B1(net231),
    .B2(net290),
    .C1(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__o221a_1 _11140_ (.A1(_06469_),
    .A2(_02429_),
    .B1(net194),
    .B2(_06461_),
    .C1(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__o221a_1 _11141_ (.A1(_00451_),
    .A2(_02432_),
    .B1(net192),
    .B2(_04046_),
    .C1(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__o21ai_1 _11142_ (.A1(_04043_),
    .A2(_04044_),
    .B1(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__o21a_1 _11143_ (.A1(net221),
    .A2(_03095_),
    .B1(_02456_),
    .X(_04052_));
 sky130_fd_sc_hd__a221o_1 _11144_ (.A1(net167),
    .A2(_04040_),
    .B1(_04052_),
    .B2(net171),
    .C1(_04051_),
    .X(_04053_));
 sky130_fd_sc_hd__a211o_1 _11145_ (.A1(net205),
    .A2(_04041_),
    .B1(_04053_),
    .C1(_04032_),
    .X(_04054_));
 sky130_fd_sc_hd__a221o_1 _11146_ (.A1(_04024_),
    .A2(_04025_),
    .B1(_04027_),
    .B2(net233),
    .C1(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__and2_1 _11147_ (.A(curr_PC[11]),
    .B(_03930_),
    .X(_04056_));
 sky130_fd_sc_hd__o21ai_1 _11148_ (.A1(curr_PC[11]),
    .A2(_03930_),
    .B1(net242),
    .Y(_04057_));
 sky130_fd_sc_hd__a2bb2o_4 _11149_ (.A1_N(_04056_),
    .A2_N(_04057_),
    .B1(net237),
    .B2(_04055_),
    .X(dest_val[11]));
 sky130_fd_sc_hd__o21ba_1 _11150_ (.A1(_04021_),
    .A2(_04022_),
    .B1_N(_03894_),
    .X(_04058_));
 sky130_fd_sc_hd__or4bb_4 _11151_ (.A(_03636_),
    .B(_03639_),
    .C_N(_03771_),
    .D_N(_04058_),
    .X(_04059_));
 sky130_fd_sc_hd__nand2_2 _11152_ (.A(_04007_),
    .B(_04009_),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_1 _11153_ (.A(_04003_),
    .B(_04005_),
    .Y(_04061_));
 sky130_fd_sc_hd__a31o_1 _11154_ (.A1(_00392_),
    .A2(net62),
    .A3(_03955_),
    .B1(_03958_),
    .X(_04062_));
 sky130_fd_sc_hd__o22a_1 _11155_ (.A1(net84),
    .A2(_00811_),
    .B1(net10),
    .B2(_00444_),
    .X(_04063_));
 sky130_fd_sc_hd__xnor2_2 _11156_ (.A(net117),
    .B(_04063_),
    .Y(_04064_));
 sky130_fd_sc_hd__nand2_1 _11157_ (.A(_00459_),
    .B(net6),
    .Y(_04065_));
 sky130_fd_sc_hd__a22o_2 _11158_ (.A1(_00458_),
    .A2(net6),
    .B1(_04065_),
    .B2(net108),
    .X(_04066_));
 sky130_fd_sc_hd__xor2_1 _11159_ (.A(_04064_),
    .B(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__a21oi_1 _11160_ (.A1(_03946_),
    .A2(_03949_),
    .B1(_04067_),
    .Y(_04068_));
 sky130_fd_sc_hd__and3_1 _11161_ (.A(_03946_),
    .B(_03949_),
    .C(_04067_),
    .X(_04069_));
 sky130_fd_sc_hd__nor2_1 _11162_ (.A(_04068_),
    .B(_04069_),
    .Y(_04070_));
 sky130_fd_sc_hd__xnor2_1 _11163_ (.A(_04062_),
    .B(_04070_),
    .Y(_04071_));
 sky130_fd_sc_hd__a22o_1 _11164_ (.A1(_00203_),
    .A2(net14),
    .B1(net30),
    .B2(_00208_),
    .X(_04072_));
 sky130_fd_sc_hd__xnor2_1 _11165_ (.A(net91),
    .B(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__o22a_1 _11166_ (.A1(net103),
    .A2(net34),
    .B1(net32),
    .B2(_00230_),
    .X(_04074_));
 sky130_fd_sc_hd__xnor2_1 _11167_ (.A(net93),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__o22a_1 _11168_ (.A1(net57),
    .A2(net38),
    .B1(net36),
    .B2(net54),
    .X(_04076_));
 sky130_fd_sc_hd__xnor2_1 _11169_ (.A(net98),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__and2_1 _11170_ (.A(_04075_),
    .B(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__nor2_1 _11171_ (.A(_04075_),
    .B(_04077_),
    .Y(_04079_));
 sky130_fd_sc_hd__or2_1 _11172_ (.A(_04078_),
    .B(_04079_),
    .X(_04080_));
 sky130_fd_sc_hd__inv_2 _11173_ (.A(_04080_),
    .Y(_04081_));
 sky130_fd_sc_hd__xor2_1 _11174_ (.A(_04073_),
    .B(_04080_),
    .X(_04082_));
 sky130_fd_sc_hd__o22a_1 _11175_ (.A1(net50),
    .A2(net29),
    .B1(net27),
    .B2(net51),
    .X(_04083_));
 sky130_fd_sc_hd__xnor2_1 _11176_ (.A(net89),
    .B(_04083_),
    .Y(_04084_));
 sky130_fd_sc_hd__o32a_1 _11177_ (.A1(net23),
    .A2(_00513_),
    .A3(_00515_),
    .B1(net25),
    .B2(net43),
    .X(_04085_));
 sky130_fd_sc_hd__xnor2_2 _11178_ (.A(net87),
    .B(_04085_),
    .Y(_04086_));
 sky130_fd_sc_hd__o22a_1 _11179_ (.A1(net47),
    .A2(net20),
    .B1(net18),
    .B2(net46),
    .X(_04087_));
 sky130_fd_sc_hd__xnor2_2 _11180_ (.A(net97),
    .B(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__nand2_1 _11181_ (.A(_04086_),
    .B(_04088_),
    .Y(_04089_));
 sky130_fd_sc_hd__xnor2_2 _11182_ (.A(_04086_),
    .B(_04088_),
    .Y(_04090_));
 sky130_fd_sc_hd__inv_2 _11183_ (.A(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__nand2_1 _11184_ (.A(_04084_),
    .B(_04091_),
    .Y(_04092_));
 sky130_fd_sc_hd__xor2_1 _11185_ (.A(_04084_),
    .B(_04090_),
    .X(_04093_));
 sky130_fd_sc_hd__a22o_1 _11186_ (.A1(net71),
    .A2(net17),
    .B1(net12),
    .B2(net73),
    .X(_04094_));
 sky130_fd_sc_hd__xnor2_1 _11187_ (.A(net65),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__a22o_1 _11188_ (.A1(_00446_),
    .A2(net9),
    .B1(net4),
    .B2(_00443_),
    .X(_04096_));
 sky130_fd_sc_hd__xnor2_1 _11189_ (.A(net59),
    .B(_04096_),
    .Y(_04097_));
 sky130_fd_sc_hd__nand2_1 _11190_ (.A(_04095_),
    .B(_04097_),
    .Y(_04098_));
 sky130_fd_sc_hd__xnor2_1 _11191_ (.A(_04095_),
    .B(_04097_),
    .Y(_04099_));
 sky130_fd_sc_hd__nor2_1 _11192_ (.A(_04093_),
    .B(_04099_),
    .Y(_04100_));
 sky130_fd_sc_hd__xor2_1 _11193_ (.A(_04093_),
    .B(_04099_),
    .X(_04101_));
 sky130_fd_sc_hd__and2b_1 _11194_ (.A_N(_04082_),
    .B(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__xnor2_1 _11195_ (.A(_04082_),
    .B(_04101_),
    .Y(_04103_));
 sky130_fd_sc_hd__o211a_1 _11196_ (.A1(_03967_),
    .A2(_03969_),
    .B1(_00397_),
    .C1(net62),
    .X(_04104_));
 sky130_fd_sc_hd__a211oi_2 _11197_ (.A1(_00397_),
    .A2(net62),
    .B1(_03967_),
    .C1(_03969_),
    .Y(_04105_));
 sky130_fd_sc_hd__a211oi_2 _11198_ (.A1(_03984_),
    .A2(_03986_),
    .B1(_04104_),
    .C1(_04105_),
    .Y(_04106_));
 sky130_fd_sc_hd__o211a_1 _11199_ (.A1(_04104_),
    .A2(_04105_),
    .B1(_03984_),
    .C1(_03986_),
    .X(_04107_));
 sky130_fd_sc_hd__nor2_1 _11200_ (.A(_04106_),
    .B(_04107_),
    .Y(_04108_));
 sky130_fd_sc_hd__nand2_1 _11201_ (.A(_04103_),
    .B(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__or2_1 _11202_ (.A(_04103_),
    .B(_04108_),
    .X(_04110_));
 sky130_fd_sc_hd__nand2_1 _11203_ (.A(_04109_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__xor2_1 _11204_ (.A(_04071_),
    .B(_04111_),
    .X(_04112_));
 sky130_fd_sc_hd__o21ai_1 _11205_ (.A1(_03978_),
    .A2(_03993_),
    .B1(_03976_),
    .Y(_04113_));
 sky130_fd_sc_hd__o21ai_1 _11206_ (.A1(_03979_),
    .A2(_03992_),
    .B1(_03990_),
    .Y(_04114_));
 sky130_fd_sc_hd__o21ba_1 _11207_ (.A1(_03951_),
    .A2(_03973_),
    .B1_N(_03972_),
    .X(_04115_));
 sky130_fd_sc_hd__a21oi_1 _11208_ (.A1(_03935_),
    .A2(_03937_),
    .B1(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__and3_1 _11209_ (.A(_03935_),
    .B(_03937_),
    .C(_04115_),
    .X(_04117_));
 sky130_fd_sc_hd__nor2_1 _11210_ (.A(_04116_),
    .B(_04117_),
    .Y(_04118_));
 sky130_fd_sc_hd__xnor2_1 _11211_ (.A(_04114_),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__a21oi_1 _11212_ (.A1(_03996_),
    .A2(_04000_),
    .B1(_03999_),
    .Y(_04120_));
 sky130_fd_sc_hd__xnor2_1 _11213_ (.A(_04119_),
    .B(_04120_),
    .Y(_04121_));
 sky130_fd_sc_hd__nand2b_1 _11214_ (.A_N(_04121_),
    .B(_04113_),
    .Y(_04122_));
 sky130_fd_sc_hd__xnor2_1 _11215_ (.A(_04113_),
    .B(_04121_),
    .Y(_04123_));
 sky130_fd_sc_hd__nand2_1 _11216_ (.A(_04112_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__xor2_1 _11217_ (.A(_04112_),
    .B(_04123_),
    .X(_04125_));
 sky130_fd_sc_hd__nand2_1 _11218_ (.A(_04061_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__or2_1 _11219_ (.A(_04061_),
    .B(_04125_),
    .X(_04127_));
 sky130_fd_sc_hd__nand2_2 _11220_ (.A(_04126_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__a21o_1 _11221_ (.A1(_04007_),
    .A2(_04009_),
    .B1(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__and3_1 _11222_ (.A(_04007_),
    .B(_04009_),
    .C(_04128_),
    .X(_04130_));
 sky130_fd_sc_hd__xor2_4 _11223_ (.A(_04060_),
    .B(_04128_),
    .X(_04131_));
 sky130_fd_sc_hd__a21oi_2 _11224_ (.A1(_03885_),
    .A2(_04012_),
    .B1(_04013_),
    .Y(_04132_));
 sky130_fd_sc_hd__nor2_1 _11225_ (.A(_03887_),
    .B(_04014_),
    .Y(_04133_));
 sky130_fd_sc_hd__a21o_1 _11226_ (.A1(_03888_),
    .A2(_04133_),
    .B1(_04132_),
    .X(_04134_));
 sky130_fd_sc_hd__nand2_1 _11227_ (.A(_03889_),
    .B(_04133_),
    .Y(_04135_));
 sky130_fd_sc_hd__o21ba_1 _11228_ (.A1(_03545_),
    .A2(_04135_),
    .B1_N(_04134_),
    .X(_04136_));
 sky130_fd_sc_hd__xor2_4 _11229_ (.A(_04131_),
    .B(_04136_),
    .X(_04137_));
 sky130_fd_sc_hd__a21o_1 _11230_ (.A1(net136),
    .A2(_04059_),
    .B1(_04137_),
    .X(_04138_));
 sky130_fd_sc_hd__nand3_1 _11231_ (.A(net144),
    .B(_04059_),
    .C(_04137_),
    .Y(_04139_));
 sky130_fd_sc_hd__a21o_1 _11232_ (.A1(_01946_),
    .A2(_01948_),
    .B1(net134),
    .X(_04140_));
 sky130_fd_sc_hd__xnor2_1 _11233_ (.A(_01951_),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__o21a_1 _11234_ (.A1(_06469_),
    .A2(_04028_),
    .B1(_06461_),
    .X(_04142_));
 sky130_fd_sc_hd__nor2_1 _11235_ (.A(net293),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__a31o_1 _11236_ (.A1(net293),
    .A2(_06443_),
    .A3(_06589_),
    .B1(_04143_),
    .X(_04144_));
 sky130_fd_sc_hd__nand2_1 _11237_ (.A(_06399_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__o211a_1 _11238_ (.A1(_06399_),
    .A2(_04144_),
    .B1(_04145_),
    .C1(net234),
    .X(_04146_));
 sky130_fd_sc_hd__mux2_1 _11239_ (.A0(_03089_),
    .A1(_03093_),
    .S(net218),
    .X(_04147_));
 sky130_fd_sc_hd__inv_2 _11240_ (.A(_04147_),
    .Y(_04148_));
 sky130_fd_sc_hd__mux2_1 _11241_ (.A0(_02937_),
    .A1(_04148_),
    .S(net220),
    .X(_04149_));
 sky130_fd_sc_hd__or2_1 _11242_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .X(_04150_));
 sky130_fd_sc_hd__nand2_1 _11243_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .Y(_04151_));
 sky130_fd_sc_hd__o211a_1 _11244_ (.A1(_04034_),
    .A2(_04037_),
    .B1(_04150_),
    .C1(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__a211o_1 _11245_ (.A1(_04150_),
    .A2(_04151_),
    .B1(_04034_),
    .C1(_04037_),
    .X(_04153_));
 sky130_fd_sc_hd__nand2_1 _11246_ (.A(net244),
    .B(_04153_),
    .Y(_04154_));
 sky130_fd_sc_hd__a2bb2o_1 _11247_ (.A1_N(_04152_),
    .A2_N(_04154_),
    .B1(net223),
    .B2(_04149_),
    .X(_04155_));
 sky130_fd_sc_hd__or3_1 _11248_ (.A(\div_res[11] ),
    .B(\div_res[10] ),
    .C(_03914_),
    .X(_04156_));
 sky130_fd_sc_hd__a21o_1 _11249_ (.A1(net139),
    .A2(_04156_),
    .B1(\div_res[12] ),
    .X(_04157_));
 sky130_fd_sc_hd__a31oi_1 _11250_ (.A1(\div_res[12] ),
    .A2(net139),
    .A3(_04156_),
    .B1(net189),
    .Y(_04158_));
 sky130_fd_sc_hd__or3_1 _11251_ (.A(\div_shifter[43] ),
    .B(\div_shifter[42] ),
    .C(_03917_),
    .X(_04159_));
 sky130_fd_sc_hd__nand3_1 _11252_ (.A(\div_shifter[44] ),
    .B(net228),
    .C(_04159_),
    .Y(_04160_));
 sky130_fd_sc_hd__a21o_1 _11253_ (.A1(net228),
    .A2(_04159_),
    .B1(\div_shifter[44] ),
    .X(_04161_));
 sky130_fd_sc_hd__o22a_1 _11254_ (.A1(_06363_),
    .A2(net203),
    .B1(net231),
    .B2(reg1_val[12]),
    .X(_04162_));
 sky130_fd_sc_hd__o21ai_1 _11255_ (.A1(_06390_),
    .A2(net194),
    .B1(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__a221o_1 _11256_ (.A1(_06399_),
    .A2(net195),
    .B1(net193),
    .B2(_06381_),
    .C1(_04163_),
    .X(_04164_));
 sky130_fd_sc_hd__a31o_2 _11257_ (.A1(_00241_),
    .A2(_00453_),
    .A3(net256),
    .B1(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__a31o_1 _11258_ (.A1(_02441_),
    .A2(_04160_),
    .A3(_04161_),
    .B1(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__o21a_1 _11259_ (.A1(net222),
    .A2(_02926_),
    .B1(_02456_),
    .X(_04167_));
 sky130_fd_sc_hd__a221o_1 _11260_ (.A1(_04157_),
    .A2(_04158_),
    .B1(_04167_),
    .B2(net171),
    .C1(_04166_),
    .X(_04168_));
 sky130_fd_sc_hd__a221o_1 _11261_ (.A1(net167),
    .A2(_04149_),
    .B1(_04155_),
    .B2(net205),
    .C1(_04168_),
    .X(_04169_));
 sky130_fd_sc_hd__a211o_1 _11262_ (.A1(net233),
    .A2(_04141_),
    .B1(_04146_),
    .C1(_04169_),
    .X(_04170_));
 sky130_fd_sc_hd__a31o_1 _11263_ (.A1(_02348_),
    .A2(_04138_),
    .A3(_04139_),
    .B1(_04170_),
    .X(_04171_));
 sky130_fd_sc_hd__or2_1 _11264_ (.A(curr_PC[12]),
    .B(_04056_),
    .X(_04172_));
 sky130_fd_sc_hd__and3_1 _11265_ (.A(curr_PC[11]),
    .B(curr_PC[12]),
    .C(_03930_),
    .X(_04173_));
 sky130_fd_sc_hd__nor2_1 _11266_ (.A(net238),
    .B(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__a22o_4 _11267_ (.A1(net238),
    .A2(_04171_),
    .B1(_04172_),
    .B2(_04174_),
    .X(dest_val[12]));
 sky130_fd_sc_hd__or2_1 _11268_ (.A(_04059_),
    .B(_04137_),
    .X(_04175_));
 sky130_fd_sc_hd__o2bb2a_1 _11269_ (.A1_N(net102),
    .A2_N(net16),
    .B1(_00797_),
    .B2(_00468_),
    .X(_04176_));
 sky130_fd_sc_hd__xnor2_1 _11270_ (.A(_00787_),
    .B(_04176_),
    .Y(_04177_));
 sky130_fd_sc_hd__o22a_1 _11271_ (.A1(net41),
    .A2(_00336_),
    .B1(_00342_),
    .B2(net57),
    .X(_04178_));
 sky130_fd_sc_hd__xnor2_1 _11272_ (.A(_00308_),
    .B(_04178_),
    .Y(_04179_));
 sky130_fd_sc_hd__nand2_1 _11273_ (.A(_04177_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__or2_1 _11274_ (.A(_04177_),
    .B(_04179_),
    .X(_04181_));
 sky130_fd_sc_hd__nand2_1 _11275_ (.A(_04180_),
    .B(_04181_),
    .Y(_04182_));
 sky130_fd_sc_hd__o22a_1 _11276_ (.A1(_00230_),
    .A2(net34),
    .B1(net32),
    .B2(_00202_),
    .X(_04183_));
 sky130_fd_sc_hd__xnor2_1 _11277_ (.A(net93),
    .B(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__nand2b_1 _11278_ (.A_N(_04182_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__xor2_1 _11279_ (.A(_04182_),
    .B(_04184_),
    .X(_04186_));
 sky130_fd_sc_hd__o22a_1 _11280_ (.A1(net83),
    .A2(net10),
    .B1(net5),
    .B2(net80),
    .X(_04187_));
 sky130_fd_sc_hd__xnor2_1 _11281_ (.A(net117),
    .B(_04187_),
    .Y(_04188_));
 sky130_fd_sc_hd__nand2_1 _11282_ (.A(_00389_),
    .B(_00516_),
    .Y(_04189_));
 sky130_fd_sc_hd__nand2_1 _11283_ (.A(_00393_),
    .B(_00812_),
    .Y(_04190_));
 sky130_fd_sc_hd__a21o_1 _11284_ (.A1(_04189_),
    .A2(_04190_),
    .B1(_00359_),
    .X(_04191_));
 sky130_fd_sc_hd__nand3_1 _11285_ (.A(_00359_),
    .B(_04189_),
    .C(_04190_),
    .Y(_04192_));
 sky130_fd_sc_hd__nand3_1 _11286_ (.A(_00431_),
    .B(_04191_),
    .C(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__a21o_1 _11287_ (.A1(_04191_),
    .A2(_04192_),
    .B1(_00431_),
    .X(_04194_));
 sky130_fd_sc_hd__and3_1 _11288_ (.A(_04188_),
    .B(_04193_),
    .C(_04194_),
    .X(_04195_));
 sky130_fd_sc_hd__a21oi_1 _11289_ (.A1(_04193_),
    .A2(_04194_),
    .B1(_04188_),
    .Y(_04196_));
 sky130_fd_sc_hd__or3_1 _11290_ (.A(_04186_),
    .B(_04195_),
    .C(_04196_),
    .X(_04197_));
 sky130_fd_sc_hd__o21ai_2 _11291_ (.A1(_04195_),
    .A2(_04196_),
    .B1(_04186_),
    .Y(_04198_));
 sky130_fd_sc_hd__o22a_1 _11292_ (.A1(net46),
    .A2(net20),
    .B1(net18),
    .B2(net50),
    .X(_04199_));
 sky130_fd_sc_hd__xnor2_2 _11293_ (.A(_00274_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__o22a_1 _11294_ (.A1(net54),
    .A2(net38),
    .B1(_00288_),
    .B2(net48),
    .X(_04201_));
 sky130_fd_sc_hd__xnor2_1 _11295_ (.A(_00262_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__o22a_1 _11296_ (.A1(net52),
    .A2(net29),
    .B1(net27),
    .B2(net43),
    .X(_04203_));
 sky130_fd_sc_hd__xnor2_1 _11297_ (.A(net90),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__nand2_1 _11298_ (.A(_04202_),
    .B(_04204_),
    .Y(_04205_));
 sky130_fd_sc_hd__or2_1 _11299_ (.A(_04202_),
    .B(_04204_),
    .X(_04206_));
 sky130_fd_sc_hd__nand2_1 _11300_ (.A(_04205_),
    .B(_04206_),
    .Y(_04207_));
 sky130_fd_sc_hd__xor2_2 _11301_ (.A(_04200_),
    .B(_04207_),
    .X(_04208_));
 sky130_fd_sc_hd__and3_1 _11302_ (.A(_04197_),
    .B(_04198_),
    .C(_04208_),
    .X(_04209_));
 sky130_fd_sc_hd__a21oi_1 _11303_ (.A1(_04197_),
    .A2(_04198_),
    .B1(_04208_),
    .Y(_04210_));
 sky130_fd_sc_hd__a22o_1 _11304_ (.A1(net73),
    .A2(net9),
    .B1(net4),
    .B2(_00446_),
    .X(_04211_));
 sky130_fd_sc_hd__xnor2_1 _11305_ (.A(net59),
    .B(_04211_),
    .Y(_04212_));
 sky130_fd_sc_hd__o21ai_1 _11306_ (.A1(_04064_),
    .A2(_04066_),
    .B1(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__or3_1 _11307_ (.A(_04064_),
    .B(_04066_),
    .C(_04212_),
    .X(_04214_));
 sky130_fd_sc_hd__nand2_1 _11308_ (.A(_04213_),
    .B(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__nand2_1 _11309_ (.A(_00443_),
    .B(net62),
    .Y(_04216_));
 sky130_fd_sc_hd__xnor2_1 _11310_ (.A(_04215_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__or3_1 _11311_ (.A(_04209_),
    .B(_04210_),
    .C(_04217_),
    .X(_04218_));
 sky130_fd_sc_hd__o21ai_1 _11312_ (.A1(_04209_),
    .A2(_04210_),
    .B1(_04217_),
    .Y(_04219_));
 sky130_fd_sc_hd__a21o_1 _11313_ (.A1(_04073_),
    .A2(_04081_),
    .B1(_04078_),
    .X(_04220_));
 sky130_fd_sc_hd__a21o_1 _11314_ (.A1(_04089_),
    .A2(_04092_),
    .B1(_04098_),
    .X(_04221_));
 sky130_fd_sc_hd__nand3_1 _11315_ (.A(_04089_),
    .B(_04092_),
    .C(_04098_),
    .Y(_04222_));
 sky130_fd_sc_hd__nand2_1 _11316_ (.A(_04221_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__nand2b_1 _11317_ (.A_N(_04223_),
    .B(_04220_),
    .Y(_04224_));
 sky130_fd_sc_hd__xnor2_1 _11318_ (.A(_04220_),
    .B(_04223_),
    .Y(_04225_));
 sky130_fd_sc_hd__and3_1 _11319_ (.A(_04218_),
    .B(_04219_),
    .C(_04225_),
    .X(_04226_));
 sky130_fd_sc_hd__a21oi_1 _11320_ (.A1(_04218_),
    .A2(_04219_),
    .B1(_04225_),
    .Y(_04227_));
 sky130_fd_sc_hd__nor2_1 _11321_ (.A(_04226_),
    .B(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__o21ai_1 _11322_ (.A1(_04071_),
    .A2(_04111_),
    .B1(_04109_),
    .Y(_04229_));
 sky130_fd_sc_hd__a21o_1 _11323_ (.A1(_04114_),
    .A2(_04118_),
    .B1(_04116_),
    .X(_04230_));
 sky130_fd_sc_hd__a21oi_1 _11324_ (.A1(_04062_),
    .A2(_04070_),
    .B1(_04068_),
    .Y(_04231_));
 sky130_fd_sc_hd__o22a_1 _11325_ (.A1(_04100_),
    .A2(_04102_),
    .B1(_04104_),
    .B2(_04106_),
    .X(_04232_));
 sky130_fd_sc_hd__or4_1 _11326_ (.A(_04100_),
    .B(_04102_),
    .C(_04104_),
    .D(_04106_),
    .X(_04233_));
 sky130_fd_sc_hd__and2b_1 _11327_ (.A_N(_04232_),
    .B(_04233_),
    .X(_04234_));
 sky130_fd_sc_hd__and2b_1 _11328_ (.A_N(_04231_),
    .B(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__xnor2_1 _11329_ (.A(_04231_),
    .B(_04234_),
    .Y(_04236_));
 sky130_fd_sc_hd__nand2_1 _11330_ (.A(_04230_),
    .B(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__xor2_1 _11331_ (.A(_04230_),
    .B(_04236_),
    .X(_04238_));
 sky130_fd_sc_hd__xor2_1 _11332_ (.A(_04229_),
    .B(_04238_),
    .X(_04239_));
 sky130_fd_sc_hd__nand2_1 _11333_ (.A(_04228_),
    .B(_04239_),
    .Y(_04240_));
 sky130_fd_sc_hd__xnor2_1 _11334_ (.A(_04228_),
    .B(_04239_),
    .Y(_04241_));
 sky130_fd_sc_hd__o21a_1 _11335_ (.A1(_04119_),
    .A2(_04120_),
    .B1(_04122_),
    .X(_04242_));
 sky130_fd_sc_hd__or2_1 _11336_ (.A(_04241_),
    .B(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__xnor2_1 _11337_ (.A(_04241_),
    .B(_04242_),
    .Y(_04244_));
 sky130_fd_sc_hd__a21oi_1 _11338_ (.A1(_04124_),
    .A2(_04126_),
    .B1(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__a21o_1 _11339_ (.A1(_04124_),
    .A2(_04126_),
    .B1(_04244_),
    .X(_04246_));
 sky130_fd_sc_hd__and3_1 _11340_ (.A(_04124_),
    .B(_04126_),
    .C(_04244_),
    .X(_04247_));
 sky130_fd_sc_hd__or2_4 _11341_ (.A(_04245_),
    .B(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__nor2_1 _11342_ (.A(_04014_),
    .B(_04131_),
    .Y(_04249_));
 sky130_fd_sc_hd__nand2_2 _11343_ (.A(_04015_),
    .B(_04249_),
    .Y(_04250_));
 sky130_fd_sc_hd__a21oi_2 _11344_ (.A1(_04012_),
    .A2(_04129_),
    .B1(_04130_),
    .Y(_04251_));
 sky130_fd_sc_hd__a21o_1 _11345_ (.A1(_04018_),
    .A2(_04249_),
    .B1(_04251_),
    .X(_04252_));
 sky130_fd_sc_hd__o21bai_4 _11346_ (.A1(_03770_),
    .A2(_04250_),
    .B1_N(_04252_),
    .Y(_04253_));
 sky130_fd_sc_hd__xnor2_4 _11347_ (.A(_04248_),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__nand3_1 _11348_ (.A(net136),
    .B(_04175_),
    .C(_04254_),
    .Y(_04255_));
 sky130_fd_sc_hd__a21o_1 _11349_ (.A1(net136),
    .A2(_04175_),
    .B1(_04254_),
    .X(_04256_));
 sky130_fd_sc_hd__a21oi_1 _11350_ (.A1(net136),
    .A2(_01952_),
    .B1(_01953_),
    .Y(_04257_));
 sky130_fd_sc_hd__a31o_1 _11351_ (.A1(net136),
    .A2(_01952_),
    .A3(_01953_),
    .B1(_02434_),
    .X(_04258_));
 sky130_fd_sc_hd__nor2_1 _11352_ (.A(_04257_),
    .B(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__o21a_1 _11353_ (.A1(_06408_),
    .A2(_04142_),
    .B1(_06390_),
    .X(_04260_));
 sky130_fd_sc_hd__nor2_1 _11354_ (.A(net294),
    .B(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__a31o_1 _11355_ (.A1(net293),
    .A2(_06372_),
    .A3(_06590_),
    .B1(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__nor2_1 _11356_ (.A(_06345_),
    .B(_04262_),
    .Y(_04263_));
 sky130_fd_sc_hd__a21o_1 _11357_ (.A1(_06345_),
    .A2(_04262_),
    .B1(_02427_),
    .X(_04264_));
 sky130_fd_sc_hd__or2_1 _11358_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .X(_04265_));
 sky130_fd_sc_hd__nand2_1 _11359_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .Y(_04266_));
 sky130_fd_sc_hd__nand2_1 _11360_ (.A(_04265_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__a21oi_1 _11361_ (.A1(reg1_val[12]),
    .A2(curr_PC[12]),
    .B1(_04152_),
    .Y(_04268_));
 sky130_fd_sc_hd__xor2_1 _11362_ (.A(_04267_),
    .B(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__mux2_1 _11363_ (.A0(_03231_),
    .A1(_03233_),
    .S(net219),
    .X(_04270_));
 sky130_fd_sc_hd__mux2_1 _11364_ (.A0(_02754_),
    .A1(_04270_),
    .S(net220),
    .X(_04271_));
 sky130_fd_sc_hd__mux2_1 _11365_ (.A0(_04269_),
    .A1(_04271_),
    .S(net224),
    .X(_04272_));
 sky130_fd_sc_hd__or2_1 _11366_ (.A(\div_res[12] ),
    .B(_04156_),
    .X(_04273_));
 sky130_fd_sc_hd__a21oi_1 _11367_ (.A1(net139),
    .A2(_04273_),
    .B1(\div_res[13] ),
    .Y(_04274_));
 sky130_fd_sc_hd__a31o_1 _11368_ (.A1(\div_res[13] ),
    .A2(net139),
    .A3(_04273_),
    .B1(net189),
    .X(_04275_));
 sky130_fd_sc_hd__or2_1 _11369_ (.A(\div_shifter[44] ),
    .B(_04159_),
    .X(_04276_));
 sky130_fd_sc_hd__a21oi_1 _11370_ (.A1(net228),
    .A2(_04276_),
    .B1(\div_shifter[45] ),
    .Y(_04277_));
 sky130_fd_sc_hd__a31o_1 _11371_ (.A1(\div_shifter[45] ),
    .A2(net227),
    .A3(_04276_),
    .B1(net191),
    .X(_04278_));
 sky130_fd_sc_hd__or3_2 _11372_ (.A(_00244_),
    .B(_00428_),
    .C(_02432_),
    .X(_04279_));
 sky130_fd_sc_hd__nand2_1 _11373_ (.A(_06327_),
    .B(net193),
    .Y(_04280_));
 sky130_fd_sc_hd__o221a_1 _11374_ (.A1(_06315_),
    .A2(net203),
    .B1(net231),
    .B2(reg1_val[13]),
    .C1(_04280_),
    .X(_04281_));
 sky130_fd_sc_hd__o221a_1 _11375_ (.A1(_06339_),
    .A2(_02429_),
    .B1(net194),
    .B2(_06333_),
    .C1(_04281_),
    .X(_04282_));
 sky130_fd_sc_hd__o211a_1 _11376_ (.A1(_04277_),
    .A2(_04278_),
    .B1(_04279_),
    .C1(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__o21ai_2 _11377_ (.A1(net221),
    .A2(_02770_),
    .B1(_02456_),
    .Y(_04284_));
 sky130_fd_sc_hd__o221ai_2 _11378_ (.A1(_04274_),
    .A2(_04275_),
    .B1(_04284_),
    .B2(net168),
    .C1(_04283_),
    .Y(_04285_));
 sky130_fd_sc_hd__a221o_1 _11379_ (.A1(net167),
    .A2(_04271_),
    .B1(_04272_),
    .B2(net205),
    .C1(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__o21bai_1 _11380_ (.A1(_04263_),
    .A2(_04264_),
    .B1_N(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__a311o_1 _11381_ (.A1(_02348_),
    .A2(_04255_),
    .A3(_04256_),
    .B1(_04259_),
    .C1(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__and3_1 _11382_ (.A(curr_PC[12]),
    .B(curr_PC[13]),
    .C(_04056_),
    .X(_04289_));
 sky130_fd_sc_hd__o21ai_1 _11383_ (.A1(curr_PC[13]),
    .A2(_04173_),
    .B1(net242),
    .Y(_04290_));
 sky130_fd_sc_hd__a2bb2o_4 _11384_ (.A1_N(_04289_),
    .A2_N(_04290_),
    .B1(net238),
    .B2(_04288_),
    .X(dest_val[13]));
 sky130_fd_sc_hd__o21ai_1 _11385_ (.A1(_04175_),
    .A2(_04254_),
    .B1(net136),
    .Y(_04291_));
 sky130_fd_sc_hd__a21bo_1 _11386_ (.A1(_04229_),
    .A2(_04238_),
    .B1_N(_04237_),
    .X(_04292_));
 sky130_fd_sc_hd__o21ai_1 _11387_ (.A1(_04200_),
    .A2(_04207_),
    .B1(_04205_),
    .Y(_04293_));
 sky130_fd_sc_hd__nand2_1 _11388_ (.A(_04180_),
    .B(_04185_),
    .Y(_04294_));
 sky130_fd_sc_hd__a21boi_1 _11389_ (.A1(_04188_),
    .A2(_04194_),
    .B1_N(_04193_),
    .Y(_04295_));
 sky130_fd_sc_hd__a21o_1 _11390_ (.A1(_04180_),
    .A2(_04185_),
    .B1(_04295_),
    .X(_04296_));
 sky130_fd_sc_hd__xnor2_1 _11391_ (.A(_04294_),
    .B(_04295_),
    .Y(_04297_));
 sky130_fd_sc_hd__xnor2_1 _11392_ (.A(_04293_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__o22a_1 _11393_ (.A1(net50),
    .A2(net20),
    .B1(net18),
    .B2(net52),
    .X(_04299_));
 sky130_fd_sc_hd__xnor2_1 _11394_ (.A(_00274_),
    .B(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__o22a_1 _11395_ (.A1(net48),
    .A2(net38),
    .B1(net36),
    .B2(net46),
    .X(_04301_));
 sky130_fd_sc_hd__xnor2_1 _11396_ (.A(_00262_),
    .B(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__o22a_1 _11397_ (.A1(net44),
    .A2(net29),
    .B1(net27),
    .B2(_00517_),
    .X(_04303_));
 sky130_fd_sc_hd__xnor2_1 _11398_ (.A(net90),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__nand2_1 _11399_ (.A(_04302_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__xnor2_1 _11400_ (.A(_04302_),
    .B(_04304_),
    .Y(_04306_));
 sky130_fd_sc_hd__xnor2_1 _11401_ (.A(_04300_),
    .B(_04306_),
    .Y(_04307_));
 sky130_fd_sc_hd__a22o_1 _11402_ (.A1(_06725_),
    .A2(net15),
    .B1(net31),
    .B2(net55),
    .X(_04308_));
 sky130_fd_sc_hd__xnor2_1 _11403_ (.A(net91),
    .B(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__o22a_1 _11404_ (.A1(_00202_),
    .A2(net34),
    .B1(net32),
    .B2(net41),
    .X(_04310_));
 sky130_fd_sc_hd__xnor2_1 _11405_ (.A(net93),
    .B(_04310_),
    .Y(_04311_));
 sky130_fd_sc_hd__nand2_1 _11406_ (.A(_04309_),
    .B(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__xnor2_1 _11407_ (.A(_04309_),
    .B(_04311_),
    .Y(_04313_));
 sky130_fd_sc_hd__o22a_1 _11408_ (.A1(net25),
    .A2(_00811_),
    .B1(_02066_),
    .B2(net23),
    .X(_04314_));
 sky130_fd_sc_hd__xnor2_1 _11409_ (.A(net87),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__or2_1 _11410_ (.A(_00439_),
    .B(net5),
    .X(_04316_));
 sky130_fd_sc_hd__a22o_2 _11411_ (.A1(_00438_),
    .A2(net7),
    .B1(_04316_),
    .B2(net117),
    .X(_04317_));
 sky130_fd_sc_hd__nor2_1 _11412_ (.A(_04315_),
    .B(_04317_),
    .Y(_04318_));
 sky130_fd_sc_hd__xor2_1 _11413_ (.A(_04315_),
    .B(_04317_),
    .X(_04319_));
 sky130_fd_sc_hd__nor2_1 _11414_ (.A(_04313_),
    .B(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__xnor2_1 _11415_ (.A(_04313_),
    .B(_04319_),
    .Y(_04321_));
 sky130_fd_sc_hd__nor2_1 _11416_ (.A(_04307_),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__and2_1 _11417_ (.A(_04307_),
    .B(_04321_),
    .X(_04323_));
 sky130_fd_sc_hd__or2_1 _11418_ (.A(_04322_),
    .B(_04323_),
    .X(_04324_));
 sky130_fd_sc_hd__a22o_1 _11419_ (.A1(net71),
    .A2(net9),
    .B1(net3),
    .B2(net73),
    .X(_04325_));
 sky130_fd_sc_hd__xnor2_1 _11420_ (.A(net62),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__a22o_1 _11421_ (.A1(net101),
    .A2(net16),
    .B1(net12),
    .B2(net102),
    .X(_04327_));
 sky130_fd_sc_hd__xnor2_1 _11422_ (.A(net64),
    .B(_04327_),
    .Y(_04328_));
 sky130_fd_sc_hd__nor2_1 _11423_ (.A(net77),
    .B(net59),
    .Y(_04329_));
 sky130_fd_sc_hd__xnor2_1 _11424_ (.A(_04328_),
    .B(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__nor2_1 _11425_ (.A(_04326_),
    .B(_04330_),
    .Y(_04331_));
 sky130_fd_sc_hd__and2_1 _11426_ (.A(_04326_),
    .B(_04330_),
    .X(_04332_));
 sky130_fd_sc_hd__or2_1 _11427_ (.A(_04331_),
    .B(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__xnor2_1 _11428_ (.A(_04324_),
    .B(_04333_),
    .Y(_04334_));
 sky130_fd_sc_hd__or2_1 _11429_ (.A(_04298_),
    .B(_04334_),
    .X(_04335_));
 sky130_fd_sc_hd__nand2_1 _11430_ (.A(_04298_),
    .B(_04334_),
    .Y(_04336_));
 sky130_fd_sc_hd__and2_1 _11431_ (.A(_04335_),
    .B(_04336_),
    .X(_04337_));
 sky130_fd_sc_hd__a21bo_1 _11432_ (.A1(_04219_),
    .A2(_04225_),
    .B1_N(_04218_),
    .X(_04338_));
 sky130_fd_sc_hd__a21boi_2 _11433_ (.A1(_04198_),
    .A2(_04208_),
    .B1_N(_04197_),
    .Y(_04339_));
 sky130_fd_sc_hd__o21a_1 _11434_ (.A1(_04215_),
    .A2(_04216_),
    .B1(_04213_),
    .X(_04340_));
 sky130_fd_sc_hd__or2_1 _11435_ (.A(_04339_),
    .B(_04340_),
    .X(_04341_));
 sky130_fd_sc_hd__xnor2_1 _11436_ (.A(_04339_),
    .B(_04340_),
    .Y(_04342_));
 sky130_fd_sc_hd__a21o_1 _11437_ (.A1(_04221_),
    .A2(_04224_),
    .B1(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__nand3_1 _11438_ (.A(_04221_),
    .B(_04224_),
    .C(_04342_),
    .Y(_04344_));
 sky130_fd_sc_hd__nand2_1 _11439_ (.A(_04343_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__nor2_1 _11440_ (.A(_04232_),
    .B(_04235_),
    .Y(_04346_));
 sky130_fd_sc_hd__xnor2_1 _11441_ (.A(_04345_),
    .B(_04346_),
    .Y(_04347_));
 sky130_fd_sc_hd__nand2b_1 _11442_ (.A_N(_04347_),
    .B(_04338_),
    .Y(_04348_));
 sky130_fd_sc_hd__xnor2_1 _11443_ (.A(_04338_),
    .B(_04347_),
    .Y(_04349_));
 sky130_fd_sc_hd__nand2_1 _11444_ (.A(_04337_),
    .B(_04349_),
    .Y(_04350_));
 sky130_fd_sc_hd__xnor2_1 _11445_ (.A(_04337_),
    .B(_04349_),
    .Y(_04351_));
 sky130_fd_sc_hd__nand2b_2 _11446_ (.A_N(_04351_),
    .B(_04292_),
    .Y(_04352_));
 sky130_fd_sc_hd__xor2_1 _11447_ (.A(_04292_),
    .B(_04351_),
    .X(_04353_));
 sky130_fd_sc_hd__a21oi_2 _11448_ (.A1(_04240_),
    .A2(_04243_),
    .B1(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__and3_1 _11449_ (.A(_04240_),
    .B(_04243_),
    .C(_04353_),
    .X(_04355_));
 sky130_fd_sc_hd__or2_4 _11450_ (.A(_04354_),
    .B(_04355_),
    .X(_04356_));
 sky130_fd_sc_hd__a21oi_2 _11451_ (.A1(_04129_),
    .A2(_04246_),
    .B1(_04247_),
    .Y(_04357_));
 sky130_fd_sc_hd__nor2_1 _11452_ (.A(_04131_),
    .B(_04248_),
    .Y(_04358_));
 sky130_fd_sc_hd__a21o_1 _11453_ (.A1(_04132_),
    .A2(_04358_),
    .B1(_04357_),
    .X(_04359_));
 sky130_fd_sc_hd__nand2_1 _11454_ (.A(_04133_),
    .B(_04358_),
    .Y(_04360_));
 sky130_fd_sc_hd__o21ba_1 _11455_ (.A1(_03893_),
    .A2(_04360_),
    .B1_N(_04359_),
    .X(_04361_));
 sky130_fd_sc_hd__xnor2_4 _11456_ (.A(_04356_),
    .B(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__inv_2 _11457_ (.A(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__or2_1 _11458_ (.A(_04291_),
    .B(_04362_),
    .X(_04364_));
 sky130_fd_sc_hd__a21oi_1 _11459_ (.A1(_04291_),
    .A2(_04362_),
    .B1(net235),
    .Y(_04365_));
 sky130_fd_sc_hd__and2_1 _11460_ (.A(net136),
    .B(_01954_),
    .X(_04366_));
 sky130_fd_sc_hd__xnor2_1 _11461_ (.A(_01959_),
    .B(_04366_),
    .Y(_04367_));
 sky130_fd_sc_hd__o21a_1 _11462_ (.A1(_06339_),
    .A2(_04260_),
    .B1(_06333_),
    .X(_04368_));
 sky130_fd_sc_hd__nor2_1 _11463_ (.A(net293),
    .B(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__a31o_1 _11464_ (.A1(net293),
    .A2(_06321_),
    .A3(_06591_),
    .B1(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__nand2_1 _11465_ (.A(_06291_),
    .B(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__o211a_1 _11466_ (.A1(_06291_),
    .A2(_04370_),
    .B1(_04371_),
    .C1(net234),
    .X(_04372_));
 sky130_fd_sc_hd__or2_1 _11467_ (.A(reg1_val[14]),
    .B(curr_PC[14]),
    .X(_04373_));
 sky130_fd_sc_hd__nand2_1 _11468_ (.A(reg1_val[14]),
    .B(curr_PC[14]),
    .Y(_04374_));
 sky130_fd_sc_hd__nand2_1 _11469_ (.A(_04373_),
    .B(_04374_),
    .Y(_04375_));
 sky130_fd_sc_hd__o21a_1 _11470_ (.A1(_04267_),
    .A2(_04268_),
    .B1(_04266_),
    .X(_04376_));
 sky130_fd_sc_hd__xor2_1 _11471_ (.A(_04375_),
    .B(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__mux2_1 _11472_ (.A0(_03368_),
    .A1(_03370_),
    .S(net219),
    .X(_04378_));
 sky130_fd_sc_hd__mux2_1 _11473_ (.A0(_02633_),
    .A1(_04378_),
    .S(net220),
    .X(_04379_));
 sky130_fd_sc_hd__mux2_1 _11474_ (.A0(_04377_),
    .A1(_04379_),
    .S(net224),
    .X(_04380_));
 sky130_fd_sc_hd__o21ai_1 _11475_ (.A1(\div_shifter[45] ),
    .A2(_04276_),
    .B1(net227),
    .Y(_04381_));
 sky130_fd_sc_hd__xnor2_1 _11476_ (.A(\div_shifter[46] ),
    .B(_04381_),
    .Y(_04382_));
 sky130_fd_sc_hd__o21ai_1 _11477_ (.A1(\div_res[13] ),
    .A2(_04273_),
    .B1(net139),
    .Y(_04383_));
 sky130_fd_sc_hd__xnor2_1 _11478_ (.A(\div_res[14] ),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__o21ai_1 _11479_ (.A1(reg1_val[14]),
    .A2(_06240_),
    .B1(net193),
    .Y(_04385_));
 sky130_fd_sc_hd__o221a_1 _11480_ (.A1(_06251_),
    .A2(net204),
    .B1(net231),
    .B2(reg1_val[14]),
    .C1(_04385_),
    .X(_04386_));
 sky130_fd_sc_hd__o221ai_4 _11481_ (.A1(_06297_),
    .A2(_02429_),
    .B1(net194),
    .B2(_06284_),
    .C1(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__a221o_1 _11482_ (.A1(_00433_),
    .A2(net257),
    .B1(_02443_),
    .B2(_04384_),
    .C1(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__a21o_1 _11483_ (.A1(_02441_),
    .A2(_04382_),
    .B1(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__o21a_1 _11484_ (.A1(net221),
    .A2(_02610_),
    .B1(_02456_),
    .X(_04390_));
 sky130_fd_sc_hd__a221o_1 _11485_ (.A1(net167),
    .A2(_04379_),
    .B1(_04390_),
    .B2(net171),
    .C1(_04389_),
    .X(_04391_));
 sky130_fd_sc_hd__a211o_1 _11486_ (.A1(net205),
    .A2(_04380_),
    .B1(_04391_),
    .C1(_04372_),
    .X(_04392_));
 sky130_fd_sc_hd__a221o_1 _11487_ (.A1(_04364_),
    .A2(_04365_),
    .B1(_04367_),
    .B2(net233),
    .C1(_04392_),
    .X(_04393_));
 sky130_fd_sc_hd__or2_1 _11488_ (.A(curr_PC[14]),
    .B(_04289_),
    .X(_04394_));
 sky130_fd_sc_hd__and2_1 _11489_ (.A(curr_PC[14]),
    .B(_04289_),
    .X(_04395_));
 sky130_fd_sc_hd__nor2_1 _11490_ (.A(net238),
    .B(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__a22o_4 _11491_ (.A1(net238),
    .A2(_04393_),
    .B1(_04394_),
    .B2(_04396_),
    .X(dest_val[14]));
 sky130_fd_sc_hd__o31ai_1 _11492_ (.A1(_04175_),
    .A2(_04254_),
    .A3(_04363_),
    .B1(net136),
    .Y(_04397_));
 sky130_fd_sc_hd__a22o_1 _11493_ (.A1(net102),
    .A2(net8),
    .B1(net3),
    .B2(net71),
    .X(_04398_));
 sky130_fd_sc_hd__xnor2_1 _11494_ (.A(net59),
    .B(_04398_),
    .Y(_04399_));
 sky130_fd_sc_hd__o22a_1 _11495_ (.A1(net41),
    .A2(net34),
    .B1(net32),
    .B2(net57),
    .X(_04400_));
 sky130_fd_sc_hd__xnor2_1 _11496_ (.A(net94),
    .B(_04400_),
    .Y(_04402_));
 sky130_fd_sc_hd__and2_1 _11497_ (.A(_04399_),
    .B(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__nor2_1 _11498_ (.A(_04399_),
    .B(_04402_),
    .Y(_04404_));
 sky130_fd_sc_hd__or2_1 _11499_ (.A(_04403_),
    .B(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__a22o_1 _11500_ (.A1(_00203_),
    .A2(net17),
    .B1(net12),
    .B2(net101),
    .X(_04406_));
 sky130_fd_sc_hd__xnor2_2 _11501_ (.A(net65),
    .B(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__and2b_1 _11502_ (.A_N(_04405_),
    .B(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__xnor2_2 _11503_ (.A(_04405_),
    .B(_04407_),
    .Y(_04409_));
 sky130_fd_sc_hd__o22a_1 _11504_ (.A1(net25),
    .A2(_02066_),
    .B1(_02176_),
    .B2(net23),
    .X(_04410_));
 sky130_fd_sc_hd__xnor2_2 _11505_ (.A(net87),
    .B(_04410_),
    .Y(_04411_));
 sky130_fd_sc_hd__o22a_1 _11506_ (.A1(net29),
    .A2(_00517_),
    .B1(_00811_),
    .B2(net27),
    .X(_04413_));
 sky130_fd_sc_hd__xnor2_2 _11507_ (.A(net90),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__xnor2_2 _11508_ (.A(net118),
    .B(_04414_),
    .Y(_04415_));
 sky130_fd_sc_hd__and2_1 _11509_ (.A(_04411_),
    .B(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__xnor2_2 _11510_ (.A(_04411_),
    .B(_04415_),
    .Y(_04417_));
 sky130_fd_sc_hd__o22a_1 _11511_ (.A1(net52),
    .A2(net20),
    .B1(net18),
    .B2(net43),
    .X(_04418_));
 sky130_fd_sc_hd__xnor2_2 _11512_ (.A(_00273_),
    .B(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__o22a_1 _11513_ (.A1(net54),
    .A2(_00336_),
    .B1(_00342_),
    .B2(net48),
    .X(_04420_));
 sky130_fd_sc_hd__xnor2_2 _11514_ (.A(_00308_),
    .B(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__nand2_1 _11515_ (.A(_04419_),
    .B(_04421_),
    .Y(_04422_));
 sky130_fd_sc_hd__xnor2_2 _11516_ (.A(_04419_),
    .B(_04421_),
    .Y(_04424_));
 sky130_fd_sc_hd__o22a_1 _11517_ (.A1(net46),
    .A2(net38),
    .B1(net36),
    .B2(net50),
    .X(_04425_));
 sky130_fd_sc_hd__xnor2_2 _11518_ (.A(net98),
    .B(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__nand2b_1 _11519_ (.A_N(_04424_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__xnor2_2 _11520_ (.A(_04424_),
    .B(_04426_),
    .Y(_04428_));
 sky130_fd_sc_hd__and3_1 _11521_ (.A(_04309_),
    .B(_04311_),
    .C(_04428_),
    .X(_04429_));
 sky130_fd_sc_hd__xnor2_2 _11522_ (.A(_04312_),
    .B(_04428_),
    .Y(_04430_));
 sky130_fd_sc_hd__and2b_1 _11523_ (.A_N(_04417_),
    .B(_04430_),
    .X(_04431_));
 sky130_fd_sc_hd__xnor2_2 _11524_ (.A(_04417_),
    .B(_04430_),
    .Y(_04432_));
 sky130_fd_sc_hd__xnor2_2 _11525_ (.A(_04409_),
    .B(_04432_),
    .Y(_04433_));
 sky130_fd_sc_hd__o21a_1 _11526_ (.A1(_04300_),
    .A2(_04306_),
    .B1(_04305_),
    .X(_04435_));
 sky130_fd_sc_hd__nand2_1 _11527_ (.A(net73),
    .B(net62),
    .Y(_04436_));
 sky130_fd_sc_hd__xnor2_1 _11528_ (.A(_04435_),
    .B(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__nor2_1 _11529_ (.A(_04318_),
    .B(_04437_),
    .Y(_04438_));
 sky130_fd_sc_hd__and2_1 _11530_ (.A(_04318_),
    .B(_04437_),
    .X(_04439_));
 sky130_fd_sc_hd__nor2_1 _11531_ (.A(_04438_),
    .B(_04439_),
    .Y(_04440_));
 sky130_fd_sc_hd__nand2b_1 _11532_ (.A_N(_04433_),
    .B(_04440_),
    .Y(_04441_));
 sky130_fd_sc_hd__xnor2_2 _11533_ (.A(_04433_),
    .B(_04440_),
    .Y(_04442_));
 sky130_fd_sc_hd__o21a_1 _11534_ (.A1(_04324_),
    .A2(_04333_),
    .B1(_04335_),
    .X(_04443_));
 sky130_fd_sc_hd__a21bo_1 _11535_ (.A1(_04293_),
    .A2(_04297_),
    .B1_N(_04296_),
    .X(_04444_));
 sky130_fd_sc_hd__a21oi_1 _11536_ (.A1(_04328_),
    .A2(_04329_),
    .B1(_04331_),
    .Y(_04446_));
 sky130_fd_sc_hd__o21ba_1 _11537_ (.A1(_04320_),
    .A2(_04322_),
    .B1_N(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__or3b_1 _11538_ (.A(_04320_),
    .B(_04322_),
    .C_N(_04446_),
    .X(_04448_));
 sky130_fd_sc_hd__and2b_1 _11539_ (.A_N(_04447_),
    .B(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__xnor2_1 _11540_ (.A(_04444_),
    .B(_04449_),
    .Y(_04450_));
 sky130_fd_sc_hd__a21oi_1 _11541_ (.A1(_04341_),
    .A2(_04343_),
    .B1(_04450_),
    .Y(_04451_));
 sky130_fd_sc_hd__and3_1 _11542_ (.A(_04341_),
    .B(_04343_),
    .C(_04450_),
    .X(_04452_));
 sky130_fd_sc_hd__nor2_1 _11543_ (.A(_04451_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__xnor2_2 _11544_ (.A(_04443_),
    .B(_04453_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand2_1 _11545_ (.A(_04442_),
    .B(_04454_),
    .Y(_04455_));
 sky130_fd_sc_hd__xnor2_2 _11546_ (.A(_04442_),
    .B(_04454_),
    .Y(_04457_));
 sky130_fd_sc_hd__o21ai_2 _11547_ (.A1(_04345_),
    .A2(_04346_),
    .B1(_04348_),
    .Y(_04458_));
 sky130_fd_sc_hd__nand2b_1 _11548_ (.A_N(_04457_),
    .B(_04458_),
    .Y(_04459_));
 sky130_fd_sc_hd__xor2_2 _11549_ (.A(_04457_),
    .B(_04458_),
    .X(_04460_));
 sky130_fd_sc_hd__a21oi_2 _11550_ (.A1(_04350_),
    .A2(_04352_),
    .B1(_04460_),
    .Y(_04461_));
 sky130_fd_sc_hd__nand3_4 _11551_ (.A(_04350_),
    .B(_04352_),
    .C(_04460_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand2b_4 _11552_ (.A_N(_04461_),
    .B(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__o21ba_1 _11553_ (.A1(_04245_),
    .A2(_04354_),
    .B1_N(_04355_),
    .X(_04464_));
 sky130_fd_sc_hd__nor2_2 _11554_ (.A(_04248_),
    .B(_04356_),
    .Y(_04465_));
 sky130_fd_sc_hd__a21oi_1 _11555_ (.A1(_04251_),
    .A2(_04465_),
    .B1(_04464_),
    .Y(_04466_));
 sky130_fd_sc_hd__nand2_2 _11556_ (.A(_04249_),
    .B(_04465_),
    .Y(_04468_));
 sky130_fd_sc_hd__a311o_1 _11557_ (.A1(_03491_),
    .A2(_03492_),
    .A3(_03494_),
    .B1(_04016_),
    .C1(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__o211ai_4 _11558_ (.A1(_04020_),
    .A2(_04468_),
    .B1(_04469_),
    .C1(_04466_),
    .Y(_04470_));
 sky130_fd_sc_hd__xor2_4 _11559_ (.A(_04463_),
    .B(_04470_),
    .X(_04471_));
 sky130_fd_sc_hd__and2_1 _11560_ (.A(_04397_),
    .B(_04471_),
    .X(_04472_));
 sky130_fd_sc_hd__nor2_1 _11561_ (.A(_04397_),
    .B(_04471_),
    .Y(_04473_));
 sky130_fd_sc_hd__or2_1 _11562_ (.A(net134),
    .B(_01960_),
    .X(_04474_));
 sky130_fd_sc_hd__o21ai_1 _11563_ (.A1(_01961_),
    .A2(_04474_),
    .B1(net233),
    .Y(_04475_));
 sky130_fd_sc_hd__a21o_1 _11564_ (.A1(_01961_),
    .A2(_04474_),
    .B1(_04475_),
    .X(_04476_));
 sky130_fd_sc_hd__o21a_1 _11565_ (.A1(_06297_),
    .A2(_04368_),
    .B1(_06284_),
    .X(_04477_));
 sky130_fd_sc_hd__nor2_1 _11566_ (.A(net294),
    .B(_04477_),
    .Y(_04479_));
 sky130_fd_sc_hd__a31o_1 _11567_ (.A1(net294),
    .A2(_06262_),
    .A3(_06592_),
    .B1(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__o21a_1 _11568_ (.A1(_06207_),
    .A2(_04480_),
    .B1(net234),
    .X(_04481_));
 sky130_fd_sc_hd__a21bo_1 _11569_ (.A1(_06207_),
    .A2(_04480_),
    .B1_N(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__or2_1 _11570_ (.A(reg1_val[15]),
    .B(curr_PC[15]),
    .X(_04483_));
 sky130_fd_sc_hd__nand2_1 _11571_ (.A(reg1_val[15]),
    .B(curr_PC[15]),
    .Y(_04484_));
 sky130_fd_sc_hd__nand2_1 _11572_ (.A(_04483_),
    .B(_04484_),
    .Y(_04485_));
 sky130_fd_sc_hd__o21a_1 _11573_ (.A1(_04375_),
    .A2(_04376_),
    .B1(_04374_),
    .X(_04486_));
 sky130_fd_sc_hd__xnor2_1 _11574_ (.A(_04485_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__mux2_1 _11575_ (.A0(_03511_),
    .A1(_03513_),
    .S(net218),
    .X(_04488_));
 sky130_fd_sc_hd__or2_1 _11576_ (.A(net220),
    .B(_02454_),
    .X(_04490_));
 sky130_fd_sc_hd__o21ai_2 _11577_ (.A1(net221),
    .A2(_04488_),
    .B1(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__mux2_1 _11578_ (.A0(_04487_),
    .A1(_04491_),
    .S(net224),
    .X(_04492_));
 sky130_fd_sc_hd__or3_2 _11579_ (.A(\div_shifter[46] ),
    .B(\div_shifter[45] ),
    .C(_04276_),
    .X(_04493_));
 sky130_fd_sc_hd__and3_1 _11580_ (.A(\div_shifter[47] ),
    .B(net227),
    .C(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__a21oi_1 _11581_ (.A1(net227),
    .A2(_04493_),
    .B1(\div_shifter[47] ),
    .Y(_04495_));
 sky130_fd_sc_hd__or3_1 _11582_ (.A(\div_res[14] ),
    .B(\div_res[13] ),
    .C(_04273_),
    .X(_04496_));
 sky130_fd_sc_hd__a21oi_1 _11583_ (.A1(net139),
    .A2(_04496_),
    .B1(\div_res[15] ),
    .Y(_04497_));
 sky130_fd_sc_hd__a31o_1 _11584_ (.A1(\div_res[15] ),
    .A2(net139),
    .A3(_04496_),
    .B1(net189),
    .X(_04498_));
 sky130_fd_sc_hd__nand2_1 _11585_ (.A(_00379_),
    .B(net256),
    .Y(_04499_));
 sky130_fd_sc_hd__nand2_1 _11586_ (.A(_06185_),
    .B(net193),
    .Y(_04501_));
 sky130_fd_sc_hd__o221a_1 _11587_ (.A1(_06196_),
    .A2(net194),
    .B1(net231),
    .B2(reg1_val[15]),
    .C1(_04501_),
    .X(_04502_));
 sky130_fd_sc_hd__o211a_1 _11588_ (.A1(_06218_),
    .A2(_02429_),
    .B1(_04499_),
    .C1(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__o21a_1 _11589_ (.A1(_04497_),
    .A2(_04498_),
    .B1(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__o31a_1 _11590_ (.A1(net191),
    .A2(_04494_),
    .A3(_04495_),
    .B1(_04504_),
    .X(_04505_));
 sky130_fd_sc_hd__o21a_1 _11591_ (.A1(net221),
    .A2(_02417_),
    .B1(_02456_),
    .X(_04506_));
 sky130_fd_sc_hd__inv_2 _11592_ (.A(_04506_),
    .Y(_04507_));
 sky130_fd_sc_hd__o221a_1 _11593_ (.A1(_02425_),
    .A2(_04491_),
    .B1(_04507_),
    .B2(net168),
    .C1(_04505_),
    .X(_04508_));
 sky130_fd_sc_hd__o211a_1 _11594_ (.A1(_06667_),
    .A2(_04492_),
    .B1(_04508_),
    .C1(_04482_),
    .X(_04509_));
 sky130_fd_sc_hd__o311a_1 _11595_ (.A1(net235),
    .A2(_04472_),
    .A3(_04473_),
    .B1(_04476_),
    .C1(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__a2bb2o_1 _11596_ (.A1_N(_06679_),
    .A2_N(_04510_),
    .B1(_06165_),
    .B2(_06677_),
    .X(_04512_));
 sky130_fd_sc_hd__and3_2 _11597_ (.A(curr_PC[14]),
    .B(curr_PC[15]),
    .C(_04289_),
    .X(_04513_));
 sky130_fd_sc_hd__o21ai_1 _11598_ (.A1(curr_PC[15]),
    .A2(_04395_),
    .B1(net242),
    .Y(_04514_));
 sky130_fd_sc_hd__a2bb2o_4 _11599_ (.A1_N(_04513_),
    .A2_N(_04514_),
    .B1(net238),
    .B2(_04512_),
    .X(dest_val[15]));
 sky130_fd_sc_hd__or4bb_1 _11600_ (.A(_04137_),
    .B(_04254_),
    .C_N(_04362_),
    .D_N(_04471_),
    .X(_04515_));
 sky130_fd_sc_hd__or2_1 _11601_ (.A(_04059_),
    .B(_04515_),
    .X(_04516_));
 sky130_fd_sc_hd__o22a_1 _11602_ (.A1(net50),
    .A2(net38),
    .B1(net36),
    .B2(net52),
    .X(_04517_));
 sky130_fd_sc_hd__xnor2_1 _11603_ (.A(_00262_),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__o22a_1 _11604_ (.A1(net43),
    .A2(net20),
    .B1(net18),
    .B2(_00517_),
    .X(_04519_));
 sky130_fd_sc_hd__xnor2_1 _11605_ (.A(net97),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _11606_ (.A(_04518_),
    .B(_04520_),
    .Y(_04522_));
 sky130_fd_sc_hd__or2_1 _11607_ (.A(_04518_),
    .B(_04520_),
    .X(_04523_));
 sky130_fd_sc_hd__nand2_1 _11608_ (.A(_04522_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__a21oi_1 _11609_ (.A1(_04422_),
    .A2(_04427_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__and3_1 _11610_ (.A(_04422_),
    .B(_04427_),
    .C(_04524_),
    .X(_04526_));
 sky130_fd_sc_hd__or2_1 _11611_ (.A(_04525_),
    .B(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__o22a_1 _11612_ (.A1(net29),
    .A2(_00811_),
    .B1(_02066_),
    .B2(net27),
    .X(_04528_));
 sky130_fd_sc_hd__xnor2_1 _11613_ (.A(net89),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__a21oi_1 _11614_ (.A1(_00386_),
    .A2(net7),
    .B1(_00359_),
    .Y(_04530_));
 sky130_fd_sc_hd__a31o_1 _11615_ (.A1(_00359_),
    .A2(_00384_),
    .A3(net7),
    .B1(_04530_),
    .X(_04531_));
 sky130_fd_sc_hd__nor2_1 _11616_ (.A(_04529_),
    .B(_04531_),
    .Y(_04533_));
 sky130_fd_sc_hd__and2_1 _11617_ (.A(_04529_),
    .B(_04531_),
    .X(_04534_));
 sky130_fd_sc_hd__nor2_1 _11618_ (.A(_04533_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__xnor2_1 _11619_ (.A(_04527_),
    .B(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__o22a_1 _11620_ (.A1(net57),
    .A2(net34),
    .B1(net32),
    .B2(net54),
    .X(_04537_));
 sky130_fd_sc_hd__xnor2_1 _11621_ (.A(net93),
    .B(_04537_),
    .Y(_04538_));
 sky130_fd_sc_hd__inv_2 _11622_ (.A(_04538_),
    .Y(_04539_));
 sky130_fd_sc_hd__a22o_1 _11623_ (.A1(_00208_),
    .A2(net17),
    .B1(net13),
    .B2(_00203_),
    .X(_04540_));
 sky130_fd_sc_hd__xnor2_1 _11624_ (.A(net65),
    .B(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__a22o_1 _11625_ (.A1(_00150_),
    .A2(net15),
    .B1(net31),
    .B2(_00161_),
    .X(_04542_));
 sky130_fd_sc_hd__xnor2_1 _11626_ (.A(net91),
    .B(_04542_),
    .Y(_04544_));
 sky130_fd_sc_hd__and2_1 _11627_ (.A(_04541_),
    .B(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__nor2_1 _11628_ (.A(_04541_),
    .B(_04544_),
    .Y(_04546_));
 sky130_fd_sc_hd__or2_1 _11629_ (.A(_04545_),
    .B(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__nor2_1 _11630_ (.A(_04539_),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__and2_1 _11631_ (.A(_04539_),
    .B(_04547_),
    .X(_04549_));
 sky130_fd_sc_hd__or2_1 _11632_ (.A(_04548_),
    .B(_04549_),
    .X(_04550_));
 sky130_fd_sc_hd__xnor2_1 _11633_ (.A(_04536_),
    .B(_04550_),
    .Y(_04551_));
 sky130_fd_sc_hd__a21o_1 _11634_ (.A1(_00381_),
    .A2(_04414_),
    .B1(_04416_),
    .X(_04552_));
 sky130_fd_sc_hd__a22o_1 _11635_ (.A1(net101),
    .A2(_02080_),
    .B1(net4),
    .B2(net102),
    .X(_04553_));
 sky130_fd_sc_hd__xnor2_1 _11636_ (.A(net59),
    .B(_04553_),
    .Y(_04555_));
 sky130_fd_sc_hd__xor2_1 _11637_ (.A(_04552_),
    .B(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__and3_1 _11638_ (.A(net71),
    .B(net62),
    .C(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__a21oi_1 _11639_ (.A1(_00467_),
    .A2(net62),
    .B1(_04556_),
    .Y(_04558_));
 sky130_fd_sc_hd__nor2_1 _11640_ (.A(_04557_),
    .B(_04558_),
    .Y(_04559_));
 sky130_fd_sc_hd__and2b_1 _11641_ (.A_N(_04551_),
    .B(_04559_),
    .X(_04560_));
 sky130_fd_sc_hd__xnor2_1 _11642_ (.A(_04551_),
    .B(_04559_),
    .Y(_04561_));
 sky130_fd_sc_hd__a21bo_1 _11643_ (.A1(_04409_),
    .A2(_04432_),
    .B1_N(_04441_),
    .X(_04562_));
 sky130_fd_sc_hd__o21bai_2 _11644_ (.A1(_04435_),
    .A2(_04436_),
    .B1_N(_04438_),
    .Y(_04563_));
 sky130_fd_sc_hd__o22ai_1 _11645_ (.A1(_04403_),
    .A2(_04408_),
    .B1(_04429_),
    .B2(_04431_),
    .Y(_04564_));
 sky130_fd_sc_hd__or4_1 _11646_ (.A(_04403_),
    .B(_04408_),
    .C(_04429_),
    .D(_04431_),
    .X(_04566_));
 sky130_fd_sc_hd__and2_1 _11647_ (.A(_04564_),
    .B(_04566_),
    .X(_04567_));
 sky130_fd_sc_hd__xnor2_2 _11648_ (.A(_04563_),
    .B(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__a21oi_2 _11649_ (.A1(_04444_),
    .A2(_04448_),
    .B1(_04447_),
    .Y(_04569_));
 sky130_fd_sc_hd__xnor2_1 _11650_ (.A(_04568_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__nand2b_1 _11651_ (.A_N(_04570_),
    .B(_04562_),
    .Y(_04571_));
 sky130_fd_sc_hd__xnor2_1 _11652_ (.A(_04562_),
    .B(_04570_),
    .Y(_04572_));
 sky130_fd_sc_hd__nand2_1 _11653_ (.A(_04561_),
    .B(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__xnor2_1 _11654_ (.A(_04561_),
    .B(_04572_),
    .Y(_04574_));
 sky130_fd_sc_hd__o21ba_1 _11655_ (.A1(_04443_),
    .A2(_04452_),
    .B1_N(_04451_),
    .X(_04575_));
 sky130_fd_sc_hd__or2_1 _11656_ (.A(_04574_),
    .B(_04575_),
    .X(_04577_));
 sky130_fd_sc_hd__nand2_1 _11657_ (.A(_04574_),
    .B(_04575_),
    .Y(_04578_));
 sky130_fd_sc_hd__nand2_1 _11658_ (.A(_04577_),
    .B(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__a21oi_2 _11659_ (.A1(_04455_),
    .A2(_04459_),
    .B1(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__nand3_2 _11660_ (.A(_04455_),
    .B(_04459_),
    .C(_04579_),
    .Y(_04581_));
 sky130_fd_sc_hd__nand2b_2 _11661_ (.A_N(_04580_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__o21a_1 _11662_ (.A1(_04354_),
    .A2(_04461_),
    .B1(_04462_),
    .X(_04583_));
 sky130_fd_sc_hd__nor2_1 _11663_ (.A(_04356_),
    .B(_04463_),
    .Y(_04584_));
 sky130_fd_sc_hd__a21o_1 _11664_ (.A1(_04357_),
    .A2(_04584_),
    .B1(_04583_),
    .X(_04585_));
 sky130_fd_sc_hd__nand2_1 _11665_ (.A(_04358_),
    .B(_04584_),
    .Y(_04586_));
 sky130_fd_sc_hd__a31oi_2 _11666_ (.A1(_04134_),
    .A2(_04358_),
    .A3(_04584_),
    .B1(_04585_),
    .Y(_04588_));
 sky130_fd_sc_hd__o31ai_4 _11667_ (.A1(_03545_),
    .A2(_04135_),
    .A3(_04586_),
    .B1(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__xnor2_4 _11668_ (.A(_04582_),
    .B(_04589_),
    .Y(_04590_));
 sky130_fd_sc_hd__a21oi_1 _11669_ (.A1(net144),
    .A2(_04516_),
    .B1(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__a31o_1 _11670_ (.A1(net144),
    .A2(_04516_),
    .A3(_04590_),
    .B1(net235),
    .X(_04592_));
 sky130_fd_sc_hd__a21o_1 _11671_ (.A1(_01960_),
    .A2(_01961_),
    .B1(net134),
    .X(_04593_));
 sky130_fd_sc_hd__xnor2_2 _11672_ (.A(_01967_),
    .B(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__o21ai_1 _11673_ (.A1(_06218_),
    .A2(_04477_),
    .B1(_06196_),
    .Y(_04595_));
 sky130_fd_sc_hd__and2_1 _11674_ (.A(net283),
    .B(_04595_),
    .X(_04596_));
 sky130_fd_sc_hd__and3_1 _11675_ (.A(net294),
    .B(_06174_),
    .C(_06593_),
    .X(_04597_));
 sky130_fd_sc_hd__o21ai_1 _11676_ (.A1(_04596_),
    .A2(_04597_),
    .B1(_06153_),
    .Y(_04599_));
 sky130_fd_sc_hd__o31a_1 _11677_ (.A1(_06153_),
    .A2(_04596_),
    .A3(_04597_),
    .B1(net234),
    .X(_04600_));
 sky130_fd_sc_hd__o21a_1 _11678_ (.A1(_04485_),
    .A2(_04486_),
    .B1(_04484_),
    .X(_04601_));
 sky130_fd_sc_hd__nor2_1 _11679_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04602_));
 sky130_fd_sc_hd__nand2_1 _11680_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04603_));
 sky130_fd_sc_hd__and2b_1 _11681_ (.A_N(_04602_),
    .B(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__xnor2_1 _11682_ (.A(_04601_),
    .B(_04604_),
    .Y(_04605_));
 sky130_fd_sc_hd__or2_1 _11683_ (.A(net244),
    .B(_04506_),
    .X(_04606_));
 sky130_fd_sc_hd__o211a_1 _11684_ (.A1(net224),
    .A2(_04605_),
    .B1(_04606_),
    .C1(net205),
    .X(_04607_));
 sky130_fd_sc_hd__o21a_1 _11685_ (.A1(\div_shifter[47] ),
    .A2(_04493_),
    .B1(net227),
    .X(_04608_));
 sky130_fd_sc_hd__o21ai_1 _11686_ (.A1(\div_shifter[48] ),
    .A2(_04608_),
    .B1(_02441_),
    .Y(_04610_));
 sky130_fd_sc_hd__a21oi_1 _11687_ (.A1(\div_shifter[48] ),
    .A2(_04608_),
    .B1(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nor2_1 _11688_ (.A(reg1_val[16]),
    .B(net232),
    .Y(_04612_));
 sky130_fd_sc_hd__a221o_1 _11689_ (.A1(_06147_),
    .A2(_02435_),
    .B1(net193),
    .B2(_06135_),
    .C1(_04612_),
    .X(_04613_));
 sky130_fd_sc_hd__a221o_1 _11690_ (.A1(_06153_),
    .A2(net196),
    .B1(net257),
    .B2(_00382_),
    .C1(_04613_),
    .X(_04614_));
 sky130_fd_sc_hd__or2_1 _11691_ (.A(\div_res[15] ),
    .B(_04496_),
    .X(_04615_));
 sky130_fd_sc_hd__a21oi_1 _11692_ (.A1(net139),
    .A2(_04615_),
    .B1(\div_res[16] ),
    .Y(_04616_));
 sky130_fd_sc_hd__a31o_1 _11693_ (.A1(\div_res[16] ),
    .A2(net139),
    .A3(_04615_),
    .B1(net189),
    .X(_04617_));
 sky130_fd_sc_hd__o22a_1 _11694_ (.A1(_02425_),
    .A2(_04507_),
    .B1(_04616_),
    .B2(_04617_),
    .X(_04618_));
 sky130_fd_sc_hd__o21ai_1 _11695_ (.A1(net168),
    .A2(_04491_),
    .B1(_04618_),
    .Y(_04619_));
 sky130_fd_sc_hd__or4_2 _11696_ (.A(_04607_),
    .B(_04611_),
    .C(_04614_),
    .D(_04619_),
    .X(_04621_));
 sky130_fd_sc_hd__a21oi_1 _11697_ (.A1(_04599_),
    .A2(_04600_),
    .B1(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__o221a_1 _11698_ (.A1(_04591_),
    .A2(_04592_),
    .B1(_04594_),
    .B2(_02434_),
    .C1(_04622_),
    .X(_04623_));
 sky130_fd_sc_hd__o22a_1 _11699_ (.A1(_06112_),
    .A2(net203),
    .B1(_06679_),
    .B2(_04623_),
    .X(_04624_));
 sky130_fd_sc_hd__or2_1 _11700_ (.A(curr_PC[16]),
    .B(_04513_),
    .X(_04625_));
 sky130_fd_sc_hd__a21oi_1 _11701_ (.A1(curr_PC[16]),
    .A2(_04513_),
    .B1(net237),
    .Y(_04626_));
 sky130_fd_sc_hd__a2bb2o_4 _11702_ (.A1_N(net243),
    .A2_N(_04624_),
    .B1(_04625_),
    .B2(_04626_),
    .X(dest_val[16]));
 sky130_fd_sc_hd__o21a_1 _11703_ (.A1(_04516_),
    .A2(_04590_),
    .B1(net138),
    .X(_04627_));
 sky130_fd_sc_hd__o22a_1 _11704_ (.A1(net29),
    .A2(_02066_),
    .B1(_02176_),
    .B2(net27),
    .X(_04628_));
 sky130_fd_sc_hd__xnor2_1 _11705_ (.A(net89),
    .B(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__o22a_1 _11706_ (.A1(net20),
    .A2(_00517_),
    .B1(_00811_),
    .B2(net18),
    .X(_04631_));
 sky130_fd_sc_hd__xnor2_1 _11707_ (.A(net97),
    .B(_04631_),
    .Y(_04632_));
 sky130_fd_sc_hd__nand2_1 _11708_ (.A(_00359_),
    .B(_04632_),
    .Y(_04633_));
 sky130_fd_sc_hd__xnor2_1 _11709_ (.A(net87),
    .B(_04632_),
    .Y(_04634_));
 sky130_fd_sc_hd__xnor2_1 _11710_ (.A(_04629_),
    .B(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__or2_1 _11711_ (.A(_04533_),
    .B(_04635_),
    .X(_04636_));
 sky130_fd_sc_hd__xor2_1 _11712_ (.A(_04533_),
    .B(_04635_),
    .X(_04637_));
 sky130_fd_sc_hd__nand2b_1 _11713_ (.A_N(_04522_),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__xnor2_1 _11714_ (.A(_04522_),
    .B(_04637_),
    .Y(_04639_));
 sky130_fd_sc_hd__a22o_1 _11715_ (.A1(_00161_),
    .A2(net15),
    .B1(net31),
    .B2(_00144_),
    .X(_04640_));
 sky130_fd_sc_hd__xnor2_1 _11716_ (.A(net91),
    .B(_04640_),
    .Y(_04642_));
 sky130_fd_sc_hd__inv_2 _11717_ (.A(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__o22a_1 _11718_ (.A1(net54),
    .A2(net34),
    .B1(net32),
    .B2(net48),
    .X(_04644_));
 sky130_fd_sc_hd__xnor2_1 _11719_ (.A(net94),
    .B(_04644_),
    .Y(_04645_));
 sky130_fd_sc_hd__o22a_1 _11720_ (.A1(net52),
    .A2(net38),
    .B1(net36),
    .B2(net43),
    .X(_04646_));
 sky130_fd_sc_hd__xnor2_1 _11721_ (.A(net98),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__xnor2_1 _11722_ (.A(_04645_),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__nor2_1 _11723_ (.A(_04643_),
    .B(_04648_),
    .Y(_04649_));
 sky130_fd_sc_hd__and2_1 _11724_ (.A(_04643_),
    .B(_04648_),
    .X(_04650_));
 sky130_fd_sc_hd__nor2_1 _11725_ (.A(_04649_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__nand2_1 _11726_ (.A(_04639_),
    .B(_04651_),
    .Y(_04653_));
 sky130_fd_sc_hd__or2_1 _11727_ (.A(_04639_),
    .B(_04651_),
    .X(_04654_));
 sky130_fd_sc_hd__a22o_1 _11728_ (.A1(_00203_),
    .A2(net8),
    .B1(net3),
    .B2(net101),
    .X(_04655_));
 sky130_fd_sc_hd__xnor2_1 _11729_ (.A(net62),
    .B(_04655_),
    .Y(_04656_));
 sky130_fd_sc_hd__a22o_1 _11730_ (.A1(_06725_),
    .A2(net17),
    .B1(net12),
    .B2(_00208_),
    .X(_04657_));
 sky130_fd_sc_hd__xnor2_1 _11731_ (.A(net65),
    .B(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__nor2_1 _11732_ (.A(net103),
    .B(net59),
    .Y(_04659_));
 sky130_fd_sc_hd__xnor2_1 _11733_ (.A(_04658_),
    .B(_04659_),
    .Y(_04660_));
 sky130_fd_sc_hd__nor2_1 _11734_ (.A(_04656_),
    .B(_04660_),
    .Y(_04661_));
 sky130_fd_sc_hd__and2_1 _11735_ (.A(_04656_),
    .B(_04660_),
    .X(_04662_));
 sky130_fd_sc_hd__nor2_1 _11736_ (.A(_04661_),
    .B(_04662_),
    .Y(_04663_));
 sky130_fd_sc_hd__and3_1 _11737_ (.A(_04653_),
    .B(_04654_),
    .C(_04663_),
    .X(_04664_));
 sky130_fd_sc_hd__a21oi_1 _11738_ (.A1(_04653_),
    .A2(_04654_),
    .B1(_04663_),
    .Y(_04665_));
 sky130_fd_sc_hd__nor2_1 _11739_ (.A(_04664_),
    .B(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__o21ba_1 _11740_ (.A1(_04536_),
    .A2(_04550_),
    .B1_N(_04560_),
    .X(_04667_));
 sky130_fd_sc_hd__a21o_1 _11741_ (.A1(_04552_),
    .A2(_04555_),
    .B1(_04557_),
    .X(_04668_));
 sky130_fd_sc_hd__o21bai_1 _11742_ (.A1(_04527_),
    .A2(_04535_),
    .B1_N(_04525_),
    .Y(_04669_));
 sky130_fd_sc_hd__nor2_1 _11743_ (.A(_04545_),
    .B(_04548_),
    .Y(_04670_));
 sky130_fd_sc_hd__o21a_1 _11744_ (.A1(_04545_),
    .A2(_04548_),
    .B1(_04669_),
    .X(_04671_));
 sky130_fd_sc_hd__xnor2_1 _11745_ (.A(_04669_),
    .B(_04670_),
    .Y(_04672_));
 sky130_fd_sc_hd__xnor2_1 _11746_ (.A(_04668_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__a21bo_1 _11747_ (.A1(_04563_),
    .A2(_04566_),
    .B1_N(_04564_),
    .X(_04674_));
 sky130_fd_sc_hd__nand2b_1 _11748_ (.A_N(_04673_),
    .B(_04674_),
    .Y(_04675_));
 sky130_fd_sc_hd__xnor2_1 _11749_ (.A(_04673_),
    .B(_04674_),
    .Y(_04676_));
 sky130_fd_sc_hd__nand2b_1 _11750_ (.A_N(_04667_),
    .B(_04676_),
    .Y(_04677_));
 sky130_fd_sc_hd__xnor2_1 _11751_ (.A(_04667_),
    .B(_04676_),
    .Y(_04678_));
 sky130_fd_sc_hd__nand2_1 _11752_ (.A(_04666_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__xnor2_1 _11753_ (.A(_04666_),
    .B(_04678_),
    .Y(_04680_));
 sky130_fd_sc_hd__o21ai_2 _11754_ (.A1(_04568_),
    .A2(_04569_),
    .B1(_04571_),
    .Y(_04681_));
 sky130_fd_sc_hd__nand2b_1 _11755_ (.A_N(_04680_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__xor2_1 _11756_ (.A(_04680_),
    .B(_04681_),
    .X(_04683_));
 sky130_fd_sc_hd__a21oi_1 _11757_ (.A1(_04573_),
    .A2(_04577_),
    .B1(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__nand3_1 _11758_ (.A(_04573_),
    .B(_04577_),
    .C(_04683_),
    .Y(_04685_));
 sky130_fd_sc_hd__nand2b_2 _11759_ (.A_N(_04684_),
    .B(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__o21a_1 _11760_ (.A1(_04461_),
    .A2(_04580_),
    .B1(_04581_),
    .X(_04687_));
 sky130_fd_sc_hd__nor2_1 _11761_ (.A(_04463_),
    .B(_04582_),
    .Y(_04688_));
 sky130_fd_sc_hd__a21o_1 _11762_ (.A1(_04464_),
    .A2(_04688_),
    .B1(_04687_),
    .X(_04689_));
 sky130_fd_sc_hd__nand2_1 _11763_ (.A(_04465_),
    .B(_04688_),
    .Y(_04690_));
 sky130_fd_sc_hd__a31oi_2 _11764_ (.A1(_04252_),
    .A2(_04465_),
    .A3(_04688_),
    .B1(_04689_),
    .Y(_04691_));
 sky130_fd_sc_hd__o31ai_4 _11765_ (.A1(_03770_),
    .A2(_04250_),
    .A3(_04690_),
    .B1(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__xnor2_4 _11766_ (.A(_04686_),
    .B(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__o21ai_1 _11767_ (.A1(_04627_),
    .A2(_04693_),
    .B1(_02348_),
    .Y(_04694_));
 sky130_fd_sc_hd__a21oi_1 _11768_ (.A1(_04627_),
    .A2(_04693_),
    .B1(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__o21ai_1 _11769_ (.A1(net135),
    .A2(_01968_),
    .B1(_01969_),
    .Y(_04696_));
 sky130_fd_sc_hd__o31a_1 _11770_ (.A1(net134),
    .A2(_01968_),
    .A3(_01969_),
    .B1(net233),
    .X(_04697_));
 sky130_fd_sc_hd__a21o_1 _11771_ (.A1(_06135_),
    .A2(_04595_),
    .B1(_06147_),
    .X(_04698_));
 sky130_fd_sc_hd__and3_1 _11772_ (.A(net294),
    .B(_06129_),
    .C(_06594_),
    .X(_04699_));
 sky130_fd_sc_hd__a21oi_1 _11773_ (.A1(net283),
    .A2(_04698_),
    .B1(_04699_),
    .Y(_04700_));
 sky130_fd_sc_hd__xnor2_2 _11774_ (.A(_06076_),
    .B(_04700_),
    .Y(_04701_));
 sky130_fd_sc_hd__o21a_1 _11775_ (.A1(_04601_),
    .A2(_04602_),
    .B1(_04603_),
    .X(_04702_));
 sky130_fd_sc_hd__nor2_1 _11776_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04703_));
 sky130_fd_sc_hd__nand2_1 _11777_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04704_));
 sky130_fd_sc_hd__nand2b_1 _11778_ (.A_N(_04703_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__xor2_1 _11779_ (.A(_04702_),
    .B(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(_04390_),
    .A1(_04706_),
    .S(net244),
    .X(_04707_));
 sky130_fd_sc_hd__o22ai_1 _11781_ (.A1(_06068_),
    .A2(_02436_),
    .B1(_02445_),
    .B2(reg1_val[17]),
    .Y(_04708_));
 sky130_fd_sc_hd__a221o_1 _11782_ (.A1(_06076_),
    .A2(net195),
    .B1(net193),
    .B2(_06059_),
    .C1(_04708_),
    .X(_04709_));
 sky130_fd_sc_hd__a31o_1 _11783_ (.A1(_00355_),
    .A2(_00356_),
    .A3(net256),
    .B1(_04709_),
    .X(_04710_));
 sky130_fd_sc_hd__a221o_1 _11784_ (.A1(net171),
    .A2(_04379_),
    .B1(_04390_),
    .B2(net167),
    .C1(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__o31a_1 _11785_ (.A1(\div_shifter[48] ),
    .A2(\div_shifter[47] ),
    .A3(_04493_),
    .B1(net227),
    .X(_04712_));
 sky130_fd_sc_hd__xor2_1 _11786_ (.A(\div_shifter[49] ),
    .B(_04712_),
    .X(_04713_));
 sky130_fd_sc_hd__o21ai_1 _11787_ (.A1(\div_res[16] ),
    .A2(_04615_),
    .B1(net141),
    .Y(_04714_));
 sky130_fd_sc_hd__xnor2_1 _11788_ (.A(\div_res[17] ),
    .B(_04714_),
    .Y(_04715_));
 sky130_fd_sc_hd__a22o_1 _11789_ (.A1(_02441_),
    .A2(_04713_),
    .B1(_04715_),
    .B2(_02443_),
    .X(_04716_));
 sky130_fd_sc_hd__a211o_1 _11790_ (.A1(net205),
    .A2(_04707_),
    .B1(_04711_),
    .C1(_04716_),
    .X(_04717_));
 sky130_fd_sc_hd__a221o_1 _11791_ (.A1(_04696_),
    .A2(_04697_),
    .B1(_04701_),
    .B2(net234),
    .C1(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__o21ba_1 _11792_ (.A1(_04695_),
    .A2(_04718_),
    .B1_N(_06679_),
    .X(_04719_));
 sky130_fd_sc_hd__nor2_1 _11793_ (.A(_06031_),
    .B(net203),
    .Y(_04720_));
 sky130_fd_sc_hd__and3_1 _11794_ (.A(curr_PC[16]),
    .B(curr_PC[17]),
    .C(_04513_),
    .X(_04721_));
 sky130_fd_sc_hd__a21oi_1 _11795_ (.A1(curr_PC[16]),
    .A2(_04513_),
    .B1(curr_PC[17]),
    .Y(_04722_));
 sky130_fd_sc_hd__o21ai_1 _11796_ (.A1(_04721_),
    .A2(_04722_),
    .B1(net242),
    .Y(_04724_));
 sky130_fd_sc_hd__o31a_4 _11797_ (.A1(net243),
    .A2(_04719_),
    .A3(_04720_),
    .B1(_04724_),
    .X(dest_val[17]));
 sky130_fd_sc_hd__or2_1 _11798_ (.A(_04590_),
    .B(_04693_),
    .X(_04725_));
 sky130_fd_sc_hd__o21a_1 _11799_ (.A1(_04516_),
    .A2(_04725_),
    .B1(net138),
    .X(_04726_));
 sky130_fd_sc_hd__or2_1 _11800_ (.A(_00364_),
    .B(net5),
    .X(_04727_));
 sky130_fd_sc_hd__a22o_2 _11801_ (.A1(_00366_),
    .A2(net7),
    .B1(_04727_),
    .B2(net89),
    .X(_04728_));
 sky130_fd_sc_hd__nand2_1 _11802_ (.A(net101),
    .B(net62),
    .Y(_04729_));
 sky130_fd_sc_hd__and2_1 _11803_ (.A(_04728_),
    .B(_04729_),
    .X(_04730_));
 sky130_fd_sc_hd__nor2_1 _11804_ (.A(_04728_),
    .B(_04729_),
    .Y(_04731_));
 sky130_fd_sc_hd__nor2_1 _11805_ (.A(_04730_),
    .B(_04731_),
    .Y(_04732_));
 sky130_fd_sc_hd__a21bo_1 _11806_ (.A1(_04629_),
    .A2(_04634_),
    .B1_N(_04633_),
    .X(_04733_));
 sky130_fd_sc_hd__xnor2_1 _11807_ (.A(_04732_),
    .B(_04733_),
    .Y(_04734_));
 sky130_fd_sc_hd__o22a_1 _11808_ (.A1(net43),
    .A2(net38),
    .B1(net36),
    .B2(_00517_),
    .X(_04735_));
 sky130_fd_sc_hd__xnor2_1 _11809_ (.A(net98),
    .B(_04735_),
    .Y(_04736_));
 sky130_fd_sc_hd__inv_2 _11810_ (.A(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__o22a_1 _11811_ (.A1(net20),
    .A2(_00811_),
    .B1(net10),
    .B2(net18),
    .X(_04738_));
 sky130_fd_sc_hd__xnor2_1 _11812_ (.A(net97),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__a22o_1 _11813_ (.A1(_00144_),
    .A2(net15),
    .B1(net31),
    .B2(_00136_),
    .X(_04740_));
 sky130_fd_sc_hd__xnor2_1 _11814_ (.A(net91),
    .B(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__and2_1 _11815_ (.A(_04739_),
    .B(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__nor2_1 _11816_ (.A(_04739_),
    .B(_04741_),
    .Y(_04743_));
 sky130_fd_sc_hd__or2_1 _11817_ (.A(_04742_),
    .B(_04743_),
    .X(_04744_));
 sky130_fd_sc_hd__nor2_1 _11818_ (.A(_04737_),
    .B(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__and2_1 _11819_ (.A(_04737_),
    .B(_04744_),
    .X(_04746_));
 sky130_fd_sc_hd__or2_1 _11820_ (.A(_04745_),
    .B(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__xnor2_1 _11821_ (.A(_04734_),
    .B(_04747_),
    .Y(_04748_));
 sky130_fd_sc_hd__a22o_1 _11822_ (.A1(net55),
    .A2(net17),
    .B1(net12),
    .B2(_06725_),
    .X(_04749_));
 sky130_fd_sc_hd__xnor2_1 _11823_ (.A(_00787_),
    .B(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__a22o_1 _11824_ (.A1(_00208_),
    .A2(net8),
    .B1(net3),
    .B2(_00203_),
    .X(_04751_));
 sky130_fd_sc_hd__xnor2_1 _11825_ (.A(net59),
    .B(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__o22a_1 _11826_ (.A1(net48),
    .A2(net34),
    .B1(net32),
    .B2(net46),
    .X(_04754_));
 sky130_fd_sc_hd__xnor2_1 _11827_ (.A(net93),
    .B(_04754_),
    .Y(_04755_));
 sky130_fd_sc_hd__nand2_1 _11828_ (.A(_04752_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__xnor2_1 _11829_ (.A(_04752_),
    .B(_04755_),
    .Y(_04757_));
 sky130_fd_sc_hd__xnor2_1 _11830_ (.A(_04750_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__or2_1 _11831_ (.A(_04748_),
    .B(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__nand2_1 _11832_ (.A(_04748_),
    .B(_04758_),
    .Y(_04760_));
 sky130_fd_sc_hd__and2_1 _11833_ (.A(_04759_),
    .B(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__a21o_1 _11834_ (.A1(_04639_),
    .A2(_04651_),
    .B1(_04664_),
    .X(_04762_));
 sky130_fd_sc_hd__a21o_1 _11835_ (.A1(_04658_),
    .A2(_04659_),
    .B1(_04661_),
    .X(_04763_));
 sky130_fd_sc_hd__a21oi_1 _11836_ (.A1(_04645_),
    .A2(_04647_),
    .B1(_04649_),
    .Y(_04765_));
 sky130_fd_sc_hd__a21o_1 _11837_ (.A1(_04636_),
    .A2(_04638_),
    .B1(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__nand3_1 _11838_ (.A(_04636_),
    .B(_04638_),
    .C(_04765_),
    .Y(_04767_));
 sky130_fd_sc_hd__and2_1 _11839_ (.A(_04766_),
    .B(_04767_),
    .X(_04768_));
 sky130_fd_sc_hd__nand2_1 _11840_ (.A(_04763_),
    .B(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__xnor2_1 _11841_ (.A(_04763_),
    .B(_04768_),
    .Y(_04770_));
 sky130_fd_sc_hd__a21oi_2 _11842_ (.A1(_04668_),
    .A2(_04672_),
    .B1(_04671_),
    .Y(_04771_));
 sky130_fd_sc_hd__xnor2_1 _11843_ (.A(_04770_),
    .B(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__and2b_1 _11844_ (.A_N(_04772_),
    .B(_04762_),
    .X(_04773_));
 sky130_fd_sc_hd__xnor2_1 _11845_ (.A(_04762_),
    .B(_04772_),
    .Y(_04774_));
 sky130_fd_sc_hd__nand2_1 _11846_ (.A(_04761_),
    .B(_04774_),
    .Y(_04776_));
 sky130_fd_sc_hd__or2_1 _11847_ (.A(_04761_),
    .B(_04774_),
    .X(_04777_));
 sky130_fd_sc_hd__nand2_1 _11848_ (.A(_04776_),
    .B(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__nand2_1 _11849_ (.A(_04675_),
    .B(_04677_),
    .Y(_04779_));
 sky130_fd_sc_hd__nand2b_1 _11850_ (.A_N(_04778_),
    .B(_04779_),
    .Y(_04780_));
 sky130_fd_sc_hd__xor2_2 _11851_ (.A(_04778_),
    .B(_04779_),
    .X(_04781_));
 sky130_fd_sc_hd__a21oi_2 _11852_ (.A1(_04679_),
    .A2(_04682_),
    .B1(_04781_),
    .Y(_04782_));
 sky130_fd_sc_hd__nand3_2 _11853_ (.A(_04679_),
    .B(_04682_),
    .C(_04781_),
    .Y(_04783_));
 sky130_fd_sc_hd__nand2b_4 _11854_ (.A_N(_04782_),
    .B(_04783_),
    .Y(_04784_));
 sky130_fd_sc_hd__o21a_1 _11855_ (.A1(_04580_),
    .A2(_04684_),
    .B1(_04685_),
    .X(_04785_));
 sky130_fd_sc_hd__nor2_1 _11856_ (.A(_04582_),
    .B(_04686_),
    .Y(_04787_));
 sky130_fd_sc_hd__and2_1 _11857_ (.A(_04584_),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__inv_2 _11858_ (.A(_04788_),
    .Y(_04789_));
 sky130_fd_sc_hd__a221oi_1 _11859_ (.A1(_04583_),
    .A2(_04787_),
    .B1(_04788_),
    .B2(_04359_),
    .C1(_04785_),
    .Y(_04790_));
 sky130_fd_sc_hd__o31a_2 _11860_ (.A1(_03893_),
    .A2(_04360_),
    .A3(_04789_),
    .B1(_04790_),
    .X(_04791_));
 sky130_fd_sc_hd__xor2_4 _11861_ (.A(_04784_),
    .B(_04791_),
    .X(_04792_));
 sky130_fd_sc_hd__nor2_1 _11862_ (.A(_04726_),
    .B(_04792_),
    .Y(_04793_));
 sky130_fd_sc_hd__a21o_1 _11863_ (.A1(_04726_),
    .A2(_04792_),
    .B1(net235),
    .X(_04794_));
 sky130_fd_sc_hd__and4_1 _11864_ (.A(net136),
    .B(_01970_),
    .C(_01974_),
    .D(_01975_),
    .X(_04795_));
 sky130_fd_sc_hd__a22o_1 _11865_ (.A1(net136),
    .A2(_01970_),
    .B1(_01974_),
    .B2(_01975_),
    .X(_04796_));
 sky130_fd_sc_hd__nand2_1 _11866_ (.A(net233),
    .B(_04796_),
    .Y(_04798_));
 sky130_fd_sc_hd__and3_1 _11867_ (.A(net294),
    .B(_06050_),
    .C(_06595_),
    .X(_04799_));
 sky130_fd_sc_hd__a21bo_1 _11868_ (.A1(_06059_),
    .A2(_04698_),
    .B1_N(_06068_),
    .X(_04800_));
 sky130_fd_sc_hd__a21o_1 _11869_ (.A1(net284),
    .A2(_04800_),
    .B1(_04799_),
    .X(_04801_));
 sky130_fd_sc_hd__o21ai_1 _11870_ (.A1(_05995_),
    .A2(_04801_),
    .B1(net234),
    .Y(_04802_));
 sky130_fd_sc_hd__a21o_1 _11871_ (.A1(_05995_),
    .A2(_04801_),
    .B1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__or2_1 _11872_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .X(_04804_));
 sky130_fd_sc_hd__nand2_1 _11873_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .Y(_04805_));
 sky130_fd_sc_hd__nand2_1 _11874_ (.A(_04804_),
    .B(_04805_),
    .Y(_04806_));
 sky130_fd_sc_hd__o21ai_1 _11875_ (.A1(_04702_),
    .A2(_04703_),
    .B1(_04704_),
    .Y(_04807_));
 sky130_fd_sc_hd__xor2_1 _11876_ (.A(_04806_),
    .B(_04807_),
    .X(_04809_));
 sky130_fd_sc_hd__mux2_1 _11877_ (.A0(_04284_),
    .A1(_04809_),
    .S(net244),
    .X(_04810_));
 sky130_fd_sc_hd__or3_1 _11878_ (.A(\div_res[17] ),
    .B(\div_res[16] ),
    .C(_04615_),
    .X(_04811_));
 sky130_fd_sc_hd__a21oi_1 _11879_ (.A1(net141),
    .A2(_04811_),
    .B1(\div_res[18] ),
    .Y(_04812_));
 sky130_fd_sc_hd__a311o_1 _11880_ (.A1(\div_res[18] ),
    .A2(net141),
    .A3(_04811_),
    .B1(_04812_),
    .C1(net189),
    .X(_04813_));
 sky130_fd_sc_hd__or4_1 _11881_ (.A(\div_shifter[49] ),
    .B(\div_shifter[48] ),
    .C(\div_shifter[47] ),
    .D(_04493_),
    .X(_04814_));
 sky130_fd_sc_hd__a21oi_1 _11882_ (.A1(net227),
    .A2(_04814_),
    .B1(\div_shifter[50] ),
    .Y(_04815_));
 sky130_fd_sc_hd__a311o_1 _11883_ (.A1(\div_shifter[50] ),
    .A2(net227),
    .A3(_04814_),
    .B1(_04815_),
    .C1(net191),
    .X(_04816_));
 sky130_fd_sc_hd__and3_1 _11884_ (.A(_00350_),
    .B(_00360_),
    .C(net256),
    .X(_04817_));
 sky130_fd_sc_hd__a2bb2o_1 _11885_ (.A1_N(reg1_val[18]),
    .A2_N(net232),
    .B1(_05949_),
    .B2(_06677_),
    .X(_04818_));
 sky130_fd_sc_hd__a221o_1 _11886_ (.A1(_05986_),
    .A2(_02435_),
    .B1(net193),
    .B2(_05978_),
    .C1(_04818_),
    .X(_04820_));
 sky130_fd_sc_hd__a211o_1 _11887_ (.A1(_05995_),
    .A2(net196),
    .B1(_04817_),
    .C1(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__o2bb2a_1 _11888_ (.A1_N(net171),
    .A2_N(_04271_),
    .B1(_04284_),
    .B2(_02425_),
    .X(_04822_));
 sky130_fd_sc_hd__and4b_1 _11889_ (.A_N(_04821_),
    .B(_04822_),
    .C(_04813_),
    .D(_04816_),
    .X(_04823_));
 sky130_fd_sc_hd__o211a_1 _11890_ (.A1(_06667_),
    .A2(_04810_),
    .B1(_04823_),
    .C1(_04803_),
    .X(_04824_));
 sky130_fd_sc_hd__o221a_1 _11891_ (.A1(_04793_),
    .A2(_04794_),
    .B1(_04795_),
    .B2(_04798_),
    .C1(_04824_),
    .X(_04825_));
 sky130_fd_sc_hd__nor2_1 _11892_ (.A(curr_PC[18]),
    .B(_04721_),
    .Y(_04826_));
 sky130_fd_sc_hd__and2_1 _11893_ (.A(curr_PC[18]),
    .B(_04721_),
    .X(_04827_));
 sky130_fd_sc_hd__or3_1 _11894_ (.A(net241),
    .B(_04826_),
    .C(_04827_),
    .X(_04828_));
 sky130_fd_sc_hd__o21ai_4 _11895_ (.A1(net242),
    .A2(_04825_),
    .B1(_04828_),
    .Y(dest_val[18]));
 sky130_fd_sc_hd__or4_2 _11896_ (.A(_04059_),
    .B(_04515_),
    .C(_04725_),
    .D(_04792_),
    .X(_04830_));
 sky130_fd_sc_hd__o21bai_2 _11897_ (.A1(_04770_),
    .A2(_04771_),
    .B1_N(_04773_),
    .Y(_04831_));
 sky130_fd_sc_hd__o22a_1 _11898_ (.A1(net46),
    .A2(net34),
    .B1(net32),
    .B2(net50),
    .X(_04832_));
 sky130_fd_sc_hd__xnor2_2 _11899_ (.A(net93),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__a22o_1 _11900_ (.A1(_00150_),
    .A2(_00562_),
    .B1(net13),
    .B2(net55),
    .X(_04834_));
 sky130_fd_sc_hd__xnor2_1 _11901_ (.A(net64),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__o22a_1 _11902_ (.A1(net52),
    .A2(_00336_),
    .B1(_00342_),
    .B2(net43),
    .X(_04836_));
 sky130_fd_sc_hd__xnor2_1 _11903_ (.A(net92),
    .B(_04836_),
    .Y(_04837_));
 sky130_fd_sc_hd__nand2_1 _11904_ (.A(_04835_),
    .B(_04837_),
    .Y(_04838_));
 sky130_fd_sc_hd__or2_1 _11905_ (.A(_04835_),
    .B(_04837_),
    .X(_04839_));
 sky130_fd_sc_hd__nand2_1 _11906_ (.A(_04838_),
    .B(_04839_),
    .Y(_04841_));
 sky130_fd_sc_hd__xnor2_2 _11907_ (.A(_04833_),
    .B(_04841_),
    .Y(_04842_));
 sky130_fd_sc_hd__o22a_1 _11908_ (.A1(net20),
    .A2(net10),
    .B1(net5),
    .B2(net18),
    .X(_04843_));
 sky130_fd_sc_hd__xnor2_1 _11909_ (.A(_00274_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__o22a_1 _11910_ (.A1(net38),
    .A2(_00517_),
    .B1(_00811_),
    .B2(net37),
    .X(_04845_));
 sky130_fd_sc_hd__xnor2_1 _11911_ (.A(net98),
    .B(_04845_),
    .Y(_04846_));
 sky130_fd_sc_hd__nand2b_1 _11912_ (.A_N(net89),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__xor2_1 _11913_ (.A(net89),
    .B(_04846_),
    .X(_04848_));
 sky130_fd_sc_hd__or2_1 _11914_ (.A(_04844_),
    .B(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__nand2_1 _11915_ (.A(_04844_),
    .B(_04848_),
    .Y(_04850_));
 sky130_fd_sc_hd__nand2_1 _11916_ (.A(_04849_),
    .B(_04850_),
    .Y(_04852_));
 sky130_fd_sc_hd__a22o_1 _11917_ (.A1(_06725_),
    .A2(net8),
    .B1(net3),
    .B2(_00208_),
    .X(_04853_));
 sky130_fd_sc_hd__xnor2_1 _11918_ (.A(net58),
    .B(_04853_),
    .Y(_04854_));
 sky130_fd_sc_hd__nand2_1 _11919_ (.A(_04728_),
    .B(_04854_),
    .Y(_04855_));
 sky130_fd_sc_hd__or2_1 _11920_ (.A(_04728_),
    .B(_04854_),
    .X(_04856_));
 sky130_fd_sc_hd__nand2_1 _11921_ (.A(_04855_),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__nand2_1 _11922_ (.A(_00203_),
    .B(net61),
    .Y(_04858_));
 sky130_fd_sc_hd__xor2_2 _11923_ (.A(_04857_),
    .B(_04858_),
    .X(_04859_));
 sky130_fd_sc_hd__xnor2_2 _11924_ (.A(_04852_),
    .B(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__xor2_2 _11925_ (.A(_04842_),
    .B(_04860_),
    .X(_04861_));
 sky130_fd_sc_hd__o21a_1 _11926_ (.A1(_04734_),
    .A2(_04747_),
    .B1(_04759_),
    .X(_04863_));
 sky130_fd_sc_hd__o21ai_1 _11927_ (.A1(_04750_),
    .A2(_04757_),
    .B1(_04756_),
    .Y(_04864_));
 sky130_fd_sc_hd__a21o_1 _11928_ (.A1(_04732_),
    .A2(_04733_),
    .B1(_04731_),
    .X(_04865_));
 sky130_fd_sc_hd__nor2_1 _11929_ (.A(_04742_),
    .B(_04745_),
    .Y(_04866_));
 sky130_fd_sc_hd__o21ai_1 _11930_ (.A1(_04742_),
    .A2(_04745_),
    .B1(_04865_),
    .Y(_04867_));
 sky130_fd_sc_hd__xnor2_1 _11931_ (.A(_04865_),
    .B(_04866_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand2_1 _11932_ (.A(_04864_),
    .B(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__xnor2_1 _11933_ (.A(_04864_),
    .B(_04868_),
    .Y(_04870_));
 sky130_fd_sc_hd__a21oi_1 _11934_ (.A1(_04766_),
    .A2(_04769_),
    .B1(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__and3_1 _11935_ (.A(_04766_),
    .B(_04769_),
    .C(_04870_),
    .X(_04872_));
 sky130_fd_sc_hd__nor2_1 _11936_ (.A(_04871_),
    .B(_04872_),
    .Y(_04874_));
 sky130_fd_sc_hd__and2b_1 _11937_ (.A_N(_04863_),
    .B(_04874_),
    .X(_04875_));
 sky130_fd_sc_hd__xnor2_2 _11938_ (.A(_04863_),
    .B(_04874_),
    .Y(_04876_));
 sky130_fd_sc_hd__and2_1 _11939_ (.A(_04861_),
    .B(_04876_),
    .X(_04877_));
 sky130_fd_sc_hd__xor2_2 _11940_ (.A(_04861_),
    .B(_04876_),
    .X(_04878_));
 sky130_fd_sc_hd__and2_1 _11941_ (.A(_04831_),
    .B(_04878_),
    .X(_04879_));
 sky130_fd_sc_hd__xnor2_2 _11942_ (.A(_04831_),
    .B(_04878_),
    .Y(_04880_));
 sky130_fd_sc_hd__a21oi_2 _11943_ (.A1(_04776_),
    .A2(_04780_),
    .B1(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__nand3_2 _11944_ (.A(_04776_),
    .B(_04780_),
    .C(_04880_),
    .Y(_04882_));
 sky130_fd_sc_hd__nand2b_4 _11945_ (.A_N(_04881_),
    .B(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__o21a_1 _11946_ (.A1(_04684_),
    .A2(_04782_),
    .B1(_04783_),
    .X(_04885_));
 sky130_fd_sc_hd__inv_2 _11947_ (.A(_04885_),
    .Y(_04886_));
 sky130_fd_sc_hd__nor2_1 _11948_ (.A(_04686_),
    .B(_04784_),
    .Y(_04887_));
 sky130_fd_sc_hd__a21oi_1 _11949_ (.A1(_04687_),
    .A2(_04887_),
    .B1(_04885_),
    .Y(_04888_));
 sky130_fd_sc_hd__and2_1 _11950_ (.A(_04688_),
    .B(_04887_),
    .X(_04889_));
 sky130_fd_sc_hd__a21bo_1 _11951_ (.A1(_04470_),
    .A2(_04889_),
    .B1_N(_04888_),
    .X(_04890_));
 sky130_fd_sc_hd__xnor2_4 _11952_ (.A(_04883_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__a21oi_1 _11953_ (.A1(net138),
    .A2(_04830_),
    .B1(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__and3_1 _11954_ (.A(net138),
    .B(_04830_),
    .C(_04891_),
    .X(_04893_));
 sky130_fd_sc_hd__or3_1 _11955_ (.A(net235),
    .B(_04892_),
    .C(_04893_),
    .X(_04894_));
 sky130_fd_sc_hd__o21a_1 _11956_ (.A1(net135),
    .A2(_01976_),
    .B1(_01977_),
    .X(_04896_));
 sky130_fd_sc_hd__nor3_1 _11957_ (.A(net135),
    .B(_01976_),
    .C(_01977_),
    .Y(_04897_));
 sky130_fd_sc_hd__and3_1 _11958_ (.A(net294),
    .B(_05959_),
    .C(_06596_),
    .X(_04898_));
 sky130_fd_sc_hd__a21o_1 _11959_ (.A1(_05995_),
    .A2(_04800_),
    .B1(_05986_),
    .X(_04899_));
 sky130_fd_sc_hd__a21o_1 _11960_ (.A1(net283),
    .A2(_04899_),
    .B1(_04898_),
    .X(_04900_));
 sky130_fd_sc_hd__nand2_1 _11961_ (.A(_05912_),
    .B(_04900_),
    .Y(_04901_));
 sky130_fd_sc_hd__o211a_1 _11962_ (.A1(_05912_),
    .A2(_04900_),
    .B1(_04901_),
    .C1(net234),
    .X(_04902_));
 sky130_fd_sc_hd__or2_1 _11963_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .X(_04903_));
 sky130_fd_sc_hd__nand2_1 _11964_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .Y(_04904_));
 sky130_fd_sc_hd__nand2_1 _11965_ (.A(_04903_),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21boi_1 _11966_ (.A1(_04804_),
    .A2(_04807_),
    .B1_N(_04805_),
    .Y(_04907_));
 sky130_fd_sc_hd__xor2_1 _11967_ (.A(_04905_),
    .B(_04907_),
    .X(_04908_));
 sky130_fd_sc_hd__mux2_1 _11968_ (.A0(_04167_),
    .A1(_04908_),
    .S(net244),
    .X(_04909_));
 sky130_fd_sc_hd__or2_1 _11969_ (.A(\div_shifter[50] ),
    .B(_04814_),
    .X(_04910_));
 sky130_fd_sc_hd__nand3_1 _11970_ (.A(\div_shifter[51] ),
    .B(net227),
    .C(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__a21o_1 _11971_ (.A1(net227),
    .A2(_04910_),
    .B1(\div_shifter[51] ),
    .X(_04912_));
 sky130_fd_sc_hd__or2_1 _11972_ (.A(\div_res[18] ),
    .B(_04811_),
    .X(_04913_));
 sky130_fd_sc_hd__a21oi_1 _11973_ (.A1(net141),
    .A2(_04913_),
    .B1(\div_res[19] ),
    .Y(_04914_));
 sky130_fd_sc_hd__a31o_1 _11974_ (.A1(\div_res[19] ),
    .A2(net141),
    .A3(_04913_),
    .B1(net189),
    .X(_04915_));
 sky130_fd_sc_hd__nor2_1 _11975_ (.A(_04914_),
    .B(_04915_),
    .Y(_04916_));
 sky130_fd_sc_hd__a2bb2o_1 _11976_ (.A1_N(reg1_val[19]),
    .A2_N(net232),
    .B1(_02435_),
    .B2(_05902_),
    .X(_04918_));
 sky130_fd_sc_hd__a2bb2o_1 _11977_ (.A1_N(_05893_),
    .A2_N(_02440_),
    .B1(net195),
    .B2(_05912_),
    .X(_04919_));
 sky130_fd_sc_hd__a31o_1 _11978_ (.A1(_00257_),
    .A2(_00351_),
    .A3(net257),
    .B1(_04916_),
    .X(_04920_));
 sky130_fd_sc_hd__a221o_1 _11979_ (.A1(net171),
    .A2(_04149_),
    .B1(_04167_),
    .B2(net167),
    .C1(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__or3_1 _11980_ (.A(_04918_),
    .B(_04919_),
    .C(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__a31o_1 _11981_ (.A1(_02441_),
    .A2(_04911_),
    .A3(_04912_),
    .B1(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__a211oi_2 _11982_ (.A1(_06666_),
    .A2(_04909_),
    .B1(_04923_),
    .C1(_04902_),
    .Y(_04924_));
 sky130_fd_sc_hd__o311a_1 _11983_ (.A1(_02434_),
    .A2(_04896_),
    .A3(_04897_),
    .B1(_04924_),
    .C1(_04894_),
    .X(_04925_));
 sky130_fd_sc_hd__o22a_1 _11984_ (.A1(_05874_),
    .A2(net203),
    .B1(_06679_),
    .B2(_04925_),
    .X(_04926_));
 sky130_fd_sc_hd__o21ai_1 _11985_ (.A1(curr_PC[19]),
    .A2(_04827_),
    .B1(net242),
    .Y(_04927_));
 sky130_fd_sc_hd__a21o_1 _11986_ (.A1(curr_PC[19]),
    .A2(_04827_),
    .B1(_04927_),
    .X(_04929_));
 sky130_fd_sc_hd__o21ai_4 _11987_ (.A1(net242),
    .A2(_04926_),
    .B1(_04929_),
    .Y(dest_val[19]));
 sky130_fd_sc_hd__or2_1 _11988_ (.A(_04830_),
    .B(_04891_),
    .X(_04930_));
 sky130_fd_sc_hd__o22a_1 _11989_ (.A1(net38),
    .A2(_00811_),
    .B1(net10),
    .B2(net36),
    .X(_04931_));
 sky130_fd_sc_hd__xnor2_1 _11990_ (.A(net98),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__or2_1 _11991_ (.A(_00405_),
    .B(net5),
    .X(_04933_));
 sky130_fd_sc_hd__a22o_1 _11992_ (.A1(_00407_),
    .A2(net7),
    .B1(_04933_),
    .B2(net97),
    .X(_04934_));
 sky130_fd_sc_hd__nor2_1 _11993_ (.A(_04932_),
    .B(_04934_),
    .Y(_04935_));
 sky130_fd_sc_hd__and2_1 _11994_ (.A(_04932_),
    .B(_04934_),
    .X(_04936_));
 sky130_fd_sc_hd__nor2_1 _11995_ (.A(_04935_),
    .B(_04936_),
    .Y(_04937_));
 sky130_fd_sc_hd__a22o_1 _11996_ (.A1(net55),
    .A2(net8),
    .B1(net3),
    .B2(_06725_),
    .X(_04939_));
 sky130_fd_sc_hd__nor2_1 _11997_ (.A(_00208_),
    .B(net58),
    .Y(_04940_));
 sky130_fd_sc_hd__xnor2_1 _11998_ (.A(_04939_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__or2_1 _11999_ (.A(_04937_),
    .B(_04941_),
    .X(_04942_));
 sky130_fd_sc_hd__nand2_1 _12000_ (.A(_04937_),
    .B(_04941_),
    .Y(_04943_));
 sky130_fd_sc_hd__nand2_1 _12001_ (.A(_04942_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__o22a_1 _12002_ (.A1(net50),
    .A2(net34),
    .B1(net32),
    .B2(net52),
    .X(_04945_));
 sky130_fd_sc_hd__xnor2_1 _12003_ (.A(net93),
    .B(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__inv_2 _12004_ (.A(_04946_),
    .Y(_04947_));
 sky130_fd_sc_hd__a22o_1 _12005_ (.A1(_00161_),
    .A2(net16),
    .B1(net12),
    .B2(_00150_),
    .X(_04948_));
 sky130_fd_sc_hd__xnor2_1 _12006_ (.A(net64),
    .B(_04948_),
    .Y(_04950_));
 sky130_fd_sc_hd__a22o_1 _12007_ (.A1(_00177_),
    .A2(net15),
    .B1(net31),
    .B2(_00516_),
    .X(_04951_));
 sky130_fd_sc_hd__xnor2_1 _12008_ (.A(net91),
    .B(_04951_),
    .Y(_04952_));
 sky130_fd_sc_hd__nand2_1 _12009_ (.A(_04950_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__xnor2_1 _12010_ (.A(_04950_),
    .B(_04952_),
    .Y(_04954_));
 sky130_fd_sc_hd__xnor2_1 _12011_ (.A(_04947_),
    .B(_04954_),
    .Y(_04955_));
 sky130_fd_sc_hd__xnor2_1 _12012_ (.A(_04944_),
    .B(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__a32o_1 _12013_ (.A1(_04849_),
    .A2(_04850_),
    .A3(_04859_),
    .B1(_04860_),
    .B2(_04842_),
    .X(_04957_));
 sky130_fd_sc_hd__nand2_1 _12014_ (.A(_04867_),
    .B(_04869_),
    .Y(_04958_));
 sky130_fd_sc_hd__a21bo_1 _12015_ (.A1(_04833_),
    .A2(_04839_),
    .B1_N(_04838_),
    .X(_04959_));
 sky130_fd_sc_hd__nand2_1 _12016_ (.A(_04847_),
    .B(_04849_),
    .Y(_04961_));
 sky130_fd_sc_hd__o21a_1 _12017_ (.A1(_04857_),
    .A2(_04858_),
    .B1(_04855_),
    .X(_04962_));
 sky130_fd_sc_hd__a21oi_1 _12018_ (.A1(_04847_),
    .A2(_04849_),
    .B1(_04962_),
    .Y(_04963_));
 sky130_fd_sc_hd__xnor2_1 _12019_ (.A(_04961_),
    .B(_04962_),
    .Y(_04964_));
 sky130_fd_sc_hd__and2_1 _12020_ (.A(_04959_),
    .B(_04964_),
    .X(_04965_));
 sky130_fd_sc_hd__nor2_1 _12021_ (.A(_04959_),
    .B(_04964_),
    .Y(_04966_));
 sky130_fd_sc_hd__or2_1 _12022_ (.A(_04965_),
    .B(_04966_),
    .X(_04967_));
 sky130_fd_sc_hd__a21oi_1 _12023_ (.A1(_04867_),
    .A2(_04869_),
    .B1(_04967_),
    .Y(_04968_));
 sky130_fd_sc_hd__xnor2_1 _12024_ (.A(_04958_),
    .B(_04967_),
    .Y(_04969_));
 sky130_fd_sc_hd__xnor2_1 _12025_ (.A(_04957_),
    .B(_04969_),
    .Y(_04970_));
 sky130_fd_sc_hd__or2_1 _12026_ (.A(_04956_),
    .B(_04970_),
    .X(_04972_));
 sky130_fd_sc_hd__xor2_1 _12027_ (.A(_04956_),
    .B(_04970_),
    .X(_04973_));
 sky130_fd_sc_hd__o21ai_1 _12028_ (.A1(_04871_),
    .A2(_04875_),
    .B1(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__or3_1 _12029_ (.A(_04871_),
    .B(_04875_),
    .C(_04973_),
    .X(_04975_));
 sky130_fd_sc_hd__and2_1 _12030_ (.A(_04974_),
    .B(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__o21a_1 _12031_ (.A1(_04877_),
    .A2(_04879_),
    .B1(_04976_),
    .X(_04977_));
 sky130_fd_sc_hd__or3_1 _12032_ (.A(_04877_),
    .B(_04879_),
    .C(_04976_),
    .X(_04978_));
 sky130_fd_sc_hd__and2b_2 _12033_ (.A_N(_04977_),
    .B(_04978_),
    .X(_04979_));
 sky130_fd_sc_hd__o21a_1 _12034_ (.A1(_04782_),
    .A2(_04881_),
    .B1(_04882_),
    .X(_04980_));
 sky130_fd_sc_hd__nor2_1 _12035_ (.A(_04784_),
    .B(_04883_),
    .Y(_04981_));
 sky130_fd_sc_hd__a21o_1 _12036_ (.A1(_04785_),
    .A2(_04981_),
    .B1(_04980_),
    .X(_04983_));
 sky130_fd_sc_hd__and2_1 _12037_ (.A(_04787_),
    .B(_04981_),
    .X(_04984_));
 sky130_fd_sc_hd__a21oi_2 _12038_ (.A1(_04589_),
    .A2(_04984_),
    .B1(_04983_),
    .Y(_04985_));
 sky130_fd_sc_hd__xnor2_4 _12039_ (.A(_04979_),
    .B(_04985_),
    .Y(_04986_));
 sky130_fd_sc_hd__a21oi_1 _12040_ (.A1(net138),
    .A2(_04930_),
    .B1(_04986_),
    .Y(_04987_));
 sky130_fd_sc_hd__a31o_1 _12041_ (.A1(net138),
    .A2(_04930_),
    .A3(_04986_),
    .B1(net235),
    .X(_04988_));
 sky130_fd_sc_hd__a21oi_1 _12042_ (.A1(_01976_),
    .A2(_01977_),
    .B1(net135),
    .Y(_04989_));
 sky130_fd_sc_hd__xnor2_1 _12043_ (.A(_01982_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__a21o_1 _12044_ (.A1(_05912_),
    .A2(_04899_),
    .B1(_05902_),
    .X(_04991_));
 sky130_fd_sc_hd__mux2_1 _12045_ (.A0(_06598_),
    .A1(_04991_),
    .S(net283),
    .X(_04992_));
 sky130_fd_sc_hd__nand2_1 _12046_ (.A(_05764_),
    .B(_04992_),
    .Y(_04994_));
 sky130_fd_sc_hd__o211a_1 _12047_ (.A1(_05764_),
    .A2(_04992_),
    .B1(_04994_),
    .C1(net234),
    .X(_04995_));
 sky130_fd_sc_hd__or2_1 _12048_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .X(_04996_));
 sky130_fd_sc_hd__nand2_1 _12049_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .Y(_04997_));
 sky130_fd_sc_hd__nand2_1 _12050_ (.A(_04996_),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__o21a_1 _12051_ (.A1(_04905_),
    .A2(_04907_),
    .B1(_04904_),
    .X(_04999_));
 sky130_fd_sc_hd__xor2_1 _12052_ (.A(_04998_),
    .B(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__mux2_1 _12053_ (.A0(_04052_),
    .A1(_05000_),
    .S(net244),
    .X(_05001_));
 sky130_fd_sc_hd__nor2_1 _12054_ (.A(\div_res[19] ),
    .B(_04913_),
    .Y(_05002_));
 sky130_fd_sc_hd__o21bai_1 _12055_ (.A1(_06681_),
    .A2(_05002_),
    .B1_N(\div_res[20] ),
    .Y(_05003_));
 sky130_fd_sc_hd__or3b_1 _12056_ (.A(_05002_),
    .B(_06681_),
    .C_N(\div_res[20] ),
    .X(_05005_));
 sky130_fd_sc_hd__or2_1 _12057_ (.A(\div_shifter[51] ),
    .B(_04910_),
    .X(_05006_));
 sky130_fd_sc_hd__and2_1 _12058_ (.A(net227),
    .B(_05006_),
    .X(_05007_));
 sky130_fd_sc_hd__o21ai_1 _12059_ (.A1(\div_shifter[52] ),
    .A2(_05007_),
    .B1(_02441_),
    .Y(_05008_));
 sky130_fd_sc_hd__a21oi_1 _12060_ (.A1(\div_shifter[52] ),
    .A2(_05007_),
    .B1(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__o22a_1 _12061_ (.A1(_05731_),
    .A2(net204),
    .B1(net232),
    .B2(reg1_val[20]),
    .X(_05010_));
 sky130_fd_sc_hd__o21ai_1 _12062_ (.A1(_05742_),
    .A2(_02440_),
    .B1(_05010_),
    .Y(_05011_));
 sky130_fd_sc_hd__a221o_1 _12063_ (.A1(_05764_),
    .A2(net196),
    .B1(_02435_),
    .B2(_05753_),
    .C1(_05011_),
    .X(_05012_));
 sky130_fd_sc_hd__a31o_1 _12064_ (.A1(_00269_),
    .A2(_00401_),
    .A3(net256),
    .B1(_05012_),
    .X(_05013_));
 sky130_fd_sc_hd__a221o_1 _12065_ (.A1(net171),
    .A2(_04040_),
    .B1(_04052_),
    .B2(net167),
    .C1(_05013_),
    .X(_05014_));
 sky130_fd_sc_hd__a311o_1 _12066_ (.A1(_02443_),
    .A2(_05003_),
    .A3(_05005_),
    .B1(_05009_),
    .C1(_05014_),
    .X(_05016_));
 sky130_fd_sc_hd__a211oi_4 _12067_ (.A1(net205),
    .A2(_05001_),
    .B1(_05016_),
    .C1(_04995_),
    .Y(_05017_));
 sky130_fd_sc_hd__o221a_1 _12068_ (.A1(_04987_),
    .A2(_04988_),
    .B1(_04990_),
    .B2(_02434_),
    .C1(_05017_),
    .X(_05018_));
 sky130_fd_sc_hd__a21oi_1 _12069_ (.A1(curr_PC[19]),
    .A2(_04827_),
    .B1(curr_PC[20]),
    .Y(_05019_));
 sky130_fd_sc_hd__and3_1 _12070_ (.A(curr_PC[19]),
    .B(curr_PC[20]),
    .C(_04827_),
    .X(_05020_));
 sky130_fd_sc_hd__or3_1 _12071_ (.A(net241),
    .B(_05019_),
    .C(_05020_),
    .X(_05021_));
 sky130_fd_sc_hd__o21ai_4 _12072_ (.A1(net242),
    .A2(_05018_),
    .B1(_05021_),
    .Y(dest_val[20]));
 sky130_fd_sc_hd__o31a_1 _12073_ (.A1(_04830_),
    .A2(_04891_),
    .A3(_04986_),
    .B1(net144),
    .X(_05022_));
 sky130_fd_sc_hd__a21o_1 _12074_ (.A1(_04957_),
    .A2(_04969_),
    .B1(_04968_),
    .X(_05023_));
 sky130_fd_sc_hd__a22o_1 _12075_ (.A1(_00144_),
    .A2(net16),
    .B1(net12),
    .B2(_00161_),
    .X(_05024_));
 sky130_fd_sc_hd__xnor2_1 _12076_ (.A(net64),
    .B(_05024_),
    .Y(_05026_));
 sky130_fd_sc_hd__a22o_1 _12077_ (.A1(_00150_),
    .A2(net8),
    .B1(net3),
    .B2(net55),
    .X(_05027_));
 sky130_fd_sc_hd__xnor2_1 _12078_ (.A(net58),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__o22a_1 _12079_ (.A1(net52),
    .A2(net35),
    .B1(net33),
    .B2(net43),
    .X(_05029_));
 sky130_fd_sc_hd__xnor2_1 _12080_ (.A(net93),
    .B(_05029_),
    .Y(_05030_));
 sky130_fd_sc_hd__nand2_1 _12081_ (.A(_05028_),
    .B(_05030_),
    .Y(_05031_));
 sky130_fd_sc_hd__or2_1 _12082_ (.A(_05028_),
    .B(_05030_),
    .X(_05032_));
 sky130_fd_sc_hd__and2_1 _12083_ (.A(_05031_),
    .B(_05032_),
    .X(_05033_));
 sky130_fd_sc_hd__nand2_1 _12084_ (.A(_05026_),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__or2_1 _12085_ (.A(_05026_),
    .B(_05033_),
    .X(_05035_));
 sky130_fd_sc_hd__nand2_1 _12086_ (.A(_05034_),
    .B(_05035_),
    .Y(_05037_));
 sky130_fd_sc_hd__nor3_1 _12087_ (.A(net41),
    .B(net58),
    .C(_04939_),
    .Y(_05038_));
 sky130_fd_sc_hd__xor2_1 _12088_ (.A(_05037_),
    .B(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__o22a_1 _12089_ (.A1(net38),
    .A2(net10),
    .B1(net5),
    .B2(net36),
    .X(_05040_));
 sky130_fd_sc_hd__xnor2_1 _12090_ (.A(net98),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__a22o_1 _12091_ (.A1(net15),
    .A2(_00516_),
    .B1(_00812_),
    .B2(net31),
    .X(_05042_));
 sky130_fd_sc_hd__xnor2_1 _12092_ (.A(net91),
    .B(_05042_),
    .Y(_05043_));
 sky130_fd_sc_hd__nand2_1 _12093_ (.A(_00274_),
    .B(_05043_),
    .Y(_05044_));
 sky130_fd_sc_hd__xnor2_1 _12094_ (.A(net97),
    .B(_05043_),
    .Y(_05045_));
 sky130_fd_sc_hd__nand2_1 _12095_ (.A(_05041_),
    .B(_05045_),
    .Y(_05046_));
 sky130_fd_sc_hd__or2_1 _12096_ (.A(_05041_),
    .B(_05045_),
    .X(_05048_));
 sky130_fd_sc_hd__nand2_1 _12097_ (.A(_05046_),
    .B(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__nor2_1 _12098_ (.A(_05039_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__and2_1 _12099_ (.A(_05039_),
    .B(_05049_),
    .X(_05051_));
 sky130_fd_sc_hd__nor2_1 _12100_ (.A(_05050_),
    .B(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__o21a_1 _12101_ (.A1(_04944_),
    .A2(_04955_),
    .B1(_04942_),
    .X(_05053_));
 sky130_fd_sc_hd__o21ai_1 _12102_ (.A1(_04947_),
    .A2(_04954_),
    .B1(_04953_),
    .Y(_05054_));
 sky130_fd_sc_hd__nor2_1 _12103_ (.A(net57),
    .B(net58),
    .Y(_05055_));
 sky130_fd_sc_hd__and2_1 _12104_ (.A(_05054_),
    .B(_05055_),
    .X(_05056_));
 sky130_fd_sc_hd__xnor2_1 _12105_ (.A(_05054_),
    .B(_05055_),
    .Y(_05057_));
 sky130_fd_sc_hd__nor2_1 _12106_ (.A(_04935_),
    .B(_05057_),
    .Y(_05059_));
 sky130_fd_sc_hd__and2_1 _12107_ (.A(_04935_),
    .B(_05057_),
    .X(_05060_));
 sky130_fd_sc_hd__nor2_1 _12108_ (.A(_05059_),
    .B(_05060_),
    .Y(_05061_));
 sky130_fd_sc_hd__o21ai_1 _12109_ (.A1(_04963_),
    .A2(_04965_),
    .B1(_05061_),
    .Y(_05062_));
 sky130_fd_sc_hd__or3_1 _12110_ (.A(_04963_),
    .B(_04965_),
    .C(_05061_),
    .X(_05063_));
 sky130_fd_sc_hd__nand2_1 _12111_ (.A(_05062_),
    .B(_05063_),
    .Y(_05064_));
 sky130_fd_sc_hd__xor2_1 _12112_ (.A(_05053_),
    .B(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__nand2_1 _12113_ (.A(_05052_),
    .B(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__or2_1 _12114_ (.A(_05052_),
    .B(_05065_),
    .X(_05067_));
 sky130_fd_sc_hd__and2_1 _12115_ (.A(_05066_),
    .B(_05067_),
    .X(_05068_));
 sky130_fd_sc_hd__nand2_1 _12116_ (.A(_05023_),
    .B(_05068_),
    .Y(_05070_));
 sky130_fd_sc_hd__xnor2_1 _12117_ (.A(_05023_),
    .B(_05068_),
    .Y(_05071_));
 sky130_fd_sc_hd__a21o_1 _12118_ (.A1(_04972_),
    .A2(_04974_),
    .B1(_05071_),
    .X(_05072_));
 sky130_fd_sc_hd__inv_2 _12119_ (.A(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__nand3_1 _12120_ (.A(_04972_),
    .B(_04974_),
    .C(_05071_),
    .Y(_05074_));
 sky130_fd_sc_hd__and2_2 _12121_ (.A(_05072_),
    .B(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__o21ai_1 _12122_ (.A1(_04881_),
    .A2(_04977_),
    .B1(_04978_),
    .Y(_05076_));
 sky130_fd_sc_hd__nand2b_1 _12123_ (.A_N(_04883_),
    .B(_04979_),
    .Y(_05077_));
 sky130_fd_sc_hd__o21ai_2 _12124_ (.A1(_04886_),
    .A2(_05077_),
    .B1(_05076_),
    .Y(_05078_));
 sky130_fd_sc_hd__and3b_1 _12125_ (.A_N(_04883_),
    .B(_04887_),
    .C(_04979_),
    .X(_05079_));
 sky130_fd_sc_hd__a21oi_2 _12126_ (.A1(_04692_),
    .A2(_05079_),
    .B1(_05078_),
    .Y(_05081_));
 sky130_fd_sc_hd__xnor2_4 _12127_ (.A(_05075_),
    .B(_05081_),
    .Y(_05082_));
 sky130_fd_sc_hd__and2_1 _12128_ (.A(_05022_),
    .B(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__nor2_1 _12129_ (.A(_05022_),
    .B(_05082_),
    .Y(_05084_));
 sky130_fd_sc_hd__and2_1 _12130_ (.A(net137),
    .B(_01983_),
    .X(_05085_));
 sky130_fd_sc_hd__nor2_1 _12131_ (.A(_01984_),
    .B(_05085_),
    .Y(_05086_));
 sky130_fd_sc_hd__a211o_1 _12132_ (.A1(_01984_),
    .A2(_05085_),
    .B1(_05086_),
    .C1(_02434_),
    .X(_05087_));
 sky130_fd_sc_hd__a21o_1 _12133_ (.A1(_05764_),
    .A2(_04991_),
    .B1(_05753_),
    .X(_05088_));
 sky130_fd_sc_hd__o21a_1 _12134_ (.A1(_05764_),
    .A2(_06598_),
    .B1(_06603_),
    .X(_05089_));
 sky130_fd_sc_hd__mux2_1 _12135_ (.A0(_05088_),
    .A1(_05089_),
    .S(net296),
    .X(_05090_));
 sky130_fd_sc_hd__nor2_1 _12136_ (.A(_05835_),
    .B(_05090_),
    .Y(_05092_));
 sky130_fd_sc_hd__a21o_1 _12137_ (.A1(_05835_),
    .A2(_05090_),
    .B1(_02427_),
    .X(_05093_));
 sky130_fd_sc_hd__or2_1 _12138_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .X(_05094_));
 sky130_fd_sc_hd__nand2_1 _12139_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .Y(_05095_));
 sky130_fd_sc_hd__nand2_1 _12140_ (.A(_05094_),
    .B(_05095_),
    .Y(_05096_));
 sky130_fd_sc_hd__o21a_1 _12141_ (.A1(_04998_),
    .A2(_04999_),
    .B1(_04997_),
    .X(_05097_));
 sky130_fd_sc_hd__xnor2_1 _12142_ (.A(_05096_),
    .B(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__nor2_1 _12143_ (.A(net245),
    .B(_03925_),
    .Y(_05099_));
 sky130_fd_sc_hd__a211o_1 _12144_ (.A1(net245),
    .A2(_05098_),
    .B1(_05099_),
    .C1(_06667_),
    .X(_05100_));
 sky130_fd_sc_hd__or2_1 _12145_ (.A(\div_shifter[52] ),
    .B(_05006_),
    .X(_05101_));
 sky130_fd_sc_hd__a21oi_1 _12146_ (.A1(net227),
    .A2(_05101_),
    .B1(\div_shifter[53] ),
    .Y(_05103_));
 sky130_fd_sc_hd__a31o_1 _12147_ (.A1(\div_shifter[53] ),
    .A2(net227),
    .A3(_05101_),
    .B1(net191),
    .X(_05104_));
 sky130_fd_sc_hd__or3_1 _12148_ (.A(\div_res[20] ),
    .B(\div_res[19] ),
    .C(_04913_),
    .X(_05105_));
 sky130_fd_sc_hd__a21oi_1 _12149_ (.A1(net141),
    .A2(_05105_),
    .B1(\div_res[21] ),
    .Y(_05106_));
 sky130_fd_sc_hd__a31o_1 _12150_ (.A1(\div_res[21] ),
    .A2(net141),
    .A3(_05105_),
    .B1(net189),
    .X(_05107_));
 sky130_fd_sc_hd__or2_1 _12151_ (.A(_05106_),
    .B(_05107_),
    .X(_05108_));
 sky130_fd_sc_hd__o22ai_1 _12152_ (.A1(_05826_),
    .A2(_02440_),
    .B1(net232),
    .B2(reg1_val[21]),
    .Y(_05109_));
 sky130_fd_sc_hd__a221o_1 _12153_ (.A1(_05835_),
    .A2(net196),
    .B1(_02435_),
    .B2(_05816_),
    .C1(_05109_),
    .X(_05110_));
 sky130_fd_sc_hd__a221o_1 _12154_ (.A1(net172),
    .A2(_03911_),
    .B1(_03925_),
    .B2(net167),
    .C1(_05110_),
    .X(_05111_));
 sky130_fd_sc_hd__a21oi_1 _12155_ (.A1(_00271_),
    .A2(net257),
    .B1(_05111_),
    .Y(_05112_));
 sky130_fd_sc_hd__o211a_1 _12156_ (.A1(_05103_),
    .A2(_05104_),
    .B1(_05108_),
    .C1(_05112_),
    .X(_05114_));
 sky130_fd_sc_hd__o211a_1 _12157_ (.A1(_05092_),
    .A2(_05093_),
    .B1(_05100_),
    .C1(_05114_),
    .X(_05115_));
 sky130_fd_sc_hd__o311a_1 _12158_ (.A1(net235),
    .A2(_05083_),
    .A3(_05084_),
    .B1(_05087_),
    .C1(_05115_),
    .X(_05116_));
 sky130_fd_sc_hd__o22a_1 _12159_ (.A1(_05796_),
    .A2(net203),
    .B1(_06679_),
    .B2(_05116_),
    .X(_05117_));
 sky130_fd_sc_hd__and2_2 _12160_ (.A(curr_PC[21]),
    .B(_05020_),
    .X(_05118_));
 sky130_fd_sc_hd__o21ai_1 _12161_ (.A1(curr_PC[21]),
    .A2(_05020_),
    .B1(net242),
    .Y(_05119_));
 sky130_fd_sc_hd__o22ai_4 _12162_ (.A1(net243),
    .A2(_05117_),
    .B1(_05118_),
    .B2(_05119_),
    .Y(dest_val[21]));
 sky130_fd_sc_hd__or3_1 _12163_ (.A(_04590_),
    .B(_04693_),
    .C(_04792_),
    .X(_05120_));
 sky130_fd_sc_hd__nor4_2 _12164_ (.A(_04891_),
    .B(_04986_),
    .C(_05082_),
    .D(_05120_),
    .Y(_05121_));
 sky130_fd_sc_hd__nand2b_1 _12165_ (.A_N(_04516_),
    .B(_05121_),
    .Y(_05122_));
 sky130_fd_sc_hd__o21ai_1 _12166_ (.A1(_05053_),
    .A2(_05064_),
    .B1(_05062_),
    .Y(_05124_));
 sky130_fd_sc_hd__o22a_1 _12167_ (.A1(net43),
    .A2(net35),
    .B1(net33),
    .B2(_00517_),
    .X(_05125_));
 sky130_fd_sc_hd__xnor2_2 _12168_ (.A(net93),
    .B(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__a22o_1 _12169_ (.A1(_00136_),
    .A2(net16),
    .B1(net12),
    .B2(_00144_),
    .X(_05127_));
 sky130_fd_sc_hd__xnor2_1 _12170_ (.A(net64),
    .B(_05127_),
    .Y(_05128_));
 sky130_fd_sc_hd__xnor2_1 _12171_ (.A(_05126_),
    .B(_05128_),
    .Y(_05129_));
 sky130_fd_sc_hd__a21o_1 _12172_ (.A1(_05031_),
    .A2(_05034_),
    .B1(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__nand3_1 _12173_ (.A(_05031_),
    .B(_05034_),
    .C(_05129_),
    .Y(_05131_));
 sky130_fd_sc_hd__nand2_1 _12174_ (.A(_05130_),
    .B(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__a22o_1 _12175_ (.A1(net15),
    .A2(_00812_),
    .B1(_02065_),
    .B2(net31),
    .X(_05133_));
 sky130_fd_sc_hd__xnor2_1 _12176_ (.A(_00309_),
    .B(_05133_),
    .Y(_05135_));
 sky130_fd_sc_hd__or2_1 _12177_ (.A(_00279_),
    .B(net5),
    .X(_05136_));
 sky130_fd_sc_hd__a22o_1 _12178_ (.A1(_00281_),
    .A2(net7),
    .B1(_05136_),
    .B2(net98),
    .X(_05137_));
 sky130_fd_sc_hd__nor2_1 _12179_ (.A(_05135_),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__and2_1 _12180_ (.A(_05135_),
    .B(_05137_),
    .X(_05139_));
 sky130_fd_sc_hd__nor2_1 _12181_ (.A(_05138_),
    .B(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__xnor2_1 _12182_ (.A(_05132_),
    .B(_05140_),
    .Y(_05141_));
 sky130_fd_sc_hd__a31o_1 _12183_ (.A1(_05034_),
    .A2(_05035_),
    .A3(_05038_),
    .B1(_05050_),
    .X(_05142_));
 sky130_fd_sc_hd__a22o_1 _12184_ (.A1(_00161_),
    .A2(net8),
    .B1(net3),
    .B2(_00150_),
    .X(_05143_));
 sky130_fd_sc_hd__xnor2_1 _12185_ (.A(net61),
    .B(_05143_),
    .Y(_05144_));
 sky130_fd_sc_hd__a21oi_1 _12186_ (.A1(_05044_),
    .A2(_05046_),
    .B1(_05144_),
    .Y(_05146_));
 sky130_fd_sc_hd__and3_1 _12187_ (.A(_05044_),
    .B(_05046_),
    .C(_05144_),
    .X(_05147_));
 sky130_fd_sc_hd__nor2_1 _12188_ (.A(_05146_),
    .B(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__nand2_1 _12189_ (.A(net55),
    .B(net61),
    .Y(_05149_));
 sky130_fd_sc_hd__xnor2_1 _12190_ (.A(_05148_),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__o21ai_1 _12191_ (.A1(_05056_),
    .A2(_05059_),
    .B1(_05150_),
    .Y(_05151_));
 sky130_fd_sc_hd__or3_1 _12192_ (.A(_05056_),
    .B(_05059_),
    .C(_05150_),
    .X(_05152_));
 sky130_fd_sc_hd__and2_1 _12193_ (.A(_05151_),
    .B(_05152_),
    .X(_05153_));
 sky130_fd_sc_hd__nand2_1 _12194_ (.A(_05142_),
    .B(_05153_),
    .Y(_05154_));
 sky130_fd_sc_hd__xnor2_1 _12195_ (.A(_05142_),
    .B(_05153_),
    .Y(_05155_));
 sky130_fd_sc_hd__or2_1 _12196_ (.A(_05141_),
    .B(_05155_),
    .X(_05157_));
 sky130_fd_sc_hd__nand2_1 _12197_ (.A(_05141_),
    .B(_05155_),
    .Y(_05158_));
 sky130_fd_sc_hd__nand2_1 _12198_ (.A(_05157_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__nand2b_1 _12199_ (.A_N(_05159_),
    .B(_05124_),
    .Y(_05160_));
 sky130_fd_sc_hd__xor2_1 _12200_ (.A(_05124_),
    .B(_05159_),
    .X(_05161_));
 sky130_fd_sc_hd__a21o_1 _12201_ (.A1(_05066_),
    .A2(_05070_),
    .B1(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__inv_2 _12202_ (.A(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__and3_1 _12203_ (.A(_05066_),
    .B(_05070_),
    .C(_05161_),
    .X(_05164_));
 sky130_fd_sc_hd__nor2_2 _12204_ (.A(_05163_),
    .B(_05164_),
    .Y(_05165_));
 sky130_fd_sc_hd__o21ai_1 _12205_ (.A1(_04977_),
    .A2(_05073_),
    .B1(_05074_),
    .Y(_05166_));
 sky130_fd_sc_hd__nand2_1 _12206_ (.A(_04979_),
    .B(_05075_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand3_1 _12207_ (.A(_04979_),
    .B(_04980_),
    .C(_05075_),
    .Y(_05169_));
 sky130_fd_sc_hd__and2_1 _12208_ (.A(_05166_),
    .B(_05169_),
    .X(_05170_));
 sky130_fd_sc_hd__o41a_2 _12209_ (.A1(_04784_),
    .A2(_04791_),
    .A3(_04883_),
    .A4(_05168_),
    .B1(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__xnor2_4 _12210_ (.A(_05165_),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__a21oi_1 _12211_ (.A1(net138),
    .A2(_05122_),
    .B1(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__a31o_1 _12212_ (.A1(net138),
    .A2(_05122_),
    .A3(_05172_),
    .B1(net235),
    .X(_05174_));
 sky130_fd_sc_hd__nand2_1 _12213_ (.A(net138),
    .B(_01987_),
    .Y(_05175_));
 sky130_fd_sc_hd__xnor2_1 _12214_ (.A(_01993_),
    .B(_05175_),
    .Y(_05176_));
 sky130_fd_sc_hd__a21o_1 _12215_ (.A1(_05835_),
    .A2(_05088_),
    .B1(_05816_),
    .X(_05177_));
 sky130_fd_sc_hd__o21a_1 _12216_ (.A1(_05835_),
    .A2(_05089_),
    .B1(_06602_),
    .X(_05179_));
 sky130_fd_sc_hd__mux2_1 _12217_ (.A0(_05177_),
    .A1(_05179_),
    .S(net296),
    .X(_05180_));
 sky130_fd_sc_hd__nand2_1 _12218_ (.A(_05699_),
    .B(_05180_),
    .Y(_05181_));
 sky130_fd_sc_hd__o21a_1 _12219_ (.A1(_05699_),
    .A2(_05180_),
    .B1(_02426_),
    .X(_05182_));
 sky130_fd_sc_hd__or2_1 _12220_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .X(_05183_));
 sky130_fd_sc_hd__nand2_1 _12221_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .Y(_05184_));
 sky130_fd_sc_hd__nand2_1 _12222_ (.A(_05183_),
    .B(_05184_),
    .Y(_05185_));
 sky130_fd_sc_hd__o21a_1 _12223_ (.A1(_05096_),
    .A2(_05097_),
    .B1(_05095_),
    .X(_05186_));
 sky130_fd_sc_hd__xor2_1 _12224_ (.A(_05185_),
    .B(_05186_),
    .X(_05187_));
 sky130_fd_sc_hd__nand2_1 _12225_ (.A(net224),
    .B(_03805_),
    .Y(_05188_));
 sky130_fd_sc_hd__o211a_1 _12226_ (.A1(net224),
    .A2(_05187_),
    .B1(_05188_),
    .C1(_06666_),
    .X(_05190_));
 sky130_fd_sc_hd__or2_1 _12227_ (.A(\div_res[21] ),
    .B(_05105_),
    .X(_05191_));
 sky130_fd_sc_hd__a21oi_1 _12228_ (.A1(net141),
    .A2(_05191_),
    .B1(\div_res[22] ),
    .Y(_05192_));
 sky130_fd_sc_hd__a31o_1 _12229_ (.A1(\div_res[22] ),
    .A2(net141),
    .A3(_05191_),
    .B1(net189),
    .X(_05193_));
 sky130_fd_sc_hd__nor2_1 _12230_ (.A(_05192_),
    .B(_05193_),
    .Y(_05194_));
 sky130_fd_sc_hd__or2_1 _12231_ (.A(\div_shifter[53] ),
    .B(_05101_),
    .X(_05195_));
 sky130_fd_sc_hd__a21oi_1 _12232_ (.A1(net230),
    .A2(_05195_),
    .B1(\div_shifter[54] ),
    .Y(_05196_));
 sky130_fd_sc_hd__a31o_1 _12233_ (.A1(\div_shifter[54] ),
    .A2(net230),
    .A3(_05195_),
    .B1(net192),
    .X(_05197_));
 sky130_fd_sc_hd__nor2_1 _12234_ (.A(_05196_),
    .B(_05197_),
    .Y(_05198_));
 sky130_fd_sc_hd__and3_1 _12235_ (.A(_00259_),
    .B(_00275_),
    .C(net256),
    .X(_05199_));
 sky130_fd_sc_hd__a21o_1 _12236_ (.A1(_04543_),
    .A2(_05656_),
    .B1(_02440_),
    .X(_05201_));
 sky130_fd_sc_hd__o221a_1 _12237_ (.A1(_05656_),
    .A2(net204),
    .B1(net232),
    .B2(reg1_val[22]),
    .C1(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__o21ai_1 _12238_ (.A1(_05677_),
    .A2(_02436_),
    .B1(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__a221o_1 _12239_ (.A1(_05699_),
    .A2(net195),
    .B1(_03806_),
    .B2(net167),
    .C1(_05203_),
    .X(_05204_));
 sky130_fd_sc_hd__a211o_1 _12240_ (.A1(net171),
    .A2(_03789_),
    .B1(_05199_),
    .C1(_05204_),
    .X(_05205_));
 sky130_fd_sc_hd__or4_1 _12241_ (.A(_05190_),
    .B(_05194_),
    .C(_05198_),
    .D(_05205_),
    .X(_05206_));
 sky130_fd_sc_hd__a21oi_1 _12242_ (.A1(_05181_),
    .A2(_05182_),
    .B1(_05206_),
    .Y(_05207_));
 sky130_fd_sc_hd__o221a_1 _12243_ (.A1(_05173_),
    .A2(_05174_),
    .B1(_05176_),
    .B2(_02434_),
    .C1(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__o21ai_1 _12244_ (.A1(curr_PC[22]),
    .A2(_05118_),
    .B1(net243),
    .Y(_05209_));
 sky130_fd_sc_hd__a21o_1 _12245_ (.A1(curr_PC[22]),
    .A2(_05118_),
    .B1(_05209_),
    .X(_05210_));
 sky130_fd_sc_hd__o21ai_4 _12246_ (.A1(net243),
    .A2(_05208_),
    .B1(_05210_),
    .Y(dest_val[22]));
 sky130_fd_sc_hd__o21a_1 _12247_ (.A1(_05122_),
    .A2(_05172_),
    .B1(net144),
    .X(_05212_));
 sky130_fd_sc_hd__a22o_1 _12248_ (.A1(net15),
    .A2(_02065_),
    .B1(net7),
    .B2(net31),
    .X(_05213_));
 sky130_fd_sc_hd__xnor2_1 _12249_ (.A(_00309_),
    .B(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__o22a_1 _12250_ (.A1(net35),
    .A2(_00517_),
    .B1(_00811_),
    .B2(net33),
    .X(_05215_));
 sky130_fd_sc_hd__xnor2_1 _12251_ (.A(net93),
    .B(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__nand2_1 _12252_ (.A(_00263_),
    .B(_05216_),
    .Y(_05217_));
 sky130_fd_sc_hd__xnor2_1 _12253_ (.A(net98),
    .B(_05216_),
    .Y(_05218_));
 sky130_fd_sc_hd__nand2_1 _12254_ (.A(_05214_),
    .B(_05218_),
    .Y(_05219_));
 sky130_fd_sc_hd__or2_1 _12255_ (.A(_05214_),
    .B(_05218_),
    .X(_05220_));
 sky130_fd_sc_hd__nand2_1 _12256_ (.A(_05219_),
    .B(_05220_),
    .Y(_05222_));
 sky130_fd_sc_hd__or2_1 _12257_ (.A(_05138_),
    .B(_05222_),
    .X(_05223_));
 sky130_fd_sc_hd__nand2_1 _12258_ (.A(_05138_),
    .B(_05222_),
    .Y(_05224_));
 sky130_fd_sc_hd__and2_1 _12259_ (.A(_05223_),
    .B(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__nand3_1 _12260_ (.A(_05126_),
    .B(_05128_),
    .C(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__a21o_1 _12261_ (.A1(_05126_),
    .A2(_05128_),
    .B1(_05225_),
    .X(_05227_));
 sky130_fd_sc_hd__and2_1 _12262_ (.A(_05226_),
    .B(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__o21a_1 _12263_ (.A1(_05132_),
    .A2(_05140_),
    .B1(_05130_),
    .X(_05229_));
 sky130_fd_sc_hd__a22o_1 _12264_ (.A1(_00144_),
    .A2(net8),
    .B1(net3),
    .B2(_00161_),
    .X(_05230_));
 sky130_fd_sc_hd__xnor2_1 _12265_ (.A(net61),
    .B(_05230_),
    .Y(_05231_));
 sky130_fd_sc_hd__a22o_1 _12266_ (.A1(_00177_),
    .A2(net16),
    .B1(net12),
    .B2(_00136_),
    .X(_05233_));
 sky130_fd_sc_hd__xnor2_1 _12267_ (.A(net64),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__nor2_1 _12268_ (.A(net48),
    .B(net58),
    .Y(_05235_));
 sky130_fd_sc_hd__nand2_1 _12269_ (.A(_05234_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__xnor2_1 _12270_ (.A(_05234_),
    .B(_05235_),
    .Y(_05237_));
 sky130_fd_sc_hd__or2_1 _12271_ (.A(_05231_),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__nand2_1 _12272_ (.A(_05231_),
    .B(_05237_),
    .Y(_05239_));
 sky130_fd_sc_hd__nand2_1 _12273_ (.A(_05238_),
    .B(_05239_),
    .Y(_05240_));
 sky130_fd_sc_hd__a31o_1 _12274_ (.A1(net55),
    .A2(net61),
    .A3(_05148_),
    .B1(_05146_),
    .X(_05241_));
 sky130_fd_sc_hd__nand2b_1 _12275_ (.A_N(_05240_),
    .B(_05241_),
    .Y(_05242_));
 sky130_fd_sc_hd__xnor2_1 _12276_ (.A(_05240_),
    .B(_05241_),
    .Y(_05244_));
 sky130_fd_sc_hd__nand2b_1 _12277_ (.A_N(_05229_),
    .B(_05244_),
    .Y(_05245_));
 sky130_fd_sc_hd__xnor2_1 _12278_ (.A(_05229_),
    .B(_05244_),
    .Y(_05246_));
 sky130_fd_sc_hd__nand2_1 _12279_ (.A(_05228_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__or2_1 _12280_ (.A(_05228_),
    .B(_05246_),
    .X(_05248_));
 sky130_fd_sc_hd__nand2_1 _12281_ (.A(_05247_),
    .B(_05248_),
    .Y(_05249_));
 sky130_fd_sc_hd__a21o_1 _12282_ (.A1(_05151_),
    .A2(_05154_),
    .B1(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__nand3_1 _12283_ (.A(_05151_),
    .B(_05154_),
    .C(_05249_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_1 _12284_ (.A(_05250_),
    .B(_05251_),
    .Y(_05252_));
 sky130_fd_sc_hd__a21o_1 _12285_ (.A1(_05157_),
    .A2(_05160_),
    .B1(_05252_),
    .X(_05253_));
 sky130_fd_sc_hd__and3_1 _12286_ (.A(_05157_),
    .B(_05160_),
    .C(_05252_),
    .X(_05255_));
 sky130_fd_sc_hd__inv_2 _12287_ (.A(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_2 _12288_ (.A(_05253_),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__nand2_1 _12289_ (.A(_05075_),
    .B(_05165_),
    .Y(_05258_));
 sky130_fd_sc_hd__nor2_1 _12290_ (.A(_05077_),
    .B(_05258_),
    .Y(_05259_));
 sky130_fd_sc_hd__a21o_1 _12291_ (.A1(_05072_),
    .A2(_05162_),
    .B1(_05164_),
    .X(_05260_));
 sky130_fd_sc_hd__o21ai_1 _12292_ (.A1(_05076_),
    .A2(_05258_),
    .B1(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__and2b_1 _12293_ (.A_N(_04888_),
    .B(_05259_),
    .X(_05262_));
 sky130_fd_sc_hd__a311o_2 _12294_ (.A1(_04470_),
    .A2(_04889_),
    .A3(_05259_),
    .B1(_05261_),
    .C1(_05262_),
    .X(_05263_));
 sky130_fd_sc_hd__xnor2_4 _12295_ (.A(_05257_),
    .B(_05263_),
    .Y(_05264_));
 sky130_fd_sc_hd__nor2_1 _12296_ (.A(_05212_),
    .B(_05264_),
    .Y(_05266_));
 sky130_fd_sc_hd__a21o_1 _12297_ (.A1(_05212_),
    .A2(_05264_),
    .B1(net235),
    .X(_05267_));
 sky130_fd_sc_hd__a21o_1 _12298_ (.A1(_01986_),
    .A2(_01993_),
    .B1(net135),
    .X(_05268_));
 sky130_fd_sc_hd__xor2_1 _12299_ (.A(_01994_),
    .B(_05268_),
    .X(_05269_));
 sky130_fd_sc_hd__o211a_1 _12300_ (.A1(_05699_),
    .A2(_05179_),
    .B1(_06601_),
    .C1(net296),
    .X(_05270_));
 sky130_fd_sc_hd__a21bo_1 _12301_ (.A1(_05699_),
    .A2(_05177_),
    .B1_N(_05677_),
    .X(_05271_));
 sky130_fd_sc_hd__a21o_1 _12302_ (.A1(net283),
    .A2(_05271_),
    .B1(_05270_),
    .X(_05272_));
 sky130_fd_sc_hd__nand2_1 _12303_ (.A(_05623_),
    .B(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__o211a_1 _12304_ (.A1(_05623_),
    .A2(_05272_),
    .B1(_05273_),
    .C1(_02426_),
    .X(_05274_));
 sky130_fd_sc_hd__nor2_1 _12305_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .Y(_05275_));
 sky130_fd_sc_hd__nand2_1 _12306_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .Y(_05277_));
 sky130_fd_sc_hd__and2b_1 _12307_ (.A_N(_05275_),
    .B(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__o21a_1 _12308_ (.A1(_05185_),
    .A2(_05186_),
    .B1(_05184_),
    .X(_05279_));
 sky130_fd_sc_hd__xnor2_1 _12309_ (.A(_05278_),
    .B(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__mux2_1 _12310_ (.A0(_03670_),
    .A1(_05280_),
    .S(net245),
    .X(_05281_));
 sky130_fd_sc_hd__o21ai_1 _12311_ (.A1(\div_res[22] ),
    .A2(_05191_),
    .B1(net141),
    .Y(_05282_));
 sky130_fd_sc_hd__xnor2_1 _12312_ (.A(\div_res[23] ),
    .B(_05282_),
    .Y(_05283_));
 sky130_fd_sc_hd__or2_1 _12313_ (.A(\div_shifter[54] ),
    .B(_05195_),
    .X(_05284_));
 sky130_fd_sc_hd__and2_1 _12314_ (.A(net230),
    .B(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__o21ai_1 _12315_ (.A1(\div_shifter[55] ),
    .A2(_05285_),
    .B1(_02441_),
    .Y(_05286_));
 sky130_fd_sc_hd__a21oi_1 _12316_ (.A1(\div_shifter[55] ),
    .A2(_05285_),
    .B1(_05286_),
    .Y(_05288_));
 sky130_fd_sc_hd__o22a_1 _12317_ (.A1(_05591_),
    .A2(net204),
    .B1(net232),
    .B2(reg1_val[23]),
    .X(_05289_));
 sky130_fd_sc_hd__o21ai_1 _12318_ (.A1(_05612_),
    .A2(_02440_),
    .B1(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__a221o_1 _12319_ (.A1(_05623_),
    .A2(net195),
    .B1(_02435_),
    .B2(_05602_),
    .C1(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__a221o_1 _12320_ (.A1(net171),
    .A2(_03656_),
    .B1(_03670_),
    .B2(net167),
    .C1(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__a31o_1 _12321_ (.A1(_00256_),
    .A2(_00260_),
    .A3(net256),
    .B1(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__a211o_1 _12322_ (.A1(_02443_),
    .A2(_05283_),
    .B1(_05288_),
    .C1(_05293_),
    .X(_05294_));
 sky130_fd_sc_hd__a211oi_1 _12323_ (.A1(_06666_),
    .A2(_05281_),
    .B1(_05294_),
    .C1(_05274_),
    .Y(_05295_));
 sky130_fd_sc_hd__o221a_1 _12324_ (.A1(_05266_),
    .A2(_05267_),
    .B1(_05269_),
    .B2(_02434_),
    .C1(_05295_),
    .X(_05296_));
 sky130_fd_sc_hd__and3_1 _12325_ (.A(curr_PC[22]),
    .B(curr_PC[23]),
    .C(_05118_),
    .X(_05297_));
 sky130_fd_sc_hd__a21oi_1 _12326_ (.A1(curr_PC[22]),
    .A2(_05118_),
    .B1(curr_PC[23]),
    .Y(_05299_));
 sky130_fd_sc_hd__or3_1 _12327_ (.A(net241),
    .B(_05297_),
    .C(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__o21ai_4 _12328_ (.A1(net243),
    .A2(_05296_),
    .B1(_05300_),
    .Y(dest_val[23]));
 sky130_fd_sc_hd__nand2_1 _12329_ (.A(_00332_),
    .B(net7),
    .Y(_05301_));
 sky130_fd_sc_hd__a22o_2 _12330_ (.A1(_00335_),
    .A2(net7),
    .B1(_05301_),
    .B2(net92),
    .X(_05302_));
 sky130_fd_sc_hd__nand2_1 _12331_ (.A(_00161_),
    .B(net61),
    .Y(_05303_));
 sky130_fd_sc_hd__xnor2_1 _12332_ (.A(_05302_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__a21o_1 _12333_ (.A1(_05217_),
    .A2(_05219_),
    .B1(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__nand3_1 _12334_ (.A(_05217_),
    .B(_05219_),
    .C(_05304_),
    .Y(_05306_));
 sky130_fd_sc_hd__and2_1 _12335_ (.A(_05305_),
    .B(_05306_),
    .X(_05307_));
 sky130_fd_sc_hd__nand2_1 _12336_ (.A(_05223_),
    .B(_05226_),
    .Y(_05309_));
 sky130_fd_sc_hd__a22o_1 _12337_ (.A1(_00516_),
    .A2(net16),
    .B1(net12),
    .B2(_00177_),
    .X(_05310_));
 sky130_fd_sc_hd__xnor2_1 _12338_ (.A(net64),
    .B(_05310_),
    .Y(_05311_));
 sky130_fd_sc_hd__a22o_1 _12339_ (.A1(_00136_),
    .A2(net8),
    .B1(net3),
    .B2(_00144_),
    .X(_05312_));
 sky130_fd_sc_hd__xnor2_1 _12340_ (.A(net58),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__o22a_1 _12341_ (.A1(net35),
    .A2(_00811_),
    .B1(net10),
    .B2(net33),
    .X(_05314_));
 sky130_fd_sc_hd__xnor2_1 _12342_ (.A(net93),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__nand2_1 _12343_ (.A(_05313_),
    .B(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__or2_1 _12344_ (.A(_05313_),
    .B(_05315_),
    .X(_05317_));
 sky130_fd_sc_hd__nand2_1 _12345_ (.A(_05316_),
    .B(_05317_),
    .Y(_05318_));
 sky130_fd_sc_hd__inv_2 _12346_ (.A(_05318_),
    .Y(_05320_));
 sky130_fd_sc_hd__nand2_1 _12347_ (.A(_05311_),
    .B(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__or2_1 _12348_ (.A(_05311_),
    .B(_05320_),
    .X(_05322_));
 sky130_fd_sc_hd__nand2_1 _12349_ (.A(_05321_),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__a21o_1 _12350_ (.A1(_05236_),
    .A2(_05238_),
    .B1(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__nand3_1 _12351_ (.A(_05236_),
    .B(_05238_),
    .C(_05323_),
    .Y(_05325_));
 sky130_fd_sc_hd__nand2_1 _12352_ (.A(_05324_),
    .B(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__xnor2_1 _12353_ (.A(_05309_),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__nand2_1 _12354_ (.A(_05307_),
    .B(_05327_),
    .Y(_05328_));
 sky130_fd_sc_hd__or2_1 _12355_ (.A(_05307_),
    .B(_05327_),
    .X(_05329_));
 sky130_fd_sc_hd__nand2_1 _12356_ (.A(_05328_),
    .B(_05329_),
    .Y(_05331_));
 sky130_fd_sc_hd__a21o_1 _12357_ (.A1(_05242_),
    .A2(_05245_),
    .B1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__nand3_1 _12358_ (.A(_05242_),
    .B(_05245_),
    .C(_05331_),
    .Y(_05333_));
 sky130_fd_sc_hd__nand2_1 _12359_ (.A(_05332_),
    .B(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__a21oi_2 _12360_ (.A1(_05247_),
    .A2(_05250_),
    .B1(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__inv_2 _12361_ (.A(_05335_),
    .Y(_05336_));
 sky130_fd_sc_hd__and3_1 _12362_ (.A(_05247_),
    .B(_05250_),
    .C(_05334_),
    .X(_05337_));
 sky130_fd_sc_hd__or2_2 _12363_ (.A(_05335_),
    .B(_05337_),
    .X(_05338_));
 sky130_fd_sc_hd__a21o_1 _12364_ (.A1(_05162_),
    .A2(_05253_),
    .B1(_05255_),
    .X(_05339_));
 sky130_fd_sc_hd__or3_2 _12365_ (.A(_05163_),
    .B(_05164_),
    .C(_05257_),
    .X(_05340_));
 sky130_fd_sc_hd__o21ai_1 _12366_ (.A1(_05166_),
    .A2(_05340_),
    .B1(_05339_),
    .Y(_05342_));
 sky130_fd_sc_hd__nor2_1 _12367_ (.A(_05168_),
    .B(_05340_),
    .Y(_05343_));
 sky130_fd_sc_hd__or3_1 _12368_ (.A(_04985_),
    .B(_05168_),
    .C(_05340_),
    .X(_05344_));
 sky130_fd_sc_hd__and2_1 _12369_ (.A(_04983_),
    .B(_05343_),
    .X(_05345_));
 sky130_fd_sc_hd__a311o_2 _12370_ (.A1(_04589_),
    .A2(_04984_),
    .A3(_05343_),
    .B1(_05345_),
    .C1(_05342_),
    .X(_05346_));
 sky130_fd_sc_hd__xor2_4 _12371_ (.A(_05338_),
    .B(_05346_),
    .X(_05347_));
 sky130_fd_sc_hd__nor4_2 _12372_ (.A(_04059_),
    .B(_04515_),
    .C(_05172_),
    .D(_05264_),
    .Y(_05348_));
 sky130_fd_sc_hd__nand2_2 _12373_ (.A(_05121_),
    .B(_05348_),
    .Y(_05349_));
 sky130_fd_sc_hd__nand2_1 _12374_ (.A(net142),
    .B(_05349_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand2_1 _12375_ (.A(_05347_),
    .B(_05350_),
    .Y(_05351_));
 sky130_fd_sc_hd__or2_1 _12376_ (.A(_05347_),
    .B(_05350_),
    .X(_05353_));
 sky130_fd_sc_hd__a21oi_1 _12377_ (.A1(net137),
    .A2(_01995_),
    .B1(_02001_),
    .Y(_05354_));
 sky130_fd_sc_hd__a31o_1 _12378_ (.A1(net137),
    .A2(_01995_),
    .A3(_02001_),
    .B1(_02434_),
    .X(_05355_));
 sky130_fd_sc_hd__nor2_2 _12379_ (.A(_05354_),
    .B(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__a21o_1 _12380_ (.A1(_05623_),
    .A2(_05271_),
    .B1(_05602_),
    .X(_05357_));
 sky130_fd_sc_hd__mux2_1 _12381_ (.A0(_06607_),
    .A1(_05357_),
    .S(net283),
    .X(_05358_));
 sky130_fd_sc_hd__nand2_1 _12382_ (.A(_05526_),
    .B(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__o211a_1 _12383_ (.A1(_05526_),
    .A2(_05358_),
    .B1(_05359_),
    .C1(_02426_),
    .X(_05360_));
 sky130_fd_sc_hd__o21a_1 _12384_ (.A1(_05275_),
    .A2(_05279_),
    .B1(_05277_),
    .X(_05361_));
 sky130_fd_sc_hd__nor2_1 _12385_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05362_));
 sky130_fd_sc_hd__nand2_1 _12386_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05364_));
 sky130_fd_sc_hd__and2b_1 _12387_ (.A_N(_05362_),
    .B(_05364_),
    .X(_05365_));
 sky130_fd_sc_hd__xnor2_1 _12388_ (.A(_05361_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__mux2_1 _12389_ (.A0(_03509_),
    .A1(_05366_),
    .S(net245),
    .X(_05367_));
 sky130_fd_sc_hd__or2_1 _12390_ (.A(\div_shifter[55] ),
    .B(_05284_),
    .X(_05368_));
 sky130_fd_sc_hd__a21oi_1 _12391_ (.A1(net230),
    .A2(_05368_),
    .B1(\div_shifter[56] ),
    .Y(_05369_));
 sky130_fd_sc_hd__a31o_1 _12392_ (.A1(\div_shifter[56] ),
    .A2(net229),
    .A3(_05368_),
    .B1(net191),
    .X(_05370_));
 sky130_fd_sc_hd__or3_1 _12393_ (.A(\div_res[23] ),
    .B(\div_res[22] ),
    .C(_05191_),
    .X(_05371_));
 sky130_fd_sc_hd__a21oi_1 _12394_ (.A1(net142),
    .A2(_05371_),
    .B1(\div_res[24] ),
    .Y(_05372_));
 sky130_fd_sc_hd__a31o_1 _12395_ (.A1(\div_res[24] ),
    .A2(net142),
    .A3(_05371_),
    .B1(net190),
    .X(_05373_));
 sky130_fd_sc_hd__o22a_1 _12396_ (.A1(_05482_),
    .A2(net204),
    .B1(net231),
    .B2(reg1_val[24]),
    .X(_05375_));
 sky130_fd_sc_hd__o21ai_1 _12397_ (.A1(_05504_),
    .A2(_02440_),
    .B1(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__a221o_1 _12398_ (.A1(_05526_),
    .A2(net196),
    .B1(_02435_),
    .B2(_05515_),
    .C1(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__a31o_1 _12399_ (.A1(_00304_),
    .A2(_00328_),
    .A3(net256),
    .B1(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__a221o_1 _12400_ (.A1(_02424_),
    .A2(_03509_),
    .B1(_03516_),
    .B2(net171),
    .C1(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__o21ba_1 _12401_ (.A1(_05372_),
    .A2(_05373_),
    .B1_N(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__o21ai_1 _12402_ (.A1(_05369_),
    .A2(_05370_),
    .B1(_05380_),
    .Y(_05381_));
 sky130_fd_sc_hd__a211o_1 _12403_ (.A1(net205),
    .A2(_05367_),
    .B1(_05381_),
    .C1(_05360_),
    .X(_05382_));
 sky130_fd_sc_hd__a311o_1 _12404_ (.A1(_02348_),
    .A2(_05351_),
    .A3(_05353_),
    .B1(_05356_),
    .C1(_05382_),
    .X(_05383_));
 sky130_fd_sc_hd__and2_1 _12405_ (.A(curr_PC[24]),
    .B(_05297_),
    .X(_05384_));
 sky130_fd_sc_hd__o21ai_1 _12406_ (.A1(curr_PC[24]),
    .A2(_05297_),
    .B1(net243),
    .Y(_05386_));
 sky130_fd_sc_hd__a2bb2o_4 _12407_ (.A1_N(_05384_),
    .A2_N(_05386_),
    .B1(net240),
    .B2(_05383_),
    .X(dest_val[24]));
 sky130_fd_sc_hd__a22o_1 _12408_ (.A1(_00177_),
    .A2(net8),
    .B1(net3),
    .B2(_00136_),
    .X(_05387_));
 sky130_fd_sc_hd__xnor2_1 _12409_ (.A(net58),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__nand2_1 _12410_ (.A(_05302_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__or2_1 _12411_ (.A(_05302_),
    .B(_05388_),
    .X(_05390_));
 sky130_fd_sc_hd__nand2_1 _12412_ (.A(_05389_),
    .B(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(_00144_),
    .B(net61),
    .Y(_05392_));
 sky130_fd_sc_hd__xor2_1 _12414_ (.A(_05391_),
    .B(_05392_),
    .X(_05393_));
 sky130_fd_sc_hd__o21ai_1 _12415_ (.A1(_05302_),
    .A2(_05303_),
    .B1(_05305_),
    .Y(_05394_));
 sky130_fd_sc_hd__o22a_1 _12416_ (.A1(net35),
    .A2(net10),
    .B1(net5),
    .B2(_00321_),
    .X(_05396_));
 sky130_fd_sc_hd__xnor2_1 _12417_ (.A(net93),
    .B(_05396_),
    .Y(_05397_));
 sky130_fd_sc_hd__a22o_1 _12418_ (.A1(_00516_),
    .A2(net12),
    .B1(_00812_),
    .B2(net16),
    .X(_05398_));
 sky130_fd_sc_hd__xnor2_1 _12419_ (.A(net64),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__nand2_1 _12420_ (.A(_00309_),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__xnor2_1 _12421_ (.A(net92),
    .B(_05399_),
    .Y(_05401_));
 sky130_fd_sc_hd__nand2_1 _12422_ (.A(_05397_),
    .B(_05401_),
    .Y(_05402_));
 sky130_fd_sc_hd__or2_1 _12423_ (.A(_05397_),
    .B(_05401_),
    .X(_05403_));
 sky130_fd_sc_hd__nand2_1 _12424_ (.A(_05402_),
    .B(_05403_),
    .Y(_05404_));
 sky130_fd_sc_hd__a21oi_1 _12425_ (.A1(_05316_),
    .A2(_05321_),
    .B1(_05404_),
    .Y(_05405_));
 sky130_fd_sc_hd__and3_1 _12426_ (.A(_05316_),
    .B(_05321_),
    .C(_05404_),
    .X(_05407_));
 sky130_fd_sc_hd__or2_1 _12427_ (.A(_05405_),
    .B(_05407_),
    .X(_05408_));
 sky130_fd_sc_hd__and2b_1 _12428_ (.A_N(_05408_),
    .B(_05394_),
    .X(_05409_));
 sky130_fd_sc_hd__xnor2_1 _12429_ (.A(_05394_),
    .B(_05408_),
    .Y(_05410_));
 sky130_fd_sc_hd__nand2_1 _12430_ (.A(_05393_),
    .B(_05410_),
    .Y(_05411_));
 sky130_fd_sc_hd__or2_1 _12431_ (.A(_05393_),
    .B(_05410_),
    .X(_05412_));
 sky130_fd_sc_hd__nand2_1 _12432_ (.A(_05411_),
    .B(_05412_),
    .Y(_05413_));
 sky130_fd_sc_hd__a21bo_1 _12433_ (.A1(_05309_),
    .A2(_05325_),
    .B1_N(_05324_),
    .X(_05414_));
 sky130_fd_sc_hd__nand2b_1 _12434_ (.A_N(_05413_),
    .B(_05414_),
    .Y(_05415_));
 sky130_fd_sc_hd__xor2_1 _12435_ (.A(_05413_),
    .B(_05414_),
    .X(_05416_));
 sky130_fd_sc_hd__a21oi_1 _12436_ (.A1(_05328_),
    .A2(_05332_),
    .B1(_05416_),
    .Y(_05418_));
 sky130_fd_sc_hd__nand3_1 _12437_ (.A(_05328_),
    .B(_05332_),
    .C(_05416_),
    .Y(_05419_));
 sky130_fd_sc_hd__nand2b_2 _12438_ (.A_N(_05418_),
    .B(_05419_),
    .Y(_05420_));
 sky130_fd_sc_hd__nor2_1 _12439_ (.A(_05257_),
    .B(_05338_),
    .Y(_05421_));
 sky130_fd_sc_hd__and3_1 _12440_ (.A(_05075_),
    .B(_05165_),
    .C(_05421_),
    .X(_05422_));
 sky130_fd_sc_hd__a21oi_1 _12441_ (.A1(_05253_),
    .A2(_05336_),
    .B1(_05337_),
    .Y(_05423_));
 sky130_fd_sc_hd__or3_1 _12442_ (.A(_05257_),
    .B(_05260_),
    .C(_05338_),
    .X(_05424_));
 sky130_fd_sc_hd__nand2b_1 _12443_ (.A_N(_05423_),
    .B(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__a21o_1 _12444_ (.A1(_05078_),
    .A2(_05422_),
    .B1(_05425_),
    .X(_05426_));
 sky130_fd_sc_hd__a31o_1 _12445_ (.A1(_04692_),
    .A2(_05079_),
    .A3(_05422_),
    .B1(_05426_),
    .X(_05427_));
 sky130_fd_sc_hd__xor2_2 _12446_ (.A(_05420_),
    .B(_05427_),
    .X(_05429_));
 sky130_fd_sc_hd__a31o_1 _12447_ (.A1(_05121_),
    .A2(_05347_),
    .A3(_05348_),
    .B1(_06681_),
    .X(_05430_));
 sky130_fd_sc_hd__o21ai_1 _12448_ (.A1(_05429_),
    .A2(_05430_),
    .B1(_02348_),
    .Y(_05431_));
 sky130_fd_sc_hd__a21oi_1 _12449_ (.A1(_05429_),
    .A2(_05430_),
    .B1(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__a21o_1 _12450_ (.A1(_05526_),
    .A2(_05357_),
    .B1(_05515_),
    .X(_05433_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(_06625_),
    .A1(_05433_),
    .S(net283),
    .X(_05434_));
 sky130_fd_sc_hd__nand2_1 _12452_ (.A(_05352_),
    .B(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__o211a_1 _12453_ (.A1(_05352_),
    .A2(_05434_),
    .B1(_05435_),
    .C1(_02426_),
    .X(_05436_));
 sky130_fd_sc_hd__o21a_1 _12454_ (.A1(_01995_),
    .A2(_02001_),
    .B1(net137),
    .X(_05437_));
 sky130_fd_sc_hd__o21ai_2 _12455_ (.A1(_01923_),
    .A2(_05437_),
    .B1(_02433_),
    .Y(_05438_));
 sky130_fd_sc_hd__a21oi_4 _12456_ (.A1(_01923_),
    .A2(_05437_),
    .B1(_05438_),
    .Y(_05440_));
 sky130_fd_sc_hd__o21a_1 _12457_ (.A1(_05361_),
    .A2(_05362_),
    .B1(_05364_),
    .X(_05441_));
 sky130_fd_sc_hd__nor2_1 _12458_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05442_));
 sky130_fd_sc_hd__nand2_1 _12459_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05443_));
 sky130_fd_sc_hd__nand2b_1 _12460_ (.A_N(_05442_),
    .B(_05443_),
    .Y(_05444_));
 sky130_fd_sc_hd__xnor2_1 _12461_ (.A(_05441_),
    .B(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__nor2_1 _12462_ (.A(net245),
    .B(_03366_),
    .Y(_05446_));
 sky130_fd_sc_hd__a211o_1 _12463_ (.A1(net245),
    .A2(_05445_),
    .B1(_05446_),
    .C1(_06667_),
    .X(_05447_));
 sky130_fd_sc_hd__or2_1 _12464_ (.A(\div_shifter[56] ),
    .B(_05368_),
    .X(_05448_));
 sky130_fd_sc_hd__a21oi_1 _12465_ (.A1(net229),
    .A2(_05448_),
    .B1(\div_shifter[57] ),
    .Y(_05449_));
 sky130_fd_sc_hd__a311o_1 _12466_ (.A1(\div_shifter[57] ),
    .A2(net229),
    .A3(_05448_),
    .B1(_05449_),
    .C1(net191),
    .X(_05451_));
 sky130_fd_sc_hd__or2_1 _12467_ (.A(\div_res[24] ),
    .B(_05371_),
    .X(_05452_));
 sky130_fd_sc_hd__a21oi_1 _12468_ (.A1(net142),
    .A2(_05452_),
    .B1(\div_res[25] ),
    .Y(_05453_));
 sky130_fd_sc_hd__a311o_1 _12469_ (.A1(\div_res[25] ),
    .A2(net142),
    .A3(_05452_),
    .B1(_05453_),
    .C1(net190),
    .X(_05454_));
 sky130_fd_sc_hd__o21ai_1 _12470_ (.A1(reg1_val[25]),
    .A2(_05308_),
    .B1(_02439_),
    .Y(_05455_));
 sky130_fd_sc_hd__o221ai_1 _12471_ (.A1(_05319_),
    .A2(net204),
    .B1(net231),
    .B2(reg1_val[25]),
    .C1(_05455_),
    .Y(_05456_));
 sky130_fd_sc_hd__a221o_1 _12472_ (.A1(_05352_),
    .A2(net196),
    .B1(_02435_),
    .B2(_05341_),
    .C1(_05456_),
    .X(_05457_));
 sky130_fd_sc_hd__a221o_1 _12473_ (.A1(_02424_),
    .A2(_03366_),
    .B1(_03372_),
    .B2(net171),
    .C1(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__a21oi_1 _12474_ (.A1(_00306_),
    .A2(net257),
    .B1(_05458_),
    .Y(_05459_));
 sky130_fd_sc_hd__and4_1 _12475_ (.A(_05447_),
    .B(_05451_),
    .C(_05454_),
    .D(_05459_),
    .X(_05460_));
 sky130_fd_sc_hd__or4b_1 _12476_ (.A(_05432_),
    .B(_05436_),
    .C(_05440_),
    .D_N(_05460_),
    .X(_05462_));
 sky130_fd_sc_hd__and3_1 _12477_ (.A(curr_PC[24]),
    .B(curr_PC[25]),
    .C(_05297_),
    .X(_05463_));
 sky130_fd_sc_hd__o21ai_1 _12478_ (.A1(curr_PC[25]),
    .A2(_05384_),
    .B1(_06652_),
    .Y(_05464_));
 sky130_fd_sc_hd__a2bb2o_4 _12479_ (.A1_N(_05463_),
    .A2_N(_05464_),
    .B1(net240),
    .B2(_05462_),
    .X(dest_val[25]));
 sky130_fd_sc_hd__nand2_1 _12480_ (.A(_05347_),
    .B(_05429_),
    .Y(_05465_));
 sky130_fd_sc_hd__o21a_1 _12481_ (.A1(_05349_),
    .A2(_05465_),
    .B1(net143),
    .X(_05466_));
 sky130_fd_sc_hd__o21ai_2 _12482_ (.A1(_05391_),
    .A2(_05392_),
    .B1(_05389_),
    .Y(_05467_));
 sky130_fd_sc_hd__a22o_1 _12483_ (.A1(net12),
    .A2(_00812_),
    .B1(_02065_),
    .B2(net16),
    .X(_05468_));
 sky130_fd_sc_hd__xnor2_1 _12484_ (.A(net64),
    .B(_05468_),
    .Y(_05469_));
 sky130_fd_sc_hd__or2_1 _12485_ (.A(_00314_),
    .B(net5),
    .X(_05470_));
 sky130_fd_sc_hd__a22o_1 _12486_ (.A1(_00316_),
    .A2(net7),
    .B1(_05470_),
    .B2(net93),
    .X(_05472_));
 sky130_fd_sc_hd__nor2_1 _12487_ (.A(_05469_),
    .B(_05472_),
    .Y(_05473_));
 sky130_fd_sc_hd__and2_1 _12488_ (.A(_05469_),
    .B(_05472_),
    .X(_05474_));
 sky130_fd_sc_hd__nor2_1 _12489_ (.A(_05473_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__a21oi_1 _12490_ (.A1(_05400_),
    .A2(_05402_),
    .B1(_05475_),
    .Y(_05476_));
 sky130_fd_sc_hd__and3_1 _12491_ (.A(_05400_),
    .B(_05402_),
    .C(_05475_),
    .X(_05477_));
 sky130_fd_sc_hd__nor2_1 _12492_ (.A(_05476_),
    .B(_05477_),
    .Y(_05478_));
 sky130_fd_sc_hd__and2_1 _12493_ (.A(_05467_),
    .B(_05478_),
    .X(_05479_));
 sky130_fd_sc_hd__xnor2_1 _12494_ (.A(_05467_),
    .B(_05478_),
    .Y(_05480_));
 sky130_fd_sc_hd__a22o_1 _12495_ (.A1(_00516_),
    .A2(net8),
    .B1(net3),
    .B2(_00177_),
    .X(_05481_));
 sky130_fd_sc_hd__nor2_1 _12496_ (.A(_00136_),
    .B(net58),
    .Y(_05483_));
 sky130_fd_sc_hd__xnor2_1 _12497_ (.A(_05481_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__nor2_1 _12498_ (.A(_05480_),
    .B(_05484_),
    .Y(_05485_));
 sky130_fd_sc_hd__and2_1 _12499_ (.A(_05480_),
    .B(_05484_),
    .X(_05486_));
 sky130_fd_sc_hd__nor2_1 _12500_ (.A(_05485_),
    .B(_05486_),
    .Y(_05487_));
 sky130_fd_sc_hd__o21a_1 _12501_ (.A1(_05405_),
    .A2(_05409_),
    .B1(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__nor3_1 _12502_ (.A(_05405_),
    .B(_05409_),
    .C(_05487_),
    .Y(_05489_));
 sky130_fd_sc_hd__or2_1 _12503_ (.A(_05488_),
    .B(_05489_),
    .X(_05490_));
 sky130_fd_sc_hd__a21oi_1 _12504_ (.A1(_05411_),
    .A2(_05415_),
    .B1(_05490_),
    .Y(_05491_));
 sky130_fd_sc_hd__and3_1 _12505_ (.A(_05411_),
    .B(_05415_),
    .C(_05490_),
    .X(_05492_));
 sky130_fd_sc_hd__or2_2 _12506_ (.A(_05491_),
    .B(_05492_),
    .X(_05494_));
 sky130_fd_sc_hd__o21ai_1 _12507_ (.A1(_05335_),
    .A2(_05418_),
    .B1(_05419_),
    .Y(_05495_));
 sky130_fd_sc_hd__or2_1 _12508_ (.A(_05338_),
    .B(_05420_),
    .X(_05496_));
 sky130_fd_sc_hd__o21a_1 _12509_ (.A1(_05339_),
    .A2(_05496_),
    .B1(_05495_),
    .X(_05497_));
 sky130_fd_sc_hd__o31a_1 _12510_ (.A1(_05171_),
    .A2(_05340_),
    .A3(_05496_),
    .B1(_05497_),
    .X(_05498_));
 sky130_fd_sc_hd__xor2_2 _12511_ (.A(_05494_),
    .B(_05498_),
    .X(_05499_));
 sky130_fd_sc_hd__and2_1 _12512_ (.A(_05466_),
    .B(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__nor2_1 _12513_ (.A(_05466_),
    .B(_05499_),
    .Y(_05501_));
 sky130_fd_sc_hd__a21oi_1 _12514_ (.A1(_05352_),
    .A2(_05433_),
    .B1(_05341_),
    .Y(_05502_));
 sky130_fd_sc_hd__mux2_1 _12515_ (.A0(_06627_),
    .A1(_05502_),
    .S(net283),
    .X(_05503_));
 sky130_fd_sc_hd__nor2_1 _12516_ (.A(_05450_),
    .B(_05503_),
    .Y(_05505_));
 sky130_fd_sc_hd__a211o_1 _12517_ (.A1(_05450_),
    .A2(_05503_),
    .B1(_05505_),
    .C1(_02427_),
    .X(_05506_));
 sky130_fd_sc_hd__a21oi_2 _12518_ (.A1(net137),
    .A2(_02002_),
    .B1(_02007_),
    .Y(_05507_));
 sky130_fd_sc_hd__a31o_1 _12519_ (.A1(net137),
    .A2(_02002_),
    .A3(_02007_),
    .B1(_02434_),
    .X(_05508_));
 sky130_fd_sc_hd__o21a_1 _12520_ (.A1(_05441_),
    .A2(_05442_),
    .B1(_05443_),
    .X(_05509_));
 sky130_fd_sc_hd__nor2_1 _12521_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05510_));
 sky130_fd_sc_hd__nand2_1 _12522_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05511_));
 sky130_fd_sc_hd__nand2b_1 _12523_ (.A_N(_05510_),
    .B(_05511_),
    .Y(_05512_));
 sky130_fd_sc_hd__xnor2_1 _12524_ (.A(_05509_),
    .B(_05512_),
    .Y(_05513_));
 sky130_fd_sc_hd__nor2_1 _12525_ (.A(net244),
    .B(_03229_),
    .Y(_05514_));
 sky130_fd_sc_hd__a211o_1 _12526_ (.A1(net244),
    .A2(_05513_),
    .B1(_05514_),
    .C1(_06667_),
    .X(_05516_));
 sky130_fd_sc_hd__or2_1 _12527_ (.A(\div_shifter[57] ),
    .B(_05448_),
    .X(_05517_));
 sky130_fd_sc_hd__a21oi_1 _12528_ (.A1(net229),
    .A2(_05517_),
    .B1(\div_shifter[58] ),
    .Y(_05518_));
 sky130_fd_sc_hd__a311o_1 _12529_ (.A1(\div_shifter[58] ),
    .A2(net229),
    .A3(_05517_),
    .B1(_05518_),
    .C1(net191),
    .X(_05519_));
 sky130_fd_sc_hd__nor2_1 _12530_ (.A(\div_res[25] ),
    .B(_05452_),
    .Y(_05520_));
 sky130_fd_sc_hd__inv_2 _12531_ (.A(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__a21oi_1 _12532_ (.A1(net142),
    .A2(_05521_),
    .B1(\div_res[26] ),
    .Y(_05522_));
 sky130_fd_sc_hd__a31o_1 _12533_ (.A1(\div_res[26] ),
    .A2(net142),
    .A3(_05521_),
    .B1(net189),
    .X(_05523_));
 sky130_fd_sc_hd__and3_1 _12534_ (.A(_00298_),
    .B(_00310_),
    .C(net257),
    .X(_05524_));
 sky130_fd_sc_hd__a2bb2o_1 _12535_ (.A1_N(reg1_val[26]),
    .A2_N(net232),
    .B1(_05395_),
    .B2(_06677_),
    .X(_05525_));
 sky130_fd_sc_hd__a221o_1 _12536_ (.A1(_05417_),
    .A2(_02435_),
    .B1(_02439_),
    .B2(_05428_),
    .C1(_05525_),
    .X(_05527_));
 sky130_fd_sc_hd__a221o_1 _12537_ (.A1(_05439_),
    .A2(net195),
    .B1(_03229_),
    .B2(net167),
    .C1(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__a211oi_1 _12538_ (.A1(net171),
    .A2(_03235_),
    .B1(_05524_),
    .C1(_05528_),
    .Y(_05529_));
 sky130_fd_sc_hd__o211a_1 _12539_ (.A1(_05522_),
    .A2(_05523_),
    .B1(_05529_),
    .C1(_05519_),
    .X(_05530_));
 sky130_fd_sc_hd__o211a_1 _12540_ (.A1(_05507_),
    .A2(_05508_),
    .B1(_05516_),
    .C1(_05530_),
    .X(_05531_));
 sky130_fd_sc_hd__o311a_1 _12541_ (.A1(_02349_),
    .A2(_05500_),
    .A3(_05501_),
    .B1(_05506_),
    .C1(_05531_),
    .X(_05532_));
 sky130_fd_sc_hd__nor2_1 _12542_ (.A(curr_PC[26]),
    .B(_05463_),
    .Y(_05533_));
 sky130_fd_sc_hd__nand2_1 _12543_ (.A(curr_PC[26]),
    .B(_05463_),
    .Y(_05534_));
 sky130_fd_sc_hd__or3b_1 _12544_ (.A(net240),
    .B(_05533_),
    .C_N(_05534_),
    .X(_05535_));
 sky130_fd_sc_hd__o21ai_4 _12545_ (.A1(_06652_),
    .A2(_05532_),
    .B1(_05535_),
    .Y(dest_val[26]));
 sky130_fd_sc_hd__nor2_1 _12546_ (.A(curr_PC[27]),
    .B(_05534_),
    .Y(_05537_));
 sky130_fd_sc_hd__a21o_1 _12547_ (.A1(curr_PC[27]),
    .A2(_05534_),
    .B1(net240),
    .X(_05538_));
 sky130_fd_sc_hd__a22o_1 _12548_ (.A1(_00812_),
    .A2(net8),
    .B1(net3),
    .B2(_00516_),
    .X(_05539_));
 sky130_fd_sc_hd__xnor2_1 _12549_ (.A(net58),
    .B(_05539_),
    .Y(_05540_));
 sky130_fd_sc_hd__and2_1 _12550_ (.A(_00302_),
    .B(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__nor2_1 _12551_ (.A(_00302_),
    .B(_05540_),
    .Y(_05542_));
 sky130_fd_sc_hd__nor2_1 _12552_ (.A(_05541_),
    .B(_05542_),
    .Y(_05543_));
 sky130_fd_sc_hd__a22o_1 _12553_ (.A1(net12),
    .A2(_02065_),
    .B1(net7),
    .B2(net16),
    .X(_05544_));
 sky130_fd_sc_hd__xnor2_1 _12554_ (.A(net64),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__xnor2_1 _12555_ (.A(_05543_),
    .B(_05545_),
    .Y(_05546_));
 sky130_fd_sc_hd__o21ai_1 _12556_ (.A1(net52),
    .A2(_05481_),
    .B1(net43),
    .Y(_05548_));
 sky130_fd_sc_hd__or4_1 _12557_ (.A(net52),
    .B(net43),
    .C(net58),
    .D(_05481_),
    .X(_05549_));
 sky130_fd_sc_hd__nand2_1 _12558_ (.A(_05548_),
    .B(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__nor2_1 _12559_ (.A(net58),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__xor2_1 _12560_ (.A(_05473_),
    .B(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__nor2_1 _12561_ (.A(_05546_),
    .B(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__and2_1 _12562_ (.A(_05546_),
    .B(_05552_),
    .X(_05554_));
 sky130_fd_sc_hd__nor2_1 _12563_ (.A(_05553_),
    .B(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__o21a_1 _12564_ (.A1(_05476_),
    .A2(_05479_),
    .B1(_05555_),
    .X(_05556_));
 sky130_fd_sc_hd__nor3_1 _12565_ (.A(_05476_),
    .B(_05479_),
    .C(_05555_),
    .Y(_05557_));
 sky130_fd_sc_hd__nor2_1 _12566_ (.A(_05556_),
    .B(_05557_),
    .Y(_05559_));
 sky130_fd_sc_hd__o21a_1 _12567_ (.A1(_05485_),
    .A2(_05488_),
    .B1(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__or3_1 _12568_ (.A(_05485_),
    .B(_05488_),
    .C(_05559_),
    .X(_05561_));
 sky130_fd_sc_hd__nand2b_2 _12569_ (.A_N(_05560_),
    .B(_05561_),
    .Y(_05562_));
 sky130_fd_sc_hd__nor2_1 _12570_ (.A(_05420_),
    .B(_05494_),
    .Y(_05563_));
 sky130_fd_sc_hd__o21ba_1 _12571_ (.A1(_05418_),
    .A2(_05491_),
    .B1_N(_05492_),
    .X(_05564_));
 sky130_fd_sc_hd__a21o_1 _12572_ (.A1(_05423_),
    .A2(_05563_),
    .B1(_05564_),
    .X(_05565_));
 sky130_fd_sc_hd__a31o_1 _12573_ (.A1(_05263_),
    .A2(_05421_),
    .A3(_05563_),
    .B1(_05565_),
    .X(_05566_));
 sky130_fd_sc_hd__xnor2_2 _12574_ (.A(_05562_),
    .B(_05566_),
    .Y(_05567_));
 sky130_fd_sc_hd__o31a_1 _12575_ (.A1(_05349_),
    .A2(_05465_),
    .A3(_05499_),
    .B1(net143),
    .X(_05568_));
 sky130_fd_sc_hd__a21oi_1 _12576_ (.A1(_05567_),
    .A2(_05568_),
    .B1(_02349_),
    .Y(_05570_));
 sky130_fd_sc_hd__o21a_1 _12577_ (.A1(_05567_),
    .A2(_05568_),
    .B1(_05570_),
    .X(_05571_));
 sky130_fd_sc_hd__and3_1 _12578_ (.A(net296),
    .B(_06612_),
    .C(_06628_),
    .X(_05572_));
 sky130_fd_sc_hd__o21ai_1 _12579_ (.A1(_05450_),
    .A2(_05502_),
    .B1(_05406_),
    .Y(_05573_));
 sky130_fd_sc_hd__a21o_1 _12580_ (.A1(net284),
    .A2(_05573_),
    .B1(_05572_),
    .X(_05574_));
 sky130_fd_sc_hd__nand2_1 _12581_ (.A(_05036_),
    .B(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hd__o211a_1 _12582_ (.A1(_05036_),
    .A2(_05574_),
    .B1(_05575_),
    .C1(_02426_),
    .X(_05576_));
 sky130_fd_sc_hd__nand2_1 _12583_ (.A(net138),
    .B(_02008_),
    .Y(_05577_));
 sky130_fd_sc_hd__xnor2_1 _12584_ (.A(_02009_),
    .B(_05577_),
    .Y(_05578_));
 sky130_fd_sc_hd__o21a_1 _12585_ (.A1(_05509_),
    .A2(_05510_),
    .B1(_05511_),
    .X(_05579_));
 sky130_fd_sc_hd__nor2_1 _12586_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05581_));
 sky130_fd_sc_hd__nand2_1 _12587_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05582_));
 sky130_fd_sc_hd__and2b_1 _12588_ (.A_N(_05581_),
    .B(_05582_),
    .X(_05583_));
 sky130_fd_sc_hd__or2_1 _12589_ (.A(_05579_),
    .B(_05583_),
    .X(_05584_));
 sky130_fd_sc_hd__a21oi_1 _12590_ (.A1(_05579_),
    .A2(_05583_),
    .B1(net224),
    .Y(_05585_));
 sky130_fd_sc_hd__a22o_1 _12591_ (.A1(net224),
    .A2(_03109_),
    .B1(_05584_),
    .B2(_05585_),
    .X(_05586_));
 sky130_fd_sc_hd__or2_1 _12592_ (.A(\div_res[26] ),
    .B(_05521_),
    .X(_05587_));
 sky130_fd_sc_hd__a21oi_1 _12593_ (.A1(net142),
    .A2(_05587_),
    .B1(\div_res[27] ),
    .Y(_05588_));
 sky130_fd_sc_hd__a31o_1 _12594_ (.A1(\div_res[27] ),
    .A2(net142),
    .A3(_05587_),
    .B1(net190),
    .X(_05589_));
 sky130_fd_sc_hd__or2_1 _12595_ (.A(\div_shifter[58] ),
    .B(_05517_),
    .X(_05590_));
 sky130_fd_sc_hd__a21oi_1 _12596_ (.A1(net229),
    .A2(_05590_),
    .B1(\div_shifter[59] ),
    .Y(_05592_));
 sky130_fd_sc_hd__a311o_1 _12597_ (.A1(\div_shifter[59] ),
    .A2(net229),
    .A3(_05590_),
    .B1(_05592_),
    .C1(net191),
    .X(_05593_));
 sky130_fd_sc_hd__or3_1 _12598_ (.A(_00296_),
    .B(_00299_),
    .C(_02432_),
    .X(_05594_));
 sky130_fd_sc_hd__a21oi_1 _12599_ (.A1(_05025_),
    .A2(net196),
    .B1(_02439_),
    .Y(_05595_));
 sky130_fd_sc_hd__o221a_1 _12600_ (.A1(_04982_),
    .A2(net204),
    .B1(net231),
    .B2(reg1_val[27]),
    .C1(net240),
    .X(_05596_));
 sky130_fd_sc_hd__o221a_1 _12601_ (.A1(_05025_),
    .A2(_02436_),
    .B1(_05595_),
    .B2(_05004_),
    .C1(_05596_),
    .X(_05597_));
 sky130_fd_sc_hd__o221a_1 _12602_ (.A1(net169),
    .A2(_03096_),
    .B1(_03109_),
    .B2(_02425_),
    .C1(_05597_),
    .X(_05598_));
 sky130_fd_sc_hd__o211a_1 _12603_ (.A1(_05588_),
    .A2(_05589_),
    .B1(_05594_),
    .C1(_05598_),
    .X(_05599_));
 sky130_fd_sc_hd__o211a_1 _12604_ (.A1(_06667_),
    .A2(_05586_),
    .B1(_05593_),
    .C1(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__o21ai_1 _12605_ (.A1(_02434_),
    .A2(_05578_),
    .B1(_05600_),
    .Y(_05601_));
 sky130_fd_sc_hd__o32a_4 _12606_ (.A1(_05571_),
    .A2(_05576_),
    .A3(_05601_),
    .B1(_05538_),
    .B2(_05537_),
    .X(dest_val[27]));
 sky130_fd_sc_hd__o31a_1 _12607_ (.A1(net58),
    .A2(_05473_),
    .A3(_05550_),
    .B1(_05549_),
    .X(_05603_));
 sky130_fd_sc_hd__a21o_1 _12608_ (.A1(_05543_),
    .A2(_05545_),
    .B1(_05541_),
    .X(_05604_));
 sky130_fd_sc_hd__a22o_1 _12609_ (.A1(_02065_),
    .A2(net8),
    .B1(net3),
    .B2(_00812_),
    .X(_05605_));
 sky130_fd_sc_hd__xnor2_1 _12610_ (.A(net58),
    .B(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__and2_1 _12611_ (.A(_05604_),
    .B(_05606_),
    .X(_05607_));
 sky130_fd_sc_hd__or2_1 _12612_ (.A(_05604_),
    .B(_05606_),
    .X(_05608_));
 sky130_fd_sc_hd__and2b_1 _12613_ (.A_N(_05607_),
    .B(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__and3_1 _12614_ (.A(_00516_),
    .B(net61),
    .C(_05609_),
    .X(_05610_));
 sky130_fd_sc_hd__a21oi_1 _12615_ (.A1(_00516_),
    .A2(net61),
    .B1(_05609_),
    .Y(_05611_));
 sky130_fd_sc_hd__or2_1 _12616_ (.A(_05610_),
    .B(_05611_),
    .X(_05613_));
 sky130_fd_sc_hd__nand2_1 _12617_ (.A(_00559_),
    .B(net7),
    .Y(_05614_));
 sky130_fd_sc_hd__a22o_1 _12618_ (.A1(_00796_),
    .A2(net7),
    .B1(_05614_),
    .B2(_00787_),
    .X(_05615_));
 sky130_fd_sc_hd__nor2_1 _12619_ (.A(_05613_),
    .B(_05615_),
    .Y(_05616_));
 sky130_fd_sc_hd__and2_1 _12620_ (.A(_05613_),
    .B(_05615_),
    .X(_05617_));
 sky130_fd_sc_hd__nor3_1 _12621_ (.A(_05603_),
    .B(_05616_),
    .C(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__o21a_1 _12622_ (.A1(_05616_),
    .A2(_05617_),
    .B1(_05603_),
    .X(_05619_));
 sky130_fd_sc_hd__nor2_1 _12623_ (.A(_05618_),
    .B(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__o21a_1 _12624_ (.A1(_05553_),
    .A2(_05556_),
    .B1(_05620_),
    .X(_05621_));
 sky130_fd_sc_hd__nor3_1 _12625_ (.A(_05553_),
    .B(_05556_),
    .C(_05620_),
    .Y(_05622_));
 sky130_fd_sc_hd__or2_2 _12626_ (.A(_05621_),
    .B(_05622_),
    .X(_05624_));
 sky130_fd_sc_hd__or2_1 _12627_ (.A(_05494_),
    .B(_05562_),
    .X(_05625_));
 sky130_fd_sc_hd__o21ai_1 _12628_ (.A1(_05491_),
    .A2(_05560_),
    .B1(_05561_),
    .Y(_05626_));
 sky130_fd_sc_hd__nand2b_1 _12629_ (.A_N(_05496_),
    .B(_05342_),
    .Y(_05627_));
 sky130_fd_sc_hd__a21o_1 _12630_ (.A1(_05495_),
    .A2(_05627_),
    .B1(_05625_),
    .X(_05628_));
 sky130_fd_sc_hd__o311a_1 _12631_ (.A1(_05344_),
    .A2(_05496_),
    .A3(_05625_),
    .B1(_05626_),
    .C1(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__xor2_2 _12632_ (.A(_05624_),
    .B(_05629_),
    .X(_05630_));
 sky130_fd_sc_hd__inv_2 _12633_ (.A(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__or2_1 _12634_ (.A(_05499_),
    .B(_05567_),
    .X(_05632_));
 sky130_fd_sc_hd__nor3_1 _12635_ (.A(_05465_),
    .B(_05499_),
    .C(_05567_),
    .Y(_05633_));
 sky130_fd_sc_hd__a31o_1 _12636_ (.A1(_05121_),
    .A2(_05348_),
    .A3(_05633_),
    .B1(_06681_),
    .X(_05635_));
 sky130_fd_sc_hd__o21ai_1 _12637_ (.A1(_05631_),
    .A2(_05635_),
    .B1(_02348_),
    .Y(_05636_));
 sky130_fd_sc_hd__a21o_1 _12638_ (.A1(_05631_),
    .A2(_05635_),
    .B1(_05636_),
    .X(_05637_));
 sky130_fd_sc_hd__a21o_1 _12639_ (.A1(_05025_),
    .A2(_05406_),
    .B1(_05004_),
    .X(_05638_));
 sky130_fd_sc_hd__o41a_1 _12640_ (.A1(_05004_),
    .A2(_05015_),
    .A3(_05450_),
    .A4(_05502_),
    .B1(_05638_),
    .X(_05639_));
 sky130_fd_sc_hd__mux2_1 _12641_ (.A0(_06630_),
    .A1(_05639_),
    .S(net284),
    .X(_05640_));
 sky130_fd_sc_hd__nor2_1 _12642_ (.A(_05276_),
    .B(_05640_),
    .Y(_05641_));
 sky130_fd_sc_hd__a211o_1 _12643_ (.A1(_05276_),
    .A2(_05640_),
    .B1(_05641_),
    .C1(_02427_),
    .X(_05642_));
 sky130_fd_sc_hd__o211a_1 _12644_ (.A1(_02014_),
    .A2(_02015_),
    .B1(net138),
    .C1(_02010_),
    .X(_05643_));
 sky130_fd_sc_hd__a211oi_1 _12645_ (.A1(net138),
    .A2(_02010_),
    .B1(_02014_),
    .C1(_02015_),
    .Y(_05644_));
 sky130_fd_sc_hd__o21ai_2 _12646_ (.A1(_05579_),
    .A2(_05581_),
    .B1(_05582_),
    .Y(_05646_));
 sky130_fd_sc_hd__xnor2_1 _12647_ (.A(_04587_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__nor2_1 _12648_ (.A(net223),
    .B(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__a211o_1 _12649_ (.A1(net223),
    .A2(_02938_),
    .B1(_05648_),
    .C1(_06667_),
    .X(_05649_));
 sky130_fd_sc_hd__or2_1 _12650_ (.A(\div_res[27] ),
    .B(_05587_),
    .X(_05650_));
 sky130_fd_sc_hd__a21oi_1 _12651_ (.A1(net143),
    .A2(_05650_),
    .B1(\div_res[28] ),
    .Y(_05651_));
 sky130_fd_sc_hd__a311o_1 _12652_ (.A1(\div_res[28] ),
    .A2(net143),
    .A3(_05650_),
    .B1(_05651_),
    .C1(net190),
    .X(_05652_));
 sky130_fd_sc_hd__or2_1 _12653_ (.A(\div_shifter[59] ),
    .B(_05590_),
    .X(_05653_));
 sky130_fd_sc_hd__a21oi_1 _12654_ (.A1(net229),
    .A2(_05653_),
    .B1(\div_shifter[60] ),
    .Y(_05654_));
 sky130_fd_sc_hd__a311o_1 _12655_ (.A1(\div_shifter[60] ),
    .A2(net229),
    .A3(_05653_),
    .B1(_05654_),
    .C1(net191),
    .X(_05655_));
 sky130_fd_sc_hd__and3_1 _12656_ (.A(_00554_),
    .B(_00555_),
    .C(net257),
    .X(_05657_));
 sky130_fd_sc_hd__o221a_1 _12657_ (.A1(_05254_),
    .A2(_02436_),
    .B1(net231),
    .B2(reg1_val[28]),
    .C1(net204),
    .X(_05658_));
 sky130_fd_sc_hd__o21ai_1 _12658_ (.A1(_05243_),
    .A2(_02440_),
    .B1(_05658_),
    .Y(_05659_));
 sky130_fd_sc_hd__a221o_1 _12659_ (.A1(_05265_),
    .A2(net196),
    .B1(_02939_),
    .B2(_02424_),
    .C1(_05659_),
    .X(_05660_));
 sky130_fd_sc_hd__a211o_1 _12660_ (.A1(net171),
    .A2(_02927_),
    .B1(_05657_),
    .C1(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__and4b_1 _12661_ (.A_N(_05661_),
    .B(_05655_),
    .C(_05652_),
    .D(_05649_),
    .X(_05662_));
 sky130_fd_sc_hd__o31a_1 _12662_ (.A1(_02434_),
    .A2(_05643_),
    .A3(_05644_),
    .B1(_05662_),
    .X(_05663_));
 sky130_fd_sc_hd__a21o_1 _12663_ (.A1(_05211_),
    .A2(_06677_),
    .B1(_06652_),
    .X(_05664_));
 sky130_fd_sc_hd__a31oi_4 _12664_ (.A1(_05637_),
    .A2(_05642_),
    .A3(_05663_),
    .B1(_05664_),
    .Y(dest_val[28]));
 sky130_fd_sc_hd__a22o_1 _12665_ (.A1(net8),
    .A2(net7),
    .B1(net3),
    .B2(_02065_),
    .X(_05665_));
 sky130_fd_sc_hd__xnor2_1 _12666_ (.A(net58),
    .B(_05665_),
    .Y(_05667_));
 sky130_fd_sc_hd__nand2_1 _12667_ (.A(_00812_),
    .B(net61),
    .Y(_05668_));
 sky130_fd_sc_hd__xnor2_1 _12668_ (.A(net64),
    .B(_05668_),
    .Y(_05669_));
 sky130_fd_sc_hd__nand2_1 _12669_ (.A(_05667_),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__or2_1 _12670_ (.A(_05667_),
    .B(_05669_),
    .X(_05671_));
 sky130_fd_sc_hd__and3_1 _12671_ (.A(_05615_),
    .B(_05670_),
    .C(_05671_),
    .X(_05672_));
 sky130_fd_sc_hd__a21oi_1 _12672_ (.A1(_05670_),
    .A2(_05671_),
    .B1(_05615_),
    .Y(_05673_));
 sky130_fd_sc_hd__nor2_1 _12673_ (.A(_05672_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__o21a_1 _12674_ (.A1(_05607_),
    .A2(_05610_),
    .B1(_05674_),
    .X(_05675_));
 sky130_fd_sc_hd__nor3_1 _12675_ (.A(_05607_),
    .B(_05610_),
    .C(_05674_),
    .Y(_05676_));
 sky130_fd_sc_hd__nor2_1 _12676_ (.A(_05675_),
    .B(_05676_),
    .Y(_05678_));
 sky130_fd_sc_hd__or3_1 _12677_ (.A(_05616_),
    .B(_05618_),
    .C(_05678_),
    .X(_05679_));
 sky130_fd_sc_hd__o21a_1 _12678_ (.A1(_05616_),
    .A2(_05618_),
    .B1(_05678_),
    .X(_05680_));
 sky130_fd_sc_hd__o21ai_1 _12679_ (.A1(_05616_),
    .A2(_05618_),
    .B1(_05678_),
    .Y(_05681_));
 sky130_fd_sc_hd__nand2_2 _12680_ (.A(_05679_),
    .B(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__nor2_1 _12681_ (.A(_05562_),
    .B(_05624_),
    .Y(_05683_));
 sky130_fd_sc_hd__and4b_1 _12682_ (.A_N(_05081_),
    .B(_05422_),
    .C(_05563_),
    .D(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__o21ba_1 _12683_ (.A1(_05560_),
    .A2(_05621_),
    .B1_N(_05622_),
    .X(_05685_));
 sky130_fd_sc_hd__a21o_1 _12684_ (.A1(_05564_),
    .A2(_05683_),
    .B1(_05685_),
    .X(_05686_));
 sky130_fd_sc_hd__a31o_1 _12685_ (.A1(_05425_),
    .A2(_05563_),
    .A3(_05683_),
    .B1(_05686_),
    .X(_05687_));
 sky130_fd_sc_hd__nor2_1 _12686_ (.A(_05684_),
    .B(_05687_),
    .Y(_05689_));
 sky130_fd_sc_hd__xor2_2 _12687_ (.A(_05682_),
    .B(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__o41a_1 _12688_ (.A1(_05349_),
    .A2(_05465_),
    .A3(_05630_),
    .A4(_05632_),
    .B1(net143),
    .X(_05691_));
 sky130_fd_sc_hd__o21ai_1 _12689_ (.A1(_05690_),
    .A2(_05691_),
    .B1(_02348_),
    .Y(_05692_));
 sky130_fd_sc_hd__a21oi_1 _12690_ (.A1(_05690_),
    .A2(_05691_),
    .B1(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_1 _12691_ (.A1(_05243_),
    .A2(_05639_),
    .B1(_05254_),
    .Y(_05694_));
 sky130_fd_sc_hd__mux2_1 _12692_ (.A0(_06631_),
    .A1(_05694_),
    .S(net284),
    .X(_05695_));
 sky130_fd_sc_hd__nand2_1 _12693_ (.A(_05178_),
    .B(_05695_),
    .Y(_05696_));
 sky130_fd_sc_hd__o211a_1 _12694_ (.A1(_05178_),
    .A2(_05695_),
    .B1(_05696_),
    .C1(_02426_),
    .X(_05697_));
 sky130_fd_sc_hd__and2_1 _12695_ (.A(net138),
    .B(_02017_),
    .X(_05698_));
 sky130_fd_sc_hd__o21ai_1 _12696_ (.A1(_01922_),
    .A2(_05698_),
    .B1(net233),
    .Y(_05700_));
 sky130_fd_sc_hd__a21oi_2 _12697_ (.A1(_01922_),
    .A2(_05698_),
    .B1(_05700_),
    .Y(_05701_));
 sky130_fd_sc_hd__and3_1 _12698_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_05646_),
    .X(_05702_));
 sky130_fd_sc_hd__a21oi_1 _12699_ (.A1(reg1_val[28]),
    .A2(_05646_),
    .B1(reg1_val[29]),
    .Y(_05703_));
 sky130_fd_sc_hd__o21a_1 _12700_ (.A1(_05702_),
    .A2(_05703_),
    .B1(net245),
    .X(_05704_));
 sky130_fd_sc_hd__a211o_1 _12701_ (.A1(net223),
    .A2(_02755_),
    .B1(_05704_),
    .C1(_06667_),
    .X(_05705_));
 sky130_fd_sc_hd__or2_1 _12702_ (.A(\div_shifter[60] ),
    .B(_05653_),
    .X(_05706_));
 sky130_fd_sc_hd__a21oi_1 _12703_ (.A1(net229),
    .A2(_05706_),
    .B1(\div_shifter[61] ),
    .Y(_05707_));
 sky130_fd_sc_hd__a31o_1 _12704_ (.A1(\div_shifter[61] ),
    .A2(net229),
    .A3(_05706_),
    .B1(net191),
    .X(_05708_));
 sky130_fd_sc_hd__or2_1 _12705_ (.A(\div_res[28] ),
    .B(_05650_),
    .X(_05709_));
 sky130_fd_sc_hd__a21oi_1 _12706_ (.A1(net142),
    .A2(_05709_),
    .B1(\div_res[29] ),
    .Y(_05711_));
 sky130_fd_sc_hd__a31o_1 _12707_ (.A1(\div_res[29] ),
    .A2(net142),
    .A3(_05709_),
    .B1(net190),
    .X(_05712_));
 sky130_fd_sc_hd__o221ai_1 _12708_ (.A1(_05145_),
    .A2(_02440_),
    .B1(net232),
    .B2(reg1_val[29]),
    .C1(net204),
    .Y(_05713_));
 sky130_fd_sc_hd__a221o_1 _12709_ (.A1(_05178_),
    .A2(net196),
    .B1(_02435_),
    .B2(_05167_),
    .C1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__a221o_1 _12710_ (.A1(_02424_),
    .A2(_02756_),
    .B1(_02771_),
    .B2(net171),
    .C1(_05714_),
    .X(_05715_));
 sky130_fd_sc_hd__a21oi_1 _12711_ (.A1(_00786_),
    .A2(net257),
    .B1(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21a_1 _12712_ (.A1(_05711_),
    .A2(_05712_),
    .B1(_05716_),
    .X(_05717_));
 sky130_fd_sc_hd__o21ai_1 _12713_ (.A1(_05707_),
    .A2(_05708_),
    .B1(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__or4b_1 _12714_ (.A(_05697_),
    .B(_05701_),
    .C(_05718_),
    .D_N(_05705_),
    .X(_05719_));
 sky130_fd_sc_hd__o221a_4 _12715_ (.A1(_05123_),
    .A2(net204),
    .B1(_05693_),
    .B2(_05719_),
    .C1(net240),
    .X(dest_val[29]));
 sky130_fd_sc_hd__o21ai_2 _12716_ (.A1(_00787_),
    .A2(_05668_),
    .B1(_05670_),
    .Y(_05721_));
 sky130_fd_sc_hd__nor2_1 _12717_ (.A(_02079_),
    .B(net5),
    .Y(_05722_));
 sky130_fd_sc_hd__nor2_1 _12718_ (.A(net5),
    .B(_02187_),
    .Y(_05723_));
 sky130_fd_sc_hd__o2bb2a_1 _12719_ (.A1_N(net10),
    .A2_N(_05723_),
    .B1(_05722_),
    .B2(net61),
    .X(_05724_));
 sky130_fd_sc_hd__o31a_1 _12720_ (.A1(net10),
    .A2(net58),
    .A3(_05723_),
    .B1(_05724_),
    .X(_05725_));
 sky130_fd_sc_hd__inv_2 _12721_ (.A(_05725_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_1 _12722_ (.A(_05721_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__xnor2_1 _12723_ (.A(_05721_),
    .B(_05725_),
    .Y(_05728_));
 sky130_fd_sc_hd__nor3_1 _12724_ (.A(_05672_),
    .B(_05675_),
    .C(_05728_),
    .Y(_05729_));
 sky130_fd_sc_hd__inv_2 _12725_ (.A(_05729_),
    .Y(_05730_));
 sky130_fd_sc_hd__o21a_1 _12726_ (.A1(_05672_),
    .A2(_05675_),
    .B1(_05728_),
    .X(_05732_));
 sky130_fd_sc_hd__or2_1 _12727_ (.A(_05729_),
    .B(_05732_),
    .X(_05733_));
 sky130_fd_sc_hd__or2_1 _12728_ (.A(_05624_),
    .B(_05682_),
    .X(_05734_));
 sky130_fd_sc_hd__a2bb2o_1 _12729_ (.A1_N(_05626_),
    .A2_N(_05734_),
    .B1(_05679_),
    .B2(_05621_),
    .X(_05735_));
 sky130_fd_sc_hd__nor3_1 _12730_ (.A(_05498_),
    .B(_05625_),
    .C(_05734_),
    .Y(_05736_));
 sky130_fd_sc_hd__or3_1 _12731_ (.A(_05680_),
    .B(_05735_),
    .C(_05736_),
    .X(_05737_));
 sky130_fd_sc_hd__xnor2_2 _12732_ (.A(_05733_),
    .B(_05737_),
    .Y(_05738_));
 sky130_fd_sc_hd__or4b_2 _12733_ (.A(_05349_),
    .B(_05630_),
    .C(_05690_),
    .D_N(_05633_),
    .X(_05739_));
 sky130_fd_sc_hd__a21oi_1 _12734_ (.A1(net143),
    .A2(_05739_),
    .B1(_05738_),
    .Y(_05740_));
 sky130_fd_sc_hd__a31o_1 _12735_ (.A1(net143),
    .A2(_05738_),
    .A3(_05739_),
    .B1(_02349_),
    .X(_05741_));
 sky130_fd_sc_hd__nor2_1 _12736_ (.A(_05740_),
    .B(_05741_),
    .Y(_05743_));
 sky130_fd_sc_hd__a21o_1 _12737_ (.A1(_05156_),
    .A2(_05694_),
    .B1(_05167_),
    .X(_05744_));
 sky130_fd_sc_hd__mux2_1 _12738_ (.A0(_06632_),
    .A1(_05744_),
    .S(net284),
    .X(_05745_));
 sky130_fd_sc_hd__nand2_1 _12739_ (.A(_05091_),
    .B(_05745_),
    .Y(_05746_));
 sky130_fd_sc_hd__nand2_1 _12740_ (.A(_05091_),
    .B(_05744_),
    .Y(_05747_));
 sky130_fd_sc_hd__o211a_1 _12741_ (.A1(_05091_),
    .A2(_05745_),
    .B1(_05746_),
    .C1(_02426_),
    .X(_05748_));
 sky130_fd_sc_hd__nor2_1 _12742_ (.A(net135),
    .B(_02018_),
    .Y(_05749_));
 sky130_fd_sc_hd__xnor2_1 _12743_ (.A(_02128_),
    .B(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__xor2_1 _12744_ (.A(net288),
    .B(_05702_),
    .X(_05751_));
 sky130_fd_sc_hd__mux2_1 _12745_ (.A0(_02635_),
    .A1(_05751_),
    .S(net245),
    .X(_05752_));
 sky130_fd_sc_hd__or2_1 _12746_ (.A(\div_shifter[61] ),
    .B(_05706_),
    .X(_05754_));
 sky130_fd_sc_hd__a21oi_1 _12747_ (.A1(net229),
    .A2(_05754_),
    .B1(\div_shifter[62] ),
    .Y(_05755_));
 sky130_fd_sc_hd__a31o_1 _12748_ (.A1(\div_shifter[62] ),
    .A2(net229),
    .A3(_05754_),
    .B1(net191),
    .X(_05756_));
 sky130_fd_sc_hd__nor2_1 _12749_ (.A(_05755_),
    .B(_05756_),
    .Y(_05757_));
 sky130_fd_sc_hd__or2_1 _12750_ (.A(\div_res[29] ),
    .B(_05709_),
    .X(_05758_));
 sky130_fd_sc_hd__a21oi_1 _12751_ (.A1(net142),
    .A2(_05758_),
    .B1(\div_res[30] ),
    .Y(_05759_));
 sky130_fd_sc_hd__a31o_1 _12752_ (.A1(\div_res[30] ),
    .A2(net142),
    .A3(_05758_),
    .B1(net190),
    .X(_05760_));
 sky130_fd_sc_hd__nor2_1 _12753_ (.A(_05759_),
    .B(_05760_),
    .Y(_05761_));
 sky130_fd_sc_hd__and3_1 _12754_ (.A(_02075_),
    .B(_02076_),
    .C(net257),
    .X(_05762_));
 sky130_fd_sc_hd__o21a_1 _12755_ (.A1(net288),
    .A2(_05069_),
    .B1(_02439_),
    .X(_05763_));
 sky130_fd_sc_hd__o21ai_1 _12756_ (.A1(net288),
    .A2(net232),
    .B1(net204),
    .Y(_05765_));
 sky130_fd_sc_hd__a311o_1 _12757_ (.A1(net288),
    .A2(_05069_),
    .A3(_02435_),
    .B1(_05763_),
    .C1(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__a221o_1 _12758_ (.A1(_05091_),
    .A2(net195),
    .B1(_02635_),
    .B2(_02424_),
    .C1(_05766_),
    .X(_05767_));
 sky130_fd_sc_hd__a2111o_1 _12759_ (.A1(net172),
    .A2(_02611_),
    .B1(_05757_),
    .C1(_05762_),
    .D1(_05767_),
    .X(_05768_));
 sky130_fd_sc_hd__a211o_1 _12760_ (.A1(net205),
    .A2(_05752_),
    .B1(_05761_),
    .C1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__a211o_1 _12761_ (.A1(_02433_),
    .A2(_05750_),
    .B1(_05769_),
    .C1(_05748_),
    .X(_05770_));
 sky130_fd_sc_hd__o221a_4 _12762_ (.A1(_05069_),
    .A2(net204),
    .B1(_05743_),
    .B2(_05770_),
    .C1(net240),
    .X(dest_val[30]));
 sky130_fd_sc_hd__o21ai_1 _12763_ (.A1(_05738_),
    .A2(_05739_),
    .B1(net142),
    .Y(_05771_));
 sky130_fd_sc_hd__nand2_1 _12764_ (.A(net5),
    .B(net61),
    .Y(_05772_));
 sky130_fd_sc_hd__nor2_1 _12765_ (.A(_05682_),
    .B(_05733_),
    .Y(_05773_));
 sky130_fd_sc_hd__a221o_1 _12766_ (.A1(_05680_),
    .A2(_05730_),
    .B1(_05773_),
    .B2(_05685_),
    .C1(_05732_),
    .X(_05775_));
 sky130_fd_sc_hd__a31o_1 _12767_ (.A1(_05566_),
    .A2(_05683_),
    .A3(_05773_),
    .B1(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__xnor2_1 _12768_ (.A(_05772_),
    .B(_05776_),
    .Y(_05777_));
 sky130_fd_sc_hd__mux2_1 _12769_ (.A0(_05721_),
    .A1(_05727_),
    .S(_05724_),
    .X(_05778_));
 sky130_fd_sc_hd__and2_1 _12770_ (.A(_05777_),
    .B(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__nand2_1 _12771_ (.A(_05777_),
    .B(_05778_),
    .Y(_05780_));
 sky130_fd_sc_hd__nor2_1 _12772_ (.A(_05777_),
    .B(_05778_),
    .Y(_05781_));
 sky130_fd_sc_hd__or2_1 _12773_ (.A(_05777_),
    .B(_05778_),
    .X(_05782_));
 sky130_fd_sc_hd__o221a_1 _12774_ (.A1(_05738_),
    .A2(_05739_),
    .B1(_05779_),
    .B2(_05781_),
    .C1(net142),
    .X(_05783_));
 sky130_fd_sc_hd__a311oi_4 _12775_ (.A1(_05771_),
    .A2(_05780_),
    .A3(_05782_),
    .B1(_05783_),
    .C1(_02349_),
    .Y(_05784_));
 sky130_fd_sc_hd__a21oi_1 _12776_ (.A1(net288),
    .A2(_05069_),
    .B1(net295),
    .Y(_05786_));
 sky130_fd_sc_hd__a22o_1 _12777_ (.A1(net295),
    .A2(_06633_),
    .B1(_05747_),
    .B2(_05786_),
    .X(_05787_));
 sky130_fd_sc_hd__xor2_1 _12778_ (.A(_04949_),
    .B(_05787_),
    .X(_05788_));
 sky130_fd_sc_hd__a21o_1 _12779_ (.A1(_02018_),
    .A2(_02128_),
    .B1(net135),
    .X(_05789_));
 sky130_fd_sc_hd__xnor2_1 _12780_ (.A(_02240_),
    .B(_05789_),
    .Y(_05790_));
 sky130_fd_sc_hd__nand2_1 _12781_ (.A(_02433_),
    .B(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__and3_1 _12782_ (.A(net288),
    .B(net245),
    .C(_05702_),
    .X(_05792_));
 sky130_fd_sc_hd__xor2_1 _12783_ (.A(_02457_),
    .B(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__o21a_1 _12784_ (.A1(\div_res[30] ),
    .A2(_05758_),
    .B1(net142),
    .X(_05794_));
 sky130_fd_sc_hd__xnor2_1 _12785_ (.A(\div_res[31] ),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__o21a_1 _12786_ (.A1(\div_shifter[62] ),
    .A2(_05754_),
    .B1(net229),
    .X(_05797_));
 sky130_fd_sc_hd__xnor2_1 _12787_ (.A(\div_shifter[63] ),
    .B(_05797_),
    .Y(_05798_));
 sky130_fd_sc_hd__a21oi_1 _12788_ (.A1(reg1_val[31]),
    .A2(_02075_),
    .B1(_02432_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21ai_1 _12789_ (.A1(reg1_val[31]),
    .A2(_02075_),
    .B1(_05799_),
    .Y(_05800_));
 sky130_fd_sc_hd__o21ai_1 _12790_ (.A1(reg1_val[31]),
    .A2(net232),
    .B1(net204),
    .Y(_05801_));
 sky130_fd_sc_hd__o21a_1 _12791_ (.A1(reg1_val[31]),
    .A2(_04917_),
    .B1(_02439_),
    .X(_05802_));
 sky130_fd_sc_hd__a311o_1 _12792_ (.A1(reg1_val[31]),
    .A2(_04917_),
    .A3(_02435_),
    .B1(_05801_),
    .C1(_05802_),
    .X(_05803_));
 sky130_fd_sc_hd__a21oi_1 _12793_ (.A1(_04949_),
    .A2(net195),
    .B1(_05803_),
    .Y(_05804_));
 sky130_fd_sc_hd__o221a_1 _12794_ (.A1(net169),
    .A2(_02419_),
    .B1(_02425_),
    .B2(_02457_),
    .C1(_05804_),
    .X(_05805_));
 sky130_fd_sc_hd__o211a_1 _12795_ (.A1(net190),
    .A2(_05795_),
    .B1(_05800_),
    .C1(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__o21a_1 _12796_ (.A1(net192),
    .A2(_05798_),
    .B1(_05806_),
    .X(_05808_));
 sky130_fd_sc_hd__o211a_1 _12797_ (.A1(_06667_),
    .A2(_05793_),
    .B1(_05808_),
    .C1(_05791_),
    .X(_05809_));
 sky130_fd_sc_hd__o21ai_1 _12798_ (.A1(_02427_),
    .A2(_05788_),
    .B1(_05809_),
    .Y(_05810_));
 sky130_fd_sc_hd__o221a_4 _12799_ (.A1(_04917_),
    .A2(net204),
    .B1(_05784_),
    .B2(_05810_),
    .C1(net240),
    .X(dest_val[31]));
 sky130_fd_sc_hd__mux2_1 _12800_ (.A0(net291),
    .A1(curr_PC[0]),
    .S(net238),
    .X(_05811_));
 sky130_fd_sc_hd__nand2_1 _12801_ (.A(_04829_),
    .B(_05811_),
    .Y(_05812_));
 sky130_fd_sc_hd__or2_1 _12802_ (.A(_04829_),
    .B(_05811_),
    .X(_05813_));
 sky130_fd_sc_hd__and2_4 _12803_ (.A(_05812_),
    .B(_05813_),
    .X(new_PC[0]));
 sky130_fd_sc_hd__mux2_1 _12804_ (.A0(net289),
    .A1(curr_PC[1]),
    .S(net237),
    .X(_05814_));
 sky130_fd_sc_hd__nand2_1 _12805_ (.A(_06085_),
    .B(_05814_),
    .Y(_05815_));
 sky130_fd_sc_hd__or2_1 _12806_ (.A(_06085_),
    .B(_05814_),
    .X(_05817_));
 sky130_fd_sc_hd__nand2_1 _12807_ (.A(_05815_),
    .B(_05817_),
    .Y(_05818_));
 sky130_fd_sc_hd__or2_1 _12808_ (.A(_05812_),
    .B(_05818_),
    .X(_05819_));
 sky130_fd_sc_hd__nand2_1 _12809_ (.A(_05812_),
    .B(_05818_),
    .Y(_05820_));
 sky130_fd_sc_hd__and2_4 _12810_ (.A(_05819_),
    .B(_05820_),
    .X(new_PC[1]));
 sky130_fd_sc_hd__mux2_1 _12811_ (.A0(reg1_val[2]),
    .A1(curr_PC[2]),
    .S(net237),
    .X(_05821_));
 sky130_fd_sc_hd__nand2_1 _12812_ (.A(_06004_),
    .B(_05821_),
    .Y(_05822_));
 sky130_fd_sc_hd__or2_1 _12813_ (.A(_06004_),
    .B(_05821_),
    .X(_05823_));
 sky130_fd_sc_hd__nand2_1 _12814_ (.A(_05822_),
    .B(_05823_),
    .Y(_05824_));
 sky130_fd_sc_hd__a21o_1 _12815_ (.A1(_05815_),
    .A2(_05819_),
    .B1(_05824_),
    .X(_05825_));
 sky130_fd_sc_hd__nand3_1 _12816_ (.A(_05815_),
    .B(_05819_),
    .C(_05824_),
    .Y(_05827_));
 sky130_fd_sc_hd__and2_4 _12817_ (.A(_05825_),
    .B(_05827_),
    .X(new_PC[2]));
 sky130_fd_sc_hd__mux2_1 _12818_ (.A0(reg1_val[3]),
    .A1(curr_PC[3]),
    .S(net237),
    .X(_05828_));
 sky130_fd_sc_hd__nand2_1 _12819_ (.A(_05921_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__or2_1 _12820_ (.A(_05921_),
    .B(_05828_),
    .X(_05830_));
 sky130_fd_sc_hd__nand2_1 _12821_ (.A(_05829_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__a21o_1 _12822_ (.A1(_05822_),
    .A2(_05825_),
    .B1(_05831_),
    .X(_05832_));
 sky130_fd_sc_hd__nand3_1 _12823_ (.A(_05822_),
    .B(_05825_),
    .C(_05831_),
    .Y(_05833_));
 sky130_fd_sc_hd__and2_4 _12824_ (.A(_05832_),
    .B(_05833_),
    .X(new_PC[3]));
 sky130_fd_sc_hd__mux2_1 _12825_ (.A0(reg1_val[4]),
    .A1(curr_PC[4]),
    .S(net237),
    .X(_05834_));
 sky130_fd_sc_hd__nand2_1 _12826_ (.A(_05854_),
    .B(_05834_),
    .Y(_05836_));
 sky130_fd_sc_hd__or2_1 _12827_ (.A(_05854_),
    .B(_05834_),
    .X(_05837_));
 sky130_fd_sc_hd__nand2_1 _12828_ (.A(_05836_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__a21o_1 _12829_ (.A1(_05829_),
    .A2(_05832_),
    .B1(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__nand3_1 _12830_ (.A(_05829_),
    .B(_05832_),
    .C(_05838_),
    .Y(_05840_));
 sky130_fd_sc_hd__and2_4 _12831_ (.A(_05839_),
    .B(_05840_),
    .X(new_PC[4]));
 sky130_fd_sc_hd__mux2_1 _12832_ (.A0(reg1_val[5]),
    .A1(curr_PC[5]),
    .S(net238),
    .X(_05841_));
 sky130_fd_sc_hd__nand2_1 _12833_ (.A(_05710_),
    .B(_05841_),
    .Y(_05842_));
 sky130_fd_sc_hd__or2_1 _12834_ (.A(_05710_),
    .B(_05841_),
    .X(_05843_));
 sky130_fd_sc_hd__nand2_1 _12835_ (.A(_05842_),
    .B(_05843_),
    .Y(_05844_));
 sky130_fd_sc_hd__a21o_1 _12836_ (.A1(_05836_),
    .A2(_05839_),
    .B1(_05844_),
    .X(_05846_));
 sky130_fd_sc_hd__nand3_1 _12837_ (.A(_05836_),
    .B(_05839_),
    .C(_05844_),
    .Y(_05847_));
 sky130_fd_sc_hd__and2_4 _12838_ (.A(_05846_),
    .B(_05847_),
    .X(new_PC[5]));
 sky130_fd_sc_hd__mux2_1 _12839_ (.A0(reg1_val[6]),
    .A1(curr_PC[6]),
    .S(net238),
    .X(_05848_));
 sky130_fd_sc_hd__nand2_1 _12840_ (.A(_05774_),
    .B(_05848_),
    .Y(_05849_));
 sky130_fd_sc_hd__or2_1 _12841_ (.A(_05774_),
    .B(_05848_),
    .X(_05850_));
 sky130_fd_sc_hd__nand2_1 _12842_ (.A(_05849_),
    .B(_05850_),
    .Y(_05851_));
 sky130_fd_sc_hd__a21o_1 _12843_ (.A1(_05842_),
    .A2(_05846_),
    .B1(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__nand3_1 _12844_ (.A(_05842_),
    .B(_05846_),
    .C(_05851_),
    .Y(_05853_));
 sky130_fd_sc_hd__and2_4 _12845_ (.A(_05852_),
    .B(_05853_),
    .X(new_PC[6]));
 sky130_fd_sc_hd__mux2_1 _12846_ (.A0(net287),
    .A1(curr_PC[7]),
    .S(net238),
    .X(_05855_));
 sky130_fd_sc_hd__nand2_1 _12847_ (.A(_05634_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__or2_1 _12848_ (.A(_05634_),
    .B(_05855_),
    .X(_05857_));
 sky130_fd_sc_hd__nand2_1 _12849_ (.A(_05856_),
    .B(_05857_),
    .Y(_05858_));
 sky130_fd_sc_hd__a21o_1 _12850_ (.A1(_05849_),
    .A2(_05852_),
    .B1(_05858_),
    .X(_05859_));
 sky130_fd_sc_hd__nand3_1 _12851_ (.A(_05849_),
    .B(_05852_),
    .C(_05858_),
    .Y(_05860_));
 sky130_fd_sc_hd__and2_4 _12852_ (.A(_05859_),
    .B(_05860_),
    .X(new_PC[7]));
 sky130_fd_sc_hd__mux2_1 _12853_ (.A0(reg1_val[8]),
    .A1(curr_PC[8]),
    .S(net238),
    .X(_05861_));
 sky130_fd_sc_hd__nand2_1 _12854_ (.A(_05569_),
    .B(_05861_),
    .Y(_05862_));
 sky130_fd_sc_hd__or2_1 _12855_ (.A(_05569_),
    .B(_05861_),
    .X(_05863_));
 sky130_fd_sc_hd__nand2_1 _12856_ (.A(_05862_),
    .B(_05863_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21o_1 _12857_ (.A1(_05856_),
    .A2(_05859_),
    .B1(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__nand3_1 _12858_ (.A(_05856_),
    .B(_05859_),
    .C(_05865_),
    .Y(_05867_));
 sky130_fd_sc_hd__and2_4 _12859_ (.A(_05866_),
    .B(_05867_),
    .X(new_PC[8]));
 sky130_fd_sc_hd__mux2_1 _12860_ (.A0(reg1_val[9]),
    .A1(curr_PC[9]),
    .S(net238),
    .X(_05868_));
 sky130_fd_sc_hd__nand2_1 _12861_ (.A(_05461_),
    .B(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__or2_1 _12862_ (.A(_05461_),
    .B(_05868_),
    .X(_05870_));
 sky130_fd_sc_hd__nand2_1 _12863_ (.A(_05869_),
    .B(_05870_),
    .Y(_05871_));
 sky130_fd_sc_hd__a21o_1 _12864_ (.A1(_05862_),
    .A2(_05866_),
    .B1(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__nand3_1 _12865_ (.A(_05862_),
    .B(_05866_),
    .C(_05871_),
    .Y(_05873_));
 sky130_fd_sc_hd__and2_4 _12866_ (.A(_05872_),
    .B(_05873_),
    .X(new_PC[9]));
 sky130_fd_sc_hd__mux2_1 _12867_ (.A0(reg1_val[10]),
    .A1(curr_PC[10]),
    .S(net238),
    .X(_05875_));
 sky130_fd_sc_hd__nand2_1 _12868_ (.A(_05287_),
    .B(_05875_),
    .Y(_05876_));
 sky130_fd_sc_hd__or2_1 _12869_ (.A(_05287_),
    .B(_05875_),
    .X(_05877_));
 sky130_fd_sc_hd__nand2_1 _12870_ (.A(_05876_),
    .B(_05877_),
    .Y(_05878_));
 sky130_fd_sc_hd__a21o_1 _12871_ (.A1(_05869_),
    .A2(_05872_),
    .B1(_05878_),
    .X(_05879_));
 sky130_fd_sc_hd__nand3_1 _12872_ (.A(_05869_),
    .B(_05872_),
    .C(_05878_),
    .Y(_05880_));
 sky130_fd_sc_hd__and2_4 _12873_ (.A(_05879_),
    .B(_05880_),
    .X(new_PC[10]));
 sky130_fd_sc_hd__mux2_1 _12874_ (.A0(net290),
    .A1(curr_PC[11]),
    .S(net239),
    .X(_05881_));
 sky130_fd_sc_hd__nand2_1 _12875_ (.A(_05363_),
    .B(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__or2_1 _12876_ (.A(_05363_),
    .B(_05881_),
    .X(_05884_));
 sky130_fd_sc_hd__nand2_1 _12877_ (.A(_05882_),
    .B(_05884_),
    .Y(_05885_));
 sky130_fd_sc_hd__a21o_1 _12878_ (.A1(_05876_),
    .A2(_05879_),
    .B1(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__nand3_1 _12879_ (.A(_05876_),
    .B(_05879_),
    .C(_05885_),
    .Y(_05887_));
 sky130_fd_sc_hd__and2_4 _12880_ (.A(_05886_),
    .B(_05887_),
    .X(new_PC[11]));
 sky130_fd_sc_hd__mux2_1 _12881_ (.A0(reg1_val[12]),
    .A1(curr_PC[12]),
    .S(net239),
    .X(_05888_));
 sky130_fd_sc_hd__nand2_1 _12882_ (.A(_04960_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__or2_1 _12883_ (.A(_04960_),
    .B(_05888_),
    .X(_05890_));
 sky130_fd_sc_hd__nand2_1 _12884_ (.A(_05889_),
    .B(_05890_),
    .Y(_05891_));
 sky130_fd_sc_hd__a21o_1 _12885_ (.A1(_05882_),
    .A2(_05886_),
    .B1(_05891_),
    .X(_05892_));
 sky130_fd_sc_hd__nand3_1 _12886_ (.A(_05882_),
    .B(_05886_),
    .C(_05891_),
    .Y(_05894_));
 sky130_fd_sc_hd__and2_4 _12887_ (.A(_05892_),
    .B(_05894_),
    .X(new_PC[12]));
 sky130_fd_sc_hd__mux2_1 _12888_ (.A0(reg1_val[13]),
    .A1(curr_PC[13]),
    .S(net239),
    .X(_05895_));
 sky130_fd_sc_hd__nand2_1 _12889_ (.A(_05189_),
    .B(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__or2_1 _12890_ (.A(_05189_),
    .B(_05895_),
    .X(_05897_));
 sky130_fd_sc_hd__nand2_1 _12891_ (.A(_05896_),
    .B(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__a21o_1 _12892_ (.A1(_05889_),
    .A2(_05892_),
    .B1(_05898_),
    .X(_05899_));
 sky130_fd_sc_hd__nand3_1 _12893_ (.A(_05889_),
    .B(_05892_),
    .C(_05898_),
    .Y(_05900_));
 sky130_fd_sc_hd__and2_4 _12894_ (.A(_05899_),
    .B(_05900_),
    .X(new_PC[13]));
 sky130_fd_sc_hd__mux2_1 _12895_ (.A0(reg1_val[14]),
    .A1(curr_PC[14]),
    .S(net239),
    .X(_05901_));
 sky130_fd_sc_hd__nand2_1 _12896_ (.A(_05102_),
    .B(_05901_),
    .Y(_05903_));
 sky130_fd_sc_hd__or2_1 _12897_ (.A(_05102_),
    .B(_05901_),
    .X(_05904_));
 sky130_fd_sc_hd__nand2_1 _12898_ (.A(_05903_),
    .B(_05904_),
    .Y(_05905_));
 sky130_fd_sc_hd__a21o_1 _12899_ (.A1(_05896_),
    .A2(_05899_),
    .B1(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__nand3_1 _12900_ (.A(_05896_),
    .B(_05899_),
    .C(_05905_),
    .Y(_05907_));
 sky130_fd_sc_hd__and2_4 _12901_ (.A(_05906_),
    .B(_05907_),
    .X(new_PC[14]));
 sky130_fd_sc_hd__mux2_1 _12902_ (.A0(reg1_val[15]),
    .A1(curr_PC[15]),
    .S(net239),
    .X(_05908_));
 sky130_fd_sc_hd__nand2_1 _12903_ (.A(_05047_),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__or2_1 _12904_ (.A(_05047_),
    .B(_05908_),
    .X(_05910_));
 sky130_fd_sc_hd__nand2_1 _12905_ (.A(_05909_),
    .B(_05910_),
    .Y(_05911_));
 sky130_fd_sc_hd__a21o_1 _12906_ (.A1(_05903_),
    .A2(_05906_),
    .B1(_05911_),
    .X(_05913_));
 sky130_fd_sc_hd__nand3_1 _12907_ (.A(_05903_),
    .B(_05906_),
    .C(_05911_),
    .Y(_05914_));
 sky130_fd_sc_hd__and2_4 _12908_ (.A(_05913_),
    .B(_05914_),
    .X(new_PC[15]));
 sky130_fd_sc_hd__mux2_2 _12909_ (.A0(reg1_val[16]),
    .A1(curr_PC[16]),
    .S(net239),
    .X(_05915_));
 sky130_fd_sc_hd__xnor2_1 _12910_ (.A(net262),
    .B(_05915_),
    .Y(_05916_));
 sky130_fd_sc_hd__a21o_1 _12911_ (.A1(_05909_),
    .A2(_05913_),
    .B1(_05916_),
    .X(_05917_));
 sky130_fd_sc_hd__nand3_1 _12912_ (.A(_05909_),
    .B(_05913_),
    .C(_05916_),
    .Y(_05918_));
 sky130_fd_sc_hd__and2_4 _12913_ (.A(_05917_),
    .B(_05918_),
    .X(new_PC[16]));
 sky130_fd_sc_hd__mux2_2 _12914_ (.A0(reg1_val[17]),
    .A1(curr_PC[17]),
    .S(net239),
    .X(_05919_));
 sky130_fd_sc_hd__xnor2_4 _12915_ (.A(net262),
    .B(_05919_),
    .Y(_05920_));
 sky130_fd_sc_hd__a21bo_1 _12916_ (.A1(net262),
    .A2(_05915_),
    .B1_N(_05917_),
    .X(_05922_));
 sky130_fd_sc_hd__xnor2_4 _12917_ (.A(_05920_),
    .B(_05922_),
    .Y(new_PC[17]));
 sky130_fd_sc_hd__mux2_1 _12918_ (.A0(reg1_val[18]),
    .A1(curr_PC[18]),
    .S(net239),
    .X(_05923_));
 sky130_fd_sc_hd__nand2_1 _12919_ (.A(net262),
    .B(_05923_),
    .Y(_05924_));
 sky130_fd_sc_hd__or2_1 _12920_ (.A(net262),
    .B(_05923_),
    .X(_05925_));
 sky130_fd_sc_hd__nand2_1 _12921_ (.A(_05924_),
    .B(_05925_),
    .Y(_05926_));
 sky130_fd_sc_hd__or2_1 _12922_ (.A(_05917_),
    .B(_05920_),
    .X(_05927_));
 sky130_fd_sc_hd__o21ai_1 _12923_ (.A1(_05915_),
    .A2(_05919_),
    .B1(net262),
    .Y(_05928_));
 sky130_fd_sc_hd__a21o_1 _12924_ (.A1(_05927_),
    .A2(_05928_),
    .B1(_05926_),
    .X(_05929_));
 sky130_fd_sc_hd__nand3_1 _12925_ (.A(_05926_),
    .B(_05927_),
    .C(_05928_),
    .Y(_05930_));
 sky130_fd_sc_hd__and2_4 _12926_ (.A(_05929_),
    .B(_05930_),
    .X(new_PC[18]));
 sky130_fd_sc_hd__mux2_1 _12927_ (.A0(reg1_val[19]),
    .A1(curr_PC[19]),
    .S(net239),
    .X(_05932_));
 sky130_fd_sc_hd__nand2_1 _12928_ (.A(net262),
    .B(_05932_),
    .Y(_05933_));
 sky130_fd_sc_hd__or2_1 _12929_ (.A(net262),
    .B(_05932_),
    .X(_05934_));
 sky130_fd_sc_hd__nand2_2 _12930_ (.A(_05933_),
    .B(_05934_),
    .Y(_05935_));
 sky130_fd_sc_hd__nand2_2 _12931_ (.A(_05924_),
    .B(_05929_),
    .Y(_05936_));
 sky130_fd_sc_hd__xnor2_4 _12932_ (.A(_05935_),
    .B(_05936_),
    .Y(new_PC[19]));
 sky130_fd_sc_hd__mux2_1 _12933_ (.A0(reg1_val[20]),
    .A1(curr_PC[20]),
    .S(net239),
    .X(_05937_));
 sky130_fd_sc_hd__nand2_1 _12934_ (.A(net262),
    .B(_05937_),
    .Y(_05938_));
 sky130_fd_sc_hd__or2_1 _12935_ (.A(net262),
    .B(_05937_),
    .X(_05939_));
 sky130_fd_sc_hd__nand2_2 _12936_ (.A(_05938_),
    .B(_05939_),
    .Y(_05941_));
 sky130_fd_sc_hd__or3_1 _12937_ (.A(_05926_),
    .B(_05927_),
    .C(_05935_),
    .X(_05942_));
 sky130_fd_sc_hd__and3_1 _12938_ (.A(_05924_),
    .B(_05928_),
    .C(_05933_),
    .X(_05943_));
 sky130_fd_sc_hd__nand2_2 _12939_ (.A(_05942_),
    .B(_05943_),
    .Y(_05944_));
 sky130_fd_sc_hd__inv_2 _12940_ (.A(_05944_),
    .Y(_05945_));
 sky130_fd_sc_hd__xnor2_4 _12941_ (.A(_05941_),
    .B(_05944_),
    .Y(new_PC[20]));
 sky130_fd_sc_hd__mux2_2 _12942_ (.A0(reg1_val[21]),
    .A1(curr_PC[21]),
    .S(net239),
    .X(_05946_));
 sky130_fd_sc_hd__xnor2_4 _12943_ (.A(net262),
    .B(_05946_),
    .Y(_05947_));
 sky130_fd_sc_hd__o21ai_2 _12944_ (.A1(_05941_),
    .A2(_05945_),
    .B1(_05938_),
    .Y(_05948_));
 sky130_fd_sc_hd__xnor2_4 _12945_ (.A(_05947_),
    .B(_05948_),
    .Y(new_PC[21]));
 sky130_fd_sc_hd__mux2_1 _12946_ (.A0(reg1_val[22]),
    .A1(curr_PC[22]),
    .S(net239),
    .X(_05950_));
 sky130_fd_sc_hd__and2_1 _12947_ (.A(net262),
    .B(_05950_),
    .X(_05951_));
 sky130_fd_sc_hd__or2_1 _12948_ (.A(net262),
    .B(_05950_),
    .X(_05952_));
 sky130_fd_sc_hd__nand2b_2 _12949_ (.A_N(_05951_),
    .B(_05952_),
    .Y(_05953_));
 sky130_fd_sc_hd__o21ai_2 _12950_ (.A1(_05937_),
    .A2(_05946_),
    .B1(net262),
    .Y(_05954_));
 sky130_fd_sc_hd__nor2_1 _12951_ (.A(_05941_),
    .B(_05947_),
    .Y(_05955_));
 sky130_fd_sc_hd__inv_2 _12952_ (.A(_05955_),
    .Y(_05956_));
 sky130_fd_sc_hd__o21ai_4 _12953_ (.A1(_05945_),
    .A2(_05956_),
    .B1(_05954_),
    .Y(_05957_));
 sky130_fd_sc_hd__xnor2_4 _12954_ (.A(_05953_),
    .B(_05957_),
    .Y(new_PC[22]));
 sky130_fd_sc_hd__mux2_2 _12955_ (.A0(reg1_val[23]),
    .A1(curr_PC[23]),
    .S(net239),
    .X(_05958_));
 sky130_fd_sc_hd__xnor2_4 _12956_ (.A(net262),
    .B(_05958_),
    .Y(_05960_));
 sky130_fd_sc_hd__a21o_1 _12957_ (.A1(_05952_),
    .A2(_05957_),
    .B1(_05951_),
    .X(_05961_));
 sky130_fd_sc_hd__xnor2_4 _12958_ (.A(_05960_),
    .B(_05961_),
    .Y(new_PC[23]));
 sky130_fd_sc_hd__mux2_2 _12959_ (.A0(reg1_val[24]),
    .A1(curr_PC[24]),
    .S(net239),
    .X(_05962_));
 sky130_fd_sc_hd__xnor2_4 _12960_ (.A(net263),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__or4_1 _12961_ (.A(_05942_),
    .B(_05953_),
    .C(_05956_),
    .D(_05960_),
    .X(_05964_));
 sky130_fd_sc_hd__o21ai_1 _12962_ (.A1(_05950_),
    .A2(_05958_),
    .B1(net262),
    .Y(_05965_));
 sky130_fd_sc_hd__and4_2 _12963_ (.A(_05943_),
    .B(_05954_),
    .C(_05964_),
    .D(_05965_),
    .X(_05966_));
 sky130_fd_sc_hd__xor2_4 _12964_ (.A(_05963_),
    .B(_05966_),
    .X(new_PC[24]));
 sky130_fd_sc_hd__mux2_1 _12965_ (.A0(reg1_val[25]),
    .A1(curr_PC[25]),
    .S(net239),
    .X(_05967_));
 sky130_fd_sc_hd__and2_1 _12966_ (.A(net263),
    .B(_05967_),
    .X(_05969_));
 sky130_fd_sc_hd__nor2_1 _12967_ (.A(net263),
    .B(_05967_),
    .Y(_05970_));
 sky130_fd_sc_hd__nor2_2 _12968_ (.A(_05969_),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__o2bb2a_2 _12969_ (.A1_N(net263),
    .A2_N(_05962_),
    .B1(_05963_),
    .B2(_05966_),
    .X(_05972_));
 sky130_fd_sc_hd__xnor2_4 _12970_ (.A(_05971_),
    .B(_05972_),
    .Y(new_PC[25]));
 sky130_fd_sc_hd__mux2_1 _12971_ (.A0(reg1_val[26]),
    .A1(curr_PC[26]),
    .S(net240),
    .X(_05973_));
 sky130_fd_sc_hd__and2_1 _12972_ (.A(net263),
    .B(_05973_),
    .X(_05974_));
 sky130_fd_sc_hd__nor2_1 _12973_ (.A(net263),
    .B(_05973_),
    .Y(_05975_));
 sky130_fd_sc_hd__nor2_2 _12974_ (.A(_05974_),
    .B(_05975_),
    .Y(_05976_));
 sky130_fd_sc_hd__o21ba_2 _12975_ (.A1(_05970_),
    .A2(_05972_),
    .B1_N(_05969_),
    .X(_05977_));
 sky130_fd_sc_hd__xnor2_4 _12976_ (.A(_05976_),
    .B(_05977_),
    .Y(new_PC[26]));
 sky130_fd_sc_hd__o21ba_2 _12977_ (.A1(_05975_),
    .A2(_05977_),
    .B1_N(_05974_),
    .X(_05979_));
 sky130_fd_sc_hd__mux2_2 _12978_ (.A0(reg1_val[27]),
    .A1(curr_PC[27]),
    .S(net239),
    .X(_05980_));
 sky130_fd_sc_hd__xor2_2 _12979_ (.A(net263),
    .B(_05980_),
    .X(_05981_));
 sky130_fd_sc_hd__xnor2_4 _12980_ (.A(_05979_),
    .B(_05981_),
    .Y(new_PC[27]));
 sky130_fd_sc_hd__and3_4 _12981_ (.A(instruction[25]),
    .B(net292),
    .C(net266),
    .X(_05982_));
 sky130_fd_sc_hd__nor2_2 _12982_ (.A(net292),
    .B(_04829_),
    .Y(_05983_));
 sky130_fd_sc_hd__nor2_8 _12983_ (.A(_05982_),
    .B(_05983_),
    .Y(loadstore_address[0]));
 sky130_fd_sc_hd__nor2_1 _12984_ (.A(_04467_),
    .B(_06094_),
    .Y(_05984_));
 sky130_fd_sc_hd__nand2_2 _12985_ (.A(_04467_),
    .B(_06094_),
    .Y(_05985_));
 sky130_fd_sc_hd__nand2b_2 _12986_ (.A_N(_05984_),
    .B(_05985_),
    .Y(_05987_));
 sky130_fd_sc_hd__xnor2_4 _12987_ (.A(_05982_),
    .B(_05987_),
    .Y(loadstore_address[1]));
 sky130_fd_sc_hd__a21oi_4 _12988_ (.A1(_05982_),
    .A2(_05985_),
    .B1(_05984_),
    .Y(_05988_));
 sky130_fd_sc_hd__nor2_1 _12989_ (.A(reg1_val[2]),
    .B(_06004_),
    .Y(_05989_));
 sky130_fd_sc_hd__nand2_1 _12990_ (.A(reg1_val[2]),
    .B(_06004_),
    .Y(_05990_));
 sky130_fd_sc_hd__nand2b_2 _12991_ (.A_N(_05989_),
    .B(_05990_),
    .Y(_05991_));
 sky130_fd_sc_hd__xor2_4 _12992_ (.A(_05988_),
    .B(_05991_),
    .X(loadstore_address[2]));
 sky130_fd_sc_hd__o21a_2 _12993_ (.A1(_05988_),
    .A2(_05989_),
    .B1(_05990_),
    .X(_05992_));
 sky130_fd_sc_hd__nor2_1 _12994_ (.A(reg1_val[3]),
    .B(_05921_),
    .Y(_05993_));
 sky130_fd_sc_hd__nand2_1 _12995_ (.A(reg1_val[3]),
    .B(_05921_),
    .Y(_05994_));
 sky130_fd_sc_hd__and2b_1 _12996_ (.A_N(_05993_),
    .B(_05994_),
    .X(_05996_));
 sky130_fd_sc_hd__xnor2_4 _12997_ (.A(_05992_),
    .B(_05996_),
    .Y(loadstore_address[3]));
 sky130_fd_sc_hd__o21a_2 _12998_ (.A1(_05992_),
    .A2(_05993_),
    .B1(_05994_),
    .X(_05997_));
 sky130_fd_sc_hd__nor2_1 _12999_ (.A(reg1_val[4]),
    .B(_05854_),
    .Y(_05998_));
 sky130_fd_sc_hd__nand2_1 _13000_ (.A(reg1_val[4]),
    .B(_05854_),
    .Y(_05999_));
 sky130_fd_sc_hd__and2b_1 _13001_ (.A_N(_05998_),
    .B(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__xnor2_4 _13002_ (.A(_05997_),
    .B(_06000_),
    .Y(loadstore_address[4]));
 sky130_fd_sc_hd__o21a_2 _13003_ (.A1(_05997_),
    .A2(_05998_),
    .B1(_05999_),
    .X(_06001_));
 sky130_fd_sc_hd__nor2_1 _13004_ (.A(reg1_val[5]),
    .B(_05710_),
    .Y(_06002_));
 sky130_fd_sc_hd__nand2_1 _13005_ (.A(reg1_val[5]),
    .B(_05710_),
    .Y(_06003_));
 sky130_fd_sc_hd__nand2b_2 _13006_ (.A_N(_06002_),
    .B(_06003_),
    .Y(_06005_));
 sky130_fd_sc_hd__xor2_4 _13007_ (.A(_06001_),
    .B(_06005_),
    .X(loadstore_address[5]));
 sky130_fd_sc_hd__o21a_2 _13008_ (.A1(_06001_),
    .A2(_06002_),
    .B1(_06003_),
    .X(_06006_));
 sky130_fd_sc_hd__nor2_1 _13009_ (.A(reg1_val[6]),
    .B(_05774_),
    .Y(_06007_));
 sky130_fd_sc_hd__nand2_1 _13010_ (.A(reg1_val[6]),
    .B(_05774_),
    .Y(_06008_));
 sky130_fd_sc_hd__and2b_1 _13011_ (.A_N(_06007_),
    .B(_06008_),
    .X(_06009_));
 sky130_fd_sc_hd__xnor2_4 _13012_ (.A(_06006_),
    .B(_06009_),
    .Y(loadstore_address[6]));
 sky130_fd_sc_hd__o21a_2 _13013_ (.A1(_06006_),
    .A2(_06007_),
    .B1(_06008_),
    .X(_06010_));
 sky130_fd_sc_hd__nor2_1 _13014_ (.A(reg1_val[7]),
    .B(_05634_),
    .Y(_06011_));
 sky130_fd_sc_hd__nand2_1 _13015_ (.A(net287),
    .B(_05634_),
    .Y(_06012_));
 sky130_fd_sc_hd__nand2b_2 _13016_ (.A_N(_06011_),
    .B(_06012_),
    .Y(_06014_));
 sky130_fd_sc_hd__xor2_4 _13017_ (.A(_06010_),
    .B(_06014_),
    .X(loadstore_address[7]));
 sky130_fd_sc_hd__o21a_2 _13018_ (.A1(_06010_),
    .A2(_06011_),
    .B1(_06012_),
    .X(_06015_));
 sky130_fd_sc_hd__nor2_1 _13019_ (.A(reg1_val[8]),
    .B(_05569_),
    .Y(_06016_));
 sky130_fd_sc_hd__nand2_1 _13020_ (.A(reg1_val[8]),
    .B(_05569_),
    .Y(_06017_));
 sky130_fd_sc_hd__nand2b_2 _13021_ (.A_N(_06016_),
    .B(_06017_),
    .Y(_06018_));
 sky130_fd_sc_hd__xor2_4 _13022_ (.A(_06015_),
    .B(_06018_),
    .X(loadstore_address[8]));
 sky130_fd_sc_hd__o21a_2 _13023_ (.A1(_06015_),
    .A2(_06016_),
    .B1(_06017_),
    .X(_06019_));
 sky130_fd_sc_hd__or2_1 _13024_ (.A(reg1_val[9]),
    .B(_05461_),
    .X(_06020_));
 sky130_fd_sc_hd__nand2_1 _13025_ (.A(reg1_val[9]),
    .B(_05461_),
    .Y(_06021_));
 sky130_fd_sc_hd__nand2_2 _13026_ (.A(_06020_),
    .B(_06021_),
    .Y(_06023_));
 sky130_fd_sc_hd__xor2_4 _13027_ (.A(_06019_),
    .B(_06023_),
    .X(loadstore_address[9]));
 sky130_fd_sc_hd__or2_1 _13028_ (.A(reg1_val[10]),
    .B(_05287_),
    .X(_06024_));
 sky130_fd_sc_hd__nand2_1 _13029_ (.A(reg1_val[10]),
    .B(_05287_),
    .Y(_06025_));
 sky130_fd_sc_hd__nand2_1 _13030_ (.A(_06024_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__nand2b_1 _13031_ (.A_N(_06019_),
    .B(_06020_),
    .Y(_06027_));
 sky130_fd_sc_hd__a21o_1 _13032_ (.A1(_06021_),
    .A2(_06027_),
    .B1(_06026_),
    .X(_06028_));
 sky130_fd_sc_hd__nand3_1 _13033_ (.A(_06021_),
    .B(_06026_),
    .C(_06027_),
    .Y(_06029_));
 sky130_fd_sc_hd__and2_4 _13034_ (.A(_06028_),
    .B(_06029_),
    .X(loadstore_address[10]));
 sky130_fd_sc_hd__or2_1 _13035_ (.A(reg1_val[11]),
    .B(_05363_),
    .X(_06030_));
 sky130_fd_sc_hd__nand2_1 _13036_ (.A(reg1_val[11]),
    .B(_05363_),
    .Y(_06032_));
 sky130_fd_sc_hd__nand2_1 _13037_ (.A(_06030_),
    .B(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__a21o_1 _13038_ (.A1(_06025_),
    .A2(_06028_),
    .B1(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__nand3_1 _13039_ (.A(_06025_),
    .B(_06028_),
    .C(_06033_),
    .Y(_06035_));
 sky130_fd_sc_hd__and2_4 _13040_ (.A(_06034_),
    .B(_06035_),
    .X(loadstore_address[11]));
 sky130_fd_sc_hd__or2_1 _13041_ (.A(reg1_val[12]),
    .B(_04960_),
    .X(_06036_));
 sky130_fd_sc_hd__nand2_1 _13042_ (.A(reg1_val[12]),
    .B(_04960_),
    .Y(_06037_));
 sky130_fd_sc_hd__nand2_1 _13043_ (.A(_06036_),
    .B(_06037_),
    .Y(_06038_));
 sky130_fd_sc_hd__a21o_1 _13044_ (.A1(_06032_),
    .A2(_06034_),
    .B1(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__nand3_1 _13045_ (.A(_06032_),
    .B(_06034_),
    .C(_06038_),
    .Y(_06040_));
 sky130_fd_sc_hd__and2_4 _13046_ (.A(_06039_),
    .B(_06040_),
    .X(loadstore_address[12]));
 sky130_fd_sc_hd__or2_1 _13047_ (.A(reg1_val[13]),
    .B(_05189_),
    .X(_06042_));
 sky130_fd_sc_hd__nand2_1 _13048_ (.A(reg1_val[13]),
    .B(_05189_),
    .Y(_06043_));
 sky130_fd_sc_hd__nand2_1 _13049_ (.A(_06042_),
    .B(_06043_),
    .Y(_06044_));
 sky130_fd_sc_hd__a21o_1 _13050_ (.A1(_06037_),
    .A2(_06039_),
    .B1(_06044_),
    .X(_06045_));
 sky130_fd_sc_hd__nand3_1 _13051_ (.A(_06037_),
    .B(_06039_),
    .C(_06044_),
    .Y(_06046_));
 sky130_fd_sc_hd__and2_4 _13052_ (.A(_06045_),
    .B(_06046_),
    .X(loadstore_address[13]));
 sky130_fd_sc_hd__or2_1 _13053_ (.A(reg1_val[14]),
    .B(_05102_),
    .X(_06047_));
 sky130_fd_sc_hd__nand2_1 _13054_ (.A(reg1_val[14]),
    .B(_05102_),
    .Y(_06048_));
 sky130_fd_sc_hd__nand2_1 _13055_ (.A(_06047_),
    .B(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__a21o_1 _13056_ (.A1(_06043_),
    .A2(_06045_),
    .B1(_06049_),
    .X(_06051_));
 sky130_fd_sc_hd__nand3_1 _13057_ (.A(_06043_),
    .B(_06045_),
    .C(_06049_),
    .Y(_06052_));
 sky130_fd_sc_hd__and2_4 _13058_ (.A(_06051_),
    .B(_06052_),
    .X(loadstore_address[14]));
 sky130_fd_sc_hd__xnor2_2 _13059_ (.A(reg1_val[15]),
    .B(_05047_),
    .Y(_06053_));
 sky130_fd_sc_hd__a21oi_4 _13060_ (.A1(_06048_),
    .A2(_06051_),
    .B1(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__and3_2 _13061_ (.A(_06048_),
    .B(_06051_),
    .C(_06053_),
    .X(_06055_));
 sky130_fd_sc_hd__nor2_8 _13062_ (.A(_06054_),
    .B(_06055_),
    .Y(loadstore_address[15]));
 sky130_fd_sc_hd__nor2_1 _13063_ (.A(reg1_val[16]),
    .B(net264),
    .Y(_06056_));
 sky130_fd_sc_hd__and2_1 _13064_ (.A(reg1_val[16]),
    .B(net264),
    .X(_06057_));
 sky130_fd_sc_hd__or2_2 _13065_ (.A(_06056_),
    .B(_06057_),
    .X(_06058_));
 sky130_fd_sc_hd__a21oi_2 _13066_ (.A1(reg1_val[15]),
    .A2(_05047_),
    .B1(_06054_),
    .Y(_06060_));
 sky130_fd_sc_hd__or2_1 _13067_ (.A(_06058_),
    .B(_06060_),
    .X(_06061_));
 sky130_fd_sc_hd__xor2_4 _13068_ (.A(_06058_),
    .B(_06060_),
    .X(loadstore_address[16]));
 sky130_fd_sc_hd__nand2b_2 _13069_ (.A_N(_06057_),
    .B(_06061_),
    .Y(_06062_));
 sky130_fd_sc_hd__xnor2_4 _13070_ (.A(reg1_val[17]),
    .B(net264),
    .Y(_06063_));
 sky130_fd_sc_hd__xnor2_4 _13071_ (.A(_06062_),
    .B(_06063_),
    .Y(loadstore_address[17]));
 sky130_fd_sc_hd__or2_1 _13072_ (.A(reg1_val[18]),
    .B(net264),
    .X(_06064_));
 sky130_fd_sc_hd__nand2_1 _13073_ (.A(reg1_val[18]),
    .B(net264),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_2 _13074_ (.A(_06064_),
    .B(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__a2bb2o_2 _13075_ (.A1_N(_06061_),
    .A2_N(_06063_),
    .B1(net264),
    .B2(_00249_),
    .X(_06067_));
 sky130_fd_sc_hd__xnor2_4 _13076_ (.A(_06066_),
    .B(_06067_),
    .Y(loadstore_address[18]));
 sky130_fd_sc_hd__a21bo_1 _13077_ (.A1(_06064_),
    .A2(_06067_),
    .B1_N(_06065_),
    .X(_06069_));
 sky130_fd_sc_hd__xnor2_2 _13078_ (.A(reg1_val[19]),
    .B(net264),
    .Y(_06070_));
 sky130_fd_sc_hd__xnor2_4 _13079_ (.A(_06069_),
    .B(_06070_),
    .Y(loadstore_address[19]));
 sky130_fd_sc_hd__xnor2_2 _13080_ (.A(reg1_val[20]),
    .B(net264),
    .Y(_06071_));
 sky130_fd_sc_hd__or4_2 _13081_ (.A(_06061_),
    .B(_06063_),
    .C(_06066_),
    .D(_06070_),
    .X(_06072_));
 sky130_fd_sc_hd__nand2_2 _13082_ (.A(_04797_),
    .B(_00251_),
    .Y(_06073_));
 sky130_fd_sc_hd__a21oi_4 _13083_ (.A1(_06072_),
    .A2(_06073_),
    .B1(_06071_),
    .Y(_06074_));
 sky130_fd_sc_hd__and3_2 _13084_ (.A(_06071_),
    .B(_06072_),
    .C(_06073_),
    .X(_06075_));
 sky130_fd_sc_hd__nor2_8 _13085_ (.A(_06074_),
    .B(_06075_),
    .Y(loadstore_address[20]));
 sky130_fd_sc_hd__nor2_1 _13086_ (.A(reg1_val[21]),
    .B(net264),
    .Y(_06077_));
 sky130_fd_sc_hd__nand2_1 _13087_ (.A(reg1_val[21]),
    .B(net264),
    .Y(_06078_));
 sky130_fd_sc_hd__nand2b_2 _13088_ (.A_N(_06077_),
    .B(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__a21oi_4 _13089_ (.A1(reg1_val[20]),
    .A2(net264),
    .B1(_06074_),
    .Y(_06080_));
 sky130_fd_sc_hd__xor2_4 _13090_ (.A(_06079_),
    .B(_06080_),
    .X(loadstore_address[21]));
 sky130_fd_sc_hd__or2_1 _13091_ (.A(reg1_val[22]),
    .B(net264),
    .X(_06081_));
 sky130_fd_sc_hd__nand2_1 _13092_ (.A(reg1_val[22]),
    .B(net264),
    .Y(_06082_));
 sky130_fd_sc_hd__nand2_2 _13093_ (.A(_06081_),
    .B(_06082_),
    .Y(_06083_));
 sky130_fd_sc_hd__o21ai_4 _13094_ (.A1(_06077_),
    .A2(_06080_),
    .B1(_06078_),
    .Y(_06084_));
 sky130_fd_sc_hd__xnor2_4 _13095_ (.A(_06083_),
    .B(_06084_),
    .Y(loadstore_address[22]));
 sky130_fd_sc_hd__a21bo_1 _13096_ (.A1(_06081_),
    .A2(_06084_),
    .B1_N(_06082_),
    .X(_06086_));
 sky130_fd_sc_hd__xnor2_4 _13097_ (.A(reg1_val[23]),
    .B(net264),
    .Y(_06087_));
 sky130_fd_sc_hd__xnor2_4 _13098_ (.A(_06086_),
    .B(_06087_),
    .Y(loadstore_address[23]));
 sky130_fd_sc_hd__or2_1 _13099_ (.A(reg1_val[24]),
    .B(net265),
    .X(_06088_));
 sky130_fd_sc_hd__nand2_1 _13100_ (.A(reg1_val[24]),
    .B(net265),
    .Y(_06089_));
 sky130_fd_sc_hd__nand2_2 _13101_ (.A(_06088_),
    .B(_06089_),
    .Y(_06090_));
 sky130_fd_sc_hd__or4_1 _13102_ (.A(_06071_),
    .B(_06079_),
    .C(_06083_),
    .D(_06087_),
    .X(_06091_));
 sky130_fd_sc_hd__a2bb2o_2 _13103_ (.A1_N(_06072_),
    .A2_N(_06091_),
    .B1(net264),
    .B2(_00255_),
    .X(_06092_));
 sky130_fd_sc_hd__nand2b_1 _13104_ (.A_N(_06090_),
    .B(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__xnor2_4 _13105_ (.A(_06090_),
    .B(_06092_),
    .Y(loadstore_address[24]));
 sky130_fd_sc_hd__nand2_2 _13106_ (.A(_06089_),
    .B(_06093_),
    .Y(_06095_));
 sky130_fd_sc_hd__xnor2_2 _13107_ (.A(reg1_val[25]),
    .B(net265),
    .Y(_06096_));
 sky130_fd_sc_hd__xnor2_4 _13108_ (.A(_06095_),
    .B(_06096_),
    .Y(loadstore_address[25]));
 sky130_fd_sc_hd__or2_1 _13109_ (.A(reg1_val[26]),
    .B(net265),
    .X(_06097_));
 sky130_fd_sc_hd__nand2_1 _13110_ (.A(reg1_val[26]),
    .B(net265),
    .Y(_06098_));
 sky130_fd_sc_hd__nand2_2 _13111_ (.A(_06097_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__or2_1 _13112_ (.A(_06093_),
    .B(_06096_),
    .X(_06100_));
 sky130_fd_sc_hd__a21bo_2 _13113_ (.A1(net265),
    .A2(_00293_),
    .B1_N(_06100_),
    .X(_06101_));
 sky130_fd_sc_hd__xnor2_4 _13114_ (.A(_06099_),
    .B(_06101_),
    .Y(loadstore_address[26]));
 sky130_fd_sc_hd__a21bo_1 _13115_ (.A1(_06097_),
    .A2(_06101_),
    .B1_N(_06098_),
    .X(_06102_));
 sky130_fd_sc_hd__xnor2_2 _13116_ (.A(reg1_val[27]),
    .B(net265),
    .Y(_06104_));
 sky130_fd_sc_hd__xnor2_4 _13117_ (.A(_06102_),
    .B(_06104_),
    .Y(loadstore_address[27]));
 sky130_fd_sc_hd__or2_1 _13118_ (.A(reg1_val[28]),
    .B(net265),
    .X(_06105_));
 sky130_fd_sc_hd__nand2_1 _13119_ (.A(reg1_val[28]),
    .B(net265),
    .Y(_06106_));
 sky130_fd_sc_hd__nand2_2 _13120_ (.A(_06105_),
    .B(_06106_),
    .Y(_06107_));
 sky130_fd_sc_hd__or2_1 _13121_ (.A(_06099_),
    .B(_06104_),
    .X(_06108_));
 sky130_fd_sc_hd__a2bb2o_2 _13122_ (.A1_N(_06100_),
    .A2_N(_06108_),
    .B1(net265),
    .B2(_00294_),
    .X(_06109_));
 sky130_fd_sc_hd__xnor2_4 _13123_ (.A(_06107_),
    .B(_06109_),
    .Y(loadstore_address[28]));
 sky130_fd_sc_hd__nand2_1 _13124_ (.A(reg1_val[29]),
    .B(net265),
    .Y(_06110_));
 sky130_fd_sc_hd__or2_1 _13125_ (.A(reg1_val[29]),
    .B(net265),
    .X(_06111_));
 sky130_fd_sc_hd__nand2_2 _13126_ (.A(_06110_),
    .B(_06111_),
    .Y(_06113_));
 sky130_fd_sc_hd__a21bo_2 _13127_ (.A1(_06105_),
    .A2(_06109_),
    .B1_N(_06106_),
    .X(_06114_));
 sky130_fd_sc_hd__xnor2_4 _13128_ (.A(_06113_),
    .B(_06114_),
    .Y(loadstore_address[29]));
 sky130_fd_sc_hd__or2_1 _13129_ (.A(net288),
    .B(net264),
    .X(_06115_));
 sky130_fd_sc_hd__nand2_1 _13130_ (.A(reg1_val[30]),
    .B(net265),
    .Y(_06116_));
 sky130_fd_sc_hd__nand2_2 _13131_ (.A(_06115_),
    .B(_06116_),
    .Y(_06117_));
 sky130_fd_sc_hd__a21bo_2 _13132_ (.A1(_06111_),
    .A2(_06114_),
    .B1_N(_06110_),
    .X(_06118_));
 sky130_fd_sc_hd__xnor2_4 _13133_ (.A(_06117_),
    .B(_06118_),
    .Y(loadstore_address[30]));
 sky130_fd_sc_hd__a21boi_2 _13134_ (.A1(_06115_),
    .A2(_06118_),
    .B1_N(_06116_),
    .Y(_06119_));
 sky130_fd_sc_hd__xnor2_4 _13135_ (.A(_04598_),
    .B(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__xnor2_4 _13136_ (.A(net265),
    .B(_06120_),
    .Y(loadstore_address[31]));
 sky130_fd_sc_hd__and3_1 _13137_ (.A(net467),
    .B(net301),
    .C(net489),
    .X(_06122_));
 sky130_fd_sc_hd__nand3_1 _13138_ (.A(net441),
    .B(net313),
    .C(_06122_),
    .Y(_06123_));
 sky130_fd_sc_hd__nor2_1 _13139_ (.A(net249),
    .B(net490),
    .Y(_06124_));
 sky130_fd_sc_hd__nor3_1 _13140_ (.A(rst),
    .B(net188),
    .C(_06124_),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_1 _13141_ (.A(net255),
    .B(_06660_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand2_1 _13142_ (.A(net249),
    .B(_06659_),
    .Y(_06126_));
 sky130_fd_sc_hd__or2_1 _13143_ (.A(net315),
    .B(net166),
    .X(_06127_));
 sky130_fd_sc_hd__o211a_1 _13144_ (.A1(net61),
    .A2(net162),
    .B1(net316),
    .C1(net280),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_1 _13145_ (.A(net211),
    .B(net165),
    .Y(_06128_));
 sky130_fd_sc_hd__o211a_1 _13146_ (.A1(net311),
    .A2(net165),
    .B1(_06128_),
    .C1(net276),
    .X(_00002_));
 sky130_fd_sc_hd__nand2_1 _13147_ (.A(_00320_),
    .B(net165),
    .Y(_06130_));
 sky130_fd_sc_hd__o211a_1 _13148_ (.A1(net309),
    .A2(net165),
    .B1(_06130_),
    .C1(net273),
    .X(_00003_));
 sky130_fd_sc_hd__nand2_1 _13149_ (.A(net151),
    .B(net165),
    .Y(_06131_));
 sky130_fd_sc_hd__o211a_1 _13150_ (.A1(net307),
    .A2(net165),
    .B1(_06131_),
    .C1(net273),
    .X(_00004_));
 sky130_fd_sc_hd__nand2_1 _13151_ (.A(_00339_),
    .B(net165),
    .Y(_06132_));
 sky130_fd_sc_hd__o211a_1 _13152_ (.A1(net305),
    .A2(net165),
    .B1(_06132_),
    .C1(net274),
    .X(_00005_));
 sky130_fd_sc_hd__or2_1 _13153_ (.A(net381),
    .B(net165),
    .X(_06133_));
 sky130_fd_sc_hd__o211a_1 _13154_ (.A1(_00266_),
    .A2(net159),
    .B1(net382),
    .C1(net276),
    .X(_00006_));
 sky130_fd_sc_hd__or2_1 _13155_ (.A(net376),
    .B(net164),
    .X(_06134_));
 sky130_fd_sc_hd__o211a_1 _13156_ (.A1(_00287_),
    .A2(net163),
    .B1(net377),
    .C1(net276),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _13157_ (.A(net333),
    .B(net164),
    .X(_06136_));
 sky130_fd_sc_hd__o211a_1 _13158_ (.A1(_00476_),
    .A2(net163),
    .B1(net334),
    .C1(net276),
    .X(_00008_));
 sky130_fd_sc_hd__or2_1 _13159_ (.A(net371),
    .B(net165),
    .X(_06137_));
 sky130_fd_sc_hd__o211a_1 _13160_ (.A1(_00412_),
    .A2(net163),
    .B1(net372),
    .C1(net276),
    .X(_00009_));
 sky130_fd_sc_hd__or2_1 _13161_ (.A(net366),
    .B(net165),
    .X(_06138_));
 sky130_fd_sc_hd__o211a_1 _13162_ (.A1(_00414_),
    .A2(net159),
    .B1(net367),
    .C1(net276),
    .X(_00010_));
 sky130_fd_sc_hd__or2_1 _13163_ (.A(net409),
    .B(net164),
    .X(_06139_));
 sky130_fd_sc_hd__o211a_1 _13164_ (.A1(net122),
    .A2(net159),
    .B1(net410),
    .C1(net275),
    .X(_00011_));
 sky130_fd_sc_hd__or2_1 _13165_ (.A(net403),
    .B(net164),
    .X(_06140_));
 sky130_fd_sc_hd__o211a_1 _13166_ (.A1(net121),
    .A2(net159),
    .B1(net404),
    .C1(net274),
    .X(_00012_));
 sky130_fd_sc_hd__or2_1 _13167_ (.A(net360),
    .B(net164),
    .X(_06142_));
 sky130_fd_sc_hd__o211a_1 _13168_ (.A1(net114),
    .A2(net159),
    .B1(net361),
    .C1(net274),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _13169_ (.A(net349),
    .B(net165),
    .X(_06143_));
 sky130_fd_sc_hd__o211a_1 _13170_ (.A1(_00397_),
    .A2(net159),
    .B1(net350),
    .C1(net272),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _13171_ (.A(net355),
    .B(net164),
    .X(_06144_));
 sky130_fd_sc_hd__o211a_1 _13172_ (.A1(net81),
    .A2(net159),
    .B1(net356),
    .C1(net274),
    .X(_00015_));
 sky130_fd_sc_hd__or2_1 _13173_ (.A(net364),
    .B(net164),
    .X(_06145_));
 sky130_fd_sc_hd__o211a_1 _13174_ (.A1(net78),
    .A2(net159),
    .B1(net365),
    .C1(net274),
    .X(_00016_));
 sky130_fd_sc_hd__or2_1 _13175_ (.A(net388),
    .B(net164),
    .X(_06146_));
 sky130_fd_sc_hd__o211a_1 _13176_ (.A1(net73),
    .A2(net159),
    .B1(net389),
    .C1(net274),
    .X(_00017_));
 sky130_fd_sc_hd__or2_1 _13177_ (.A(net424),
    .B(net164),
    .X(_06148_));
 sky130_fd_sc_hd__o211a_1 _13178_ (.A1(net71),
    .A2(net159),
    .B1(net425),
    .C1(net275),
    .X(_00018_));
 sky130_fd_sc_hd__or2_1 _13179_ (.A(net353),
    .B(net164),
    .X(_06149_));
 sky130_fd_sc_hd__o211a_1 _13180_ (.A1(net102),
    .A2(net159),
    .B1(net354),
    .C1(net275),
    .X(_00019_));
 sky130_fd_sc_hd__or2_1 _13181_ (.A(net335),
    .B(net164),
    .X(_06150_));
 sky130_fd_sc_hd__o211a_1 _13182_ (.A1(net101),
    .A2(net159),
    .B1(net336),
    .C1(net275),
    .X(_00020_));
 sky130_fd_sc_hd__or2_1 _13183_ (.A(net414),
    .B(net164),
    .X(_06151_));
 sky130_fd_sc_hd__o211a_1 _13184_ (.A1(_00203_),
    .A2(net159),
    .B1(net415),
    .C1(net275),
    .X(_00021_));
 sky130_fd_sc_hd__or2_1 _13185_ (.A(net432),
    .B(net164),
    .X(_06152_));
 sky130_fd_sc_hd__o211a_1 _13186_ (.A1(_00208_),
    .A2(net159),
    .B1(net433),
    .C1(net275),
    .X(_00022_));
 sky130_fd_sc_hd__or2_1 _13187_ (.A(net383),
    .B(net164),
    .X(_06154_));
 sky130_fd_sc_hd__o211a_1 _13188_ (.A1(_06725_),
    .A2(net163),
    .B1(net384),
    .C1(net277),
    .X(_00023_));
 sky130_fd_sc_hd__or2_1 _13189_ (.A(net346),
    .B(net164),
    .X(_06155_));
 sky130_fd_sc_hd__o211a_1 _13190_ (.A1(net55),
    .A2(net163),
    .B1(net347),
    .C1(net277),
    .X(_00024_));
 sky130_fd_sc_hd__or2_1 _13191_ (.A(net401),
    .B(net164),
    .X(_06156_));
 sky130_fd_sc_hd__o211a_1 _13192_ (.A1(_00150_),
    .A2(net159),
    .B1(net402),
    .C1(net277),
    .X(_00025_));
 sky130_fd_sc_hd__or2_1 _13193_ (.A(net416),
    .B(net165),
    .X(_06157_));
 sky130_fd_sc_hd__o211a_1 _13194_ (.A1(_00161_),
    .A2(net159),
    .B1(net417),
    .C1(net277),
    .X(_00026_));
 sky130_fd_sc_hd__or2_1 _13195_ (.A(net337),
    .B(net166),
    .X(_06158_));
 sky130_fd_sc_hd__o211a_1 _13196_ (.A1(_00144_),
    .A2(net163),
    .B1(net338),
    .C1(net277),
    .X(_00027_));
 sky130_fd_sc_hd__or2_1 _13197_ (.A(net344),
    .B(net166),
    .X(_06160_));
 sky130_fd_sc_hd__o211a_1 _13198_ (.A1(_00136_),
    .A2(net162),
    .B1(net345),
    .C1(net281),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _13199_ (.A(net340),
    .B(net166),
    .X(_06161_));
 sky130_fd_sc_hd__o211a_1 _13200_ (.A1(_00177_),
    .A2(net162),
    .B1(net341),
    .C1(net280),
    .X(_00029_));
 sky130_fd_sc_hd__or2_1 _13201_ (.A(net326),
    .B(net166),
    .X(_06162_));
 sky130_fd_sc_hd__o211a_1 _13202_ (.A1(_00516_),
    .A2(net162),
    .B1(net327),
    .C1(net280),
    .X(_00030_));
 sky130_fd_sc_hd__or2_1 _13203_ (.A(net328),
    .B(net166),
    .X(_06163_));
 sky130_fd_sc_hd__o211a_1 _13204_ (.A1(_00812_),
    .A2(net162),
    .B1(net329),
    .C1(net280),
    .X(_00031_));
 sky130_fd_sc_hd__or2_1 _13205_ (.A(net342),
    .B(net166),
    .X(_06164_));
 sky130_fd_sc_hd__o211a_1 _13206_ (.A1(_02065_),
    .A2(net162),
    .B1(net343),
    .C1(net280),
    .X(_00032_));
 sky130_fd_sc_hd__or2_1 _13207_ (.A(net470),
    .B(net166),
    .X(_06166_));
 sky130_fd_sc_hd__o211a_1 _13208_ (.A1(net7),
    .A2(net162),
    .B1(net471),
    .C1(net280),
    .X(_00033_));
 sky130_fd_sc_hd__nand2b_1 _13209_ (.A_N(net342),
    .B(net566),
    .Y(_06167_));
 sky130_fd_sc_hd__nand2b_1 _13210_ (.A_N(net566),
    .B(net342),
    .Y(_06168_));
 sky130_fd_sc_hd__nand2_1 _13211_ (.A(_06167_),
    .B(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__and2b_1 _13212_ (.A_N(net328),
    .B(net545),
    .X(_06170_));
 sky130_fd_sc_hd__and2b_1 _13213_ (.A_N(net545),
    .B(net328),
    .X(_06171_));
 sky130_fd_sc_hd__nor2_1 _13214_ (.A(_06170_),
    .B(_06171_),
    .Y(_06172_));
 sky130_fd_sc_hd__and2b_1 _13215_ (.A_N(net326),
    .B(net547),
    .X(_06173_));
 sky130_fd_sc_hd__and2b_1 _13216_ (.A_N(\div_shifter[59] ),
    .B(net326),
    .X(_06175_));
 sky130_fd_sc_hd__nor2_1 _13217_ (.A(_06173_),
    .B(_06175_),
    .Y(_06176_));
 sky130_fd_sc_hd__and2b_1 _13218_ (.A_N(net340),
    .B(\div_shifter[58] ),
    .X(_06177_));
 sky130_fd_sc_hd__nand2b_1 _13219_ (.A_N(\div_shifter[58] ),
    .B(net340),
    .Y(_06178_));
 sky130_fd_sc_hd__and2b_1 _13220_ (.A_N(net344),
    .B(\div_shifter[57] ),
    .X(_06179_));
 sky130_fd_sc_hd__and2b_1 _13221_ (.A_N(\div_shifter[57] ),
    .B(net344),
    .X(_06180_));
 sky130_fd_sc_hd__nor2_1 _13222_ (.A(_06179_),
    .B(_06180_),
    .Y(_06181_));
 sky130_fd_sc_hd__and2b_1 _13223_ (.A_N(net337),
    .B(net567),
    .X(_06182_));
 sky130_fd_sc_hd__and2b_1 _13224_ (.A_N(net567),
    .B(net337),
    .X(_06183_));
 sky130_fd_sc_hd__nor2_1 _13225_ (.A(_06182_),
    .B(_06183_),
    .Y(_06184_));
 sky130_fd_sc_hd__and2b_1 _13226_ (.A_N(net416),
    .B(\div_shifter[55] ),
    .X(_06186_));
 sky130_fd_sc_hd__nand2b_1 _13227_ (.A_N(\div_shifter[55] ),
    .B(net416),
    .Y(_06187_));
 sky130_fd_sc_hd__nand2b_1 _13228_ (.A_N(_06186_),
    .B(_06187_),
    .Y(_06188_));
 sky130_fd_sc_hd__and2b_1 _13229_ (.A_N(net401),
    .B(net553),
    .X(_06189_));
 sky130_fd_sc_hd__nand2b_1 _13230_ (.A_N(net553),
    .B(net401),
    .Y(_06190_));
 sky130_fd_sc_hd__and2b_1 _13231_ (.A_N(net346),
    .B(net564),
    .X(_06191_));
 sky130_fd_sc_hd__and2b_1 _13232_ (.A_N(net564),
    .B(net346),
    .X(_06192_));
 sky130_fd_sc_hd__nor2_1 _13233_ (.A(_06191_),
    .B(_06192_),
    .Y(_06193_));
 sky130_fd_sc_hd__and2b_1 _13234_ (.A_N(net383),
    .B(\div_shifter[52] ),
    .X(_06194_));
 sky130_fd_sc_hd__and2b_1 _13235_ (.A_N(\div_shifter[52] ),
    .B(net383),
    .X(_06195_));
 sky130_fd_sc_hd__nor2_1 _13236_ (.A(_06194_),
    .B(_06195_),
    .Y(_06197_));
 sky130_fd_sc_hd__and2b_1 _13237_ (.A_N(net432),
    .B(net559),
    .X(_06198_));
 sky130_fd_sc_hd__nand2b_1 _13238_ (.A_N(net559),
    .B(net432),
    .Y(_06199_));
 sky130_fd_sc_hd__nand2b_1 _13239_ (.A_N(_06198_),
    .B(_06199_),
    .Y(_06200_));
 sky130_fd_sc_hd__and2b_1 _13240_ (.A_N(net414),
    .B(net557),
    .X(_06201_));
 sky130_fd_sc_hd__nand2b_1 _13241_ (.A_N(net557),
    .B(net414),
    .Y(_06202_));
 sky130_fd_sc_hd__and2b_1 _13242_ (.A_N(net335),
    .B(net555),
    .X(_06203_));
 sky130_fd_sc_hd__and2b_1 _13243_ (.A_N(net555),
    .B(net335),
    .X(_06204_));
 sky130_fd_sc_hd__nor2_1 _13244_ (.A(_06203_),
    .B(_06204_),
    .Y(_06205_));
 sky130_fd_sc_hd__and2b_1 _13245_ (.A_N(net353),
    .B(\div_shifter[48] ),
    .X(_06206_));
 sky130_fd_sc_hd__and2b_1 _13246_ (.A_N(\div_shifter[48] ),
    .B(net353),
    .X(_06208_));
 sky130_fd_sc_hd__nor2_1 _13247_ (.A(_06206_),
    .B(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__and2b_1 _13248_ (.A_N(net424),
    .B(\div_shifter[47] ),
    .X(_06210_));
 sky130_fd_sc_hd__nand2b_1 _13249_ (.A_N(\div_shifter[47] ),
    .B(net424),
    .Y(_06211_));
 sky130_fd_sc_hd__nand2b_1 _13250_ (.A_N(_06210_),
    .B(_06211_),
    .Y(_06212_));
 sky130_fd_sc_hd__and2b_1 _13251_ (.A_N(net388),
    .B(net549),
    .X(_06213_));
 sky130_fd_sc_hd__nand2b_1 _13252_ (.A_N(net549),
    .B(net388),
    .Y(_06214_));
 sky130_fd_sc_hd__and2b_1 _13253_ (.A_N(net364),
    .B(net587),
    .X(_06215_));
 sky130_fd_sc_hd__nand2b_1 _13254_ (.A_N(net587),
    .B(net364),
    .Y(_06216_));
 sky130_fd_sc_hd__and2b_1 _13255_ (.A_N(net355),
    .B(net569),
    .X(_06217_));
 sky130_fd_sc_hd__nand2b_1 _13256_ (.A_N(net569),
    .B(net355),
    .Y(_06219_));
 sky130_fd_sc_hd__and2b_1 _13257_ (.A_N(net349),
    .B(\div_shifter[43] ),
    .X(_06220_));
 sky130_fd_sc_hd__nand2b_1 _13258_ (.A_N(\div_shifter[43] ),
    .B(net349),
    .Y(_06221_));
 sky130_fd_sc_hd__and2b_1 _13259_ (.A_N(net360),
    .B(net578),
    .X(_06222_));
 sky130_fd_sc_hd__nand2b_1 _13260_ (.A_N(net578),
    .B(net360),
    .Y(_06223_));
 sky130_fd_sc_hd__and2b_1 _13261_ (.A_N(net403),
    .B(net551),
    .X(_06224_));
 sky130_fd_sc_hd__nand2b_1 _13262_ (.A_N(net551),
    .B(net403),
    .Y(_06225_));
 sky130_fd_sc_hd__and2b_1 _13263_ (.A_N(net409),
    .B(\div_shifter[40] ),
    .X(_06226_));
 sky130_fd_sc_hd__nand2b_1 _13264_ (.A_N(\div_shifter[40] ),
    .B(net409),
    .Y(_06227_));
 sky130_fd_sc_hd__and2b_1 _13265_ (.A_N(net366),
    .B(net574),
    .X(_06228_));
 sky130_fd_sc_hd__nand2b_1 _13266_ (.A_N(net574),
    .B(net366),
    .Y(_06230_));
 sky130_fd_sc_hd__and2b_1 _13267_ (.A_N(net371),
    .B(net585),
    .X(_06231_));
 sky130_fd_sc_hd__nand2b_1 _13268_ (.A_N(net585),
    .B(net371),
    .Y(_06232_));
 sky130_fd_sc_hd__and2b_1 _13269_ (.A_N(net333),
    .B(\div_shifter[37] ),
    .X(_06233_));
 sky130_fd_sc_hd__nand2b_1 _13270_ (.A_N(\div_shifter[37] ),
    .B(net333),
    .Y(_06234_));
 sky130_fd_sc_hd__and2b_1 _13271_ (.A_N(net376),
    .B(net581),
    .X(_06235_));
 sky130_fd_sc_hd__nand2b_1 _13272_ (.A_N(net581),
    .B(net376),
    .Y(_06236_));
 sky130_fd_sc_hd__nand2b_1 _13273_ (.A_N(_06235_),
    .B(_06236_),
    .Y(_06237_));
 sky130_fd_sc_hd__and2b_1 _13274_ (.A_N(net381),
    .B(net562),
    .X(_06238_));
 sky130_fd_sc_hd__nand2b_1 _13275_ (.A_N(net562),
    .B(net381),
    .Y(_06239_));
 sky130_fd_sc_hd__nand2b_1 _13276_ (.A_N(_06238_),
    .B(_06239_),
    .Y(_06241_));
 sky130_fd_sc_hd__and2b_1 _13277_ (.A_N(net305),
    .B(\div_shifter[34] ),
    .X(_06242_));
 sky130_fd_sc_hd__nand2b_1 _13278_ (.A_N(\div_shifter[34] ),
    .B(net305),
    .Y(_06243_));
 sky130_fd_sc_hd__and2b_1 _13279_ (.A_N(net307),
    .B(net560),
    .X(_06244_));
 sky130_fd_sc_hd__nand2b_1 _13280_ (.A_N(net560),
    .B(net307),
    .Y(_06245_));
 sky130_fd_sc_hd__nand2b_1 _13281_ (.A_N(net309),
    .B(net543),
    .Y(_06246_));
 sky130_fd_sc_hd__xor2_1 _13282_ (.A(net543),
    .B(net309),
    .X(_06247_));
 sky130_fd_sc_hd__and2b_1 _13283_ (.A_N(\div_shifter[31] ),
    .B(net311),
    .X(_06248_));
 sky130_fd_sc_hd__o21ai_1 _13284_ (.A1(_06247_),
    .A2(_06248_),
    .B1(_06246_),
    .Y(_06249_));
 sky130_fd_sc_hd__a21o_1 _13285_ (.A1(_06245_),
    .A2(_06249_),
    .B1(_06244_),
    .X(_06250_));
 sky130_fd_sc_hd__a21o_1 _13286_ (.A1(_06243_),
    .A2(_06250_),
    .B1(_06242_),
    .X(_06252_));
 sky130_fd_sc_hd__a21o_1 _13287_ (.A1(_06239_),
    .A2(_06252_),
    .B1(_06238_),
    .X(_06253_));
 sky130_fd_sc_hd__a21o_1 _13288_ (.A1(_06236_),
    .A2(_06253_),
    .B1(_06235_),
    .X(_06254_));
 sky130_fd_sc_hd__a21o_1 _13289_ (.A1(_06234_),
    .A2(_06254_),
    .B1(_06233_),
    .X(_06255_));
 sky130_fd_sc_hd__a21o_1 _13290_ (.A1(_06232_),
    .A2(_06255_),
    .B1(_06231_),
    .X(_06256_));
 sky130_fd_sc_hd__a21o_1 _13291_ (.A1(_06230_),
    .A2(_06256_),
    .B1(_06228_),
    .X(_06257_));
 sky130_fd_sc_hd__a21o_1 _13292_ (.A1(_06227_),
    .A2(_06257_),
    .B1(_06226_),
    .X(_06258_));
 sky130_fd_sc_hd__a21o_1 _13293_ (.A1(_06225_),
    .A2(_06258_),
    .B1(_06224_),
    .X(_06259_));
 sky130_fd_sc_hd__a21o_1 _13294_ (.A1(_06223_),
    .A2(_06259_),
    .B1(_06222_),
    .X(_06260_));
 sky130_fd_sc_hd__a21o_1 _13295_ (.A1(_06221_),
    .A2(_06260_),
    .B1(_06220_),
    .X(_06261_));
 sky130_fd_sc_hd__a21o_1 _13296_ (.A1(_06219_),
    .A2(_06261_),
    .B1(_06217_),
    .X(_06263_));
 sky130_fd_sc_hd__a21o_1 _13297_ (.A1(_06216_),
    .A2(_06263_),
    .B1(_06215_),
    .X(_06264_));
 sky130_fd_sc_hd__a21o_1 _13298_ (.A1(_06214_),
    .A2(_06264_),
    .B1(_06213_),
    .X(_06265_));
 sky130_fd_sc_hd__a21o_1 _13299_ (.A1(_06211_),
    .A2(_06265_),
    .B1(_06210_),
    .X(_06266_));
 sky130_fd_sc_hd__a21oi_1 _13300_ (.A1(_06209_),
    .A2(_06266_),
    .B1(_06206_),
    .Y(_06267_));
 sky130_fd_sc_hd__o21bai_1 _13301_ (.A1(_06204_),
    .A2(_06267_),
    .B1_N(_06203_),
    .Y(_06268_));
 sky130_fd_sc_hd__a21o_1 _13302_ (.A1(_06202_),
    .A2(_06268_),
    .B1(_06201_),
    .X(_06269_));
 sky130_fd_sc_hd__a21o_1 _13303_ (.A1(_06199_),
    .A2(_06269_),
    .B1(_06198_),
    .X(_06270_));
 sky130_fd_sc_hd__a21oi_1 _13304_ (.A1(_06197_),
    .A2(_06270_),
    .B1(_06194_),
    .Y(_06271_));
 sky130_fd_sc_hd__o21bai_1 _13305_ (.A1(_06192_),
    .A2(_06271_),
    .B1_N(_06191_),
    .Y(_06272_));
 sky130_fd_sc_hd__a21o_1 _13306_ (.A1(_06190_),
    .A2(_06272_),
    .B1(_06189_),
    .X(_06274_));
 sky130_fd_sc_hd__a21o_1 _13307_ (.A1(_06187_),
    .A2(_06274_),
    .B1(_06186_),
    .X(_06275_));
 sky130_fd_sc_hd__a21oi_2 _13308_ (.A1(_06184_),
    .A2(_06275_),
    .B1(_06182_),
    .Y(_06276_));
 sky130_fd_sc_hd__o21bai_2 _13309_ (.A1(_06180_),
    .A2(_06276_),
    .B1_N(_06179_),
    .Y(_06277_));
 sky130_fd_sc_hd__a21oi_1 _13310_ (.A1(_06178_),
    .A2(_06277_),
    .B1(_06177_),
    .Y(_06278_));
 sky130_fd_sc_hd__and2b_1 _13311_ (.A_N(_06278_),
    .B(_06176_),
    .X(_06279_));
 sky130_fd_sc_hd__o21a_1 _13312_ (.A1(_06173_),
    .A2(_06279_),
    .B1(_06172_),
    .X(_06280_));
 sky130_fd_sc_hd__nor2_1 _13313_ (.A(_06170_),
    .B(_06280_),
    .Y(_06281_));
 sky130_fd_sc_hd__o21ai_1 _13314_ (.A1(_06169_),
    .A2(_06281_),
    .B1(_06167_),
    .Y(_06282_));
 sky130_fd_sc_hd__and2b_1 _13315_ (.A_N(net470),
    .B(net531),
    .X(_06283_));
 sky130_fd_sc_hd__nand2b_1 _13316_ (.A_N(net531),
    .B(net470),
    .Y(_06285_));
 sky130_fd_sc_hd__a21o_1 _13317_ (.A1(_06282_),
    .A2(_06285_),
    .B1(_06283_),
    .X(_06286_));
 sky130_fd_sc_hd__a22o_1 _13318_ (.A1(net486),
    .A2(net185),
    .B1(net1),
    .B2(net251),
    .X(_06287_));
 sky130_fd_sc_hd__and2_1 _13319_ (.A(net273),
    .B(_06287_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _13320_ (.A1(net486),
    .A2(net251),
    .B1(net185),
    .B2(\div_res[1] ),
    .X(_06288_));
 sky130_fd_sc_hd__and2_1 _13321_ (.A(net273),
    .B(net487),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_1 _13322_ (.A1(\div_res[1] ),
    .A2(net251),
    .B1(net185),
    .B2(net541),
    .X(_06289_));
 sky130_fd_sc_hd__and2_1 _13323_ (.A(net273),
    .B(net542),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_1 _13324_ (.A1(\div_res[2] ),
    .A2(net251),
    .B1(net185),
    .B2(net524),
    .X(_06290_));
 sky130_fd_sc_hd__and2_1 _13325_ (.A(net273),
    .B(net525),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _13326_ (.A1(net524),
    .A2(net251),
    .B1(net185),
    .B2(net536),
    .X(_06292_));
 sky130_fd_sc_hd__and2_1 _13327_ (.A(net273),
    .B(net537),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _13328_ (.A1(\div_res[4] ),
    .A2(net250),
    .B1(net184),
    .B2(net480),
    .X(_06293_));
 sky130_fd_sc_hd__and2_1 _13329_ (.A(net272),
    .B(net481),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_1 _13330_ (.A1(net480),
    .A2(net250),
    .B1(net184),
    .B2(net520),
    .X(_06294_));
 sky130_fd_sc_hd__and2_1 _13331_ (.A(net272),
    .B(net521),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_1 _13332_ (.A1(net520),
    .A2(net250),
    .B1(net184),
    .B2(net478),
    .X(_06295_));
 sky130_fd_sc_hd__and2_1 _13333_ (.A(net272),
    .B(_06295_),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_1 _13334_ (.A1(net478),
    .A2(net250),
    .B1(net184),
    .B2(net461),
    .X(_06296_));
 sky130_fd_sc_hd__and2_1 _13335_ (.A(net272),
    .B(net479),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_1 _13336_ (.A1(net461),
    .A2(net250),
    .B1(net184),
    .B2(\div_res[9] ),
    .X(_06298_));
 sky130_fd_sc_hd__and2_1 _13337_ (.A(net272),
    .B(net462),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_1 _13338_ (.A1(net538),
    .A2(net250),
    .B1(net184),
    .B2(\div_res[10] ),
    .X(_06299_));
 sky130_fd_sc_hd__and2_1 _13339_ (.A(net272),
    .B(net539),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_1 _13340_ (.A1(\div_res[10] ),
    .A2(net250),
    .B1(net184),
    .B2(net507),
    .X(_06300_));
 sky130_fd_sc_hd__and2_1 _13341_ (.A(net272),
    .B(net508),
    .X(_00045_));
 sky130_fd_sc_hd__a22o_1 _13342_ (.A1(net507),
    .A2(net250),
    .B1(net184),
    .B2(net512),
    .X(_06301_));
 sky130_fd_sc_hd__and2_1 _13343_ (.A(net272),
    .B(net513),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _13344_ (.A1(net512),
    .A2(net250),
    .B1(net184),
    .B2(net533),
    .X(_06302_));
 sky130_fd_sc_hd__and2_1 _13345_ (.A(net273),
    .B(net534),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _13346_ (.A1(net595),
    .A2(net250),
    .B1(net184),
    .B2(net491),
    .X(_06304_));
 sky130_fd_sc_hd__and2_1 _13347_ (.A(net272),
    .B(net492),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _13348_ (.A1(net491),
    .A2(net250),
    .B1(net184),
    .B2(net493),
    .X(_06305_));
 sky130_fd_sc_hd__and2_1 _13349_ (.A(net272),
    .B(net494),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _13350_ (.A1(net493),
    .A2(net251),
    .B1(net185),
    .B2(net529),
    .X(_06306_));
 sky130_fd_sc_hd__and2_1 _13351_ (.A(net272),
    .B(net530),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_1 _13352_ (.A1(\div_res[16] ),
    .A2(net250),
    .B1(net184),
    .B2(net498),
    .X(_06307_));
 sky130_fd_sc_hd__and2_1 _13353_ (.A(net272),
    .B(net499),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_1 _13354_ (.A1(net498),
    .A2(net250),
    .B1(net185),
    .B2(net483),
    .X(_06308_));
 sky130_fd_sc_hd__and2_1 _13355_ (.A(net272),
    .B(net502),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_1 _13356_ (.A1(net483),
    .A2(net250),
    .B1(net184),
    .B2(\div_res[19] ),
    .X(_06310_));
 sky130_fd_sc_hd__and2_1 _13357_ (.A(net272),
    .B(net484),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_1 _13358_ (.A1(\div_res[19] ),
    .A2(net251),
    .B1(net184),
    .B2(net475),
    .X(_06311_));
 sky130_fd_sc_hd__and2_1 _13359_ (.A(net272),
    .B(net476),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_1 _13360_ (.A1(net475),
    .A2(net251),
    .B1(net185),
    .B2(net472),
    .X(_06312_));
 sky130_fd_sc_hd__and2_1 _13361_ (.A(net274),
    .B(net511),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_1 _13362_ (.A1(net472),
    .A2(net252),
    .B1(net186),
    .B2(\div_res[22] ),
    .X(_06313_));
 sky130_fd_sc_hd__and2_1 _13363_ (.A(net274),
    .B(net473),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_1 _13364_ (.A1(\div_res[22] ),
    .A2(net252),
    .B1(net186),
    .B2(net503),
    .X(_06314_));
 sky130_fd_sc_hd__and2_1 _13365_ (.A(net274),
    .B(net504),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _13366_ (.A1(net503),
    .A2(net252),
    .B1(net187),
    .B2(net514),
    .X(_06316_));
 sky130_fd_sc_hd__and2_1 _13367_ (.A(net276),
    .B(net528),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _13368_ (.A1(net514),
    .A2(net253),
    .B1(net187),
    .B2(net505),
    .X(_06317_));
 sky130_fd_sc_hd__and2_1 _13369_ (.A(net276),
    .B(net515),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _13370_ (.A1(net505),
    .A2(net253),
    .B1(net188),
    .B2(net464),
    .X(_06318_));
 sky130_fd_sc_hd__and2_1 _13371_ (.A(net276),
    .B(net506),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_1 _13372_ (.A1(net464),
    .A2(net252),
    .B1(net188),
    .B2(\div_res[27] ),
    .X(_06319_));
 sky130_fd_sc_hd__and2_1 _13373_ (.A(net276),
    .B(net465),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_1 _13374_ (.A1(\div_res[27] ),
    .A2(net254),
    .B1(net188),
    .B2(net517),
    .X(_06320_));
 sky130_fd_sc_hd__and2_1 _13375_ (.A(net276),
    .B(net518),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _13376_ (.A1(\div_res[28] ),
    .A2(net254),
    .B1(net188),
    .B2(net495),
    .X(_06322_));
 sky130_fd_sc_hd__and2_1 _13377_ (.A(net280),
    .B(net496),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_1 _13378_ (.A1(net495),
    .A2(net254),
    .B1(net188),
    .B2(net522),
    .X(_06323_));
 sky130_fd_sc_hd__and2_1 _13379_ (.A(net280),
    .B(net523),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_1 _13380_ (.A1(\div_res[30] ),
    .A2(net254),
    .B1(net188),
    .B2(net452),
    .X(_06324_));
 sky130_fd_sc_hd__and2_1 _13381_ (.A(net280),
    .B(net453),
    .X(_00065_));
 sky130_fd_sc_hd__a22o_1 _13382_ (.A1(net447),
    .A2(_06661_),
    .B1(net166),
    .B2(net292),
    .X(_06325_));
 sky130_fd_sc_hd__and2_1 _13383_ (.A(net278),
    .B(net448),
    .X(_00066_));
 sky130_fd_sc_hd__o221a_1 _13384_ (.A1(net447),
    .A2(net248),
    .B1(net199),
    .B2(net160),
    .C1(net278),
    .X(_06326_));
 sky130_fd_sc_hd__o21a_1 _13385_ (.A1(net299),
    .A2(net183),
    .B1(_06326_),
    .X(_00067_));
 sky130_fd_sc_hd__o221a_1 _13386_ (.A1(net299),
    .A2(net248),
    .B1(net183),
    .B2(net374),
    .C1(net278),
    .X(_06328_));
 sky130_fd_sc_hd__o21a_1 _13387_ (.A1(_00153_),
    .A2(net160),
    .B1(net375),
    .X(_00068_));
 sky130_fd_sc_hd__o221a_1 _13388_ (.A1(net374),
    .A2(net248),
    .B1(net182),
    .B2(net399),
    .C1(net278),
    .X(_06329_));
 sky130_fd_sc_hd__o21a_1 _13389_ (.A1(net200),
    .A2(net160),
    .B1(net400),
    .X(_00069_));
 sky130_fd_sc_hd__o221a_1 _13390_ (.A1(net399),
    .A2(net248),
    .B1(net182),
    .B2(net426),
    .C1(net278),
    .X(_06330_));
 sky130_fd_sc_hd__o21a_1 _13391_ (.A1(_06696_),
    .A2(net160),
    .B1(net427),
    .X(_00070_));
 sky130_fd_sc_hd__o221a_1 _13392_ (.A1(\div_shifter[4] ),
    .A2(net248),
    .B1(net182),
    .B2(net396),
    .C1(net279),
    .X(_06331_));
 sky130_fd_sc_hd__o21a_1 _13393_ (.A1(net179),
    .A2(net160),
    .B1(net397),
    .X(_00071_));
 sky130_fd_sc_hd__o221a_1 _13394_ (.A1(net396),
    .A2(net248),
    .B1(net182),
    .B2(net459),
    .C1(net278),
    .X(_06332_));
 sky130_fd_sc_hd__a21boi_1 _13395_ (.A1(_00192_),
    .A2(net166),
    .B1_N(net460),
    .Y(_00072_));
 sky130_fd_sc_hd__a21oi_1 _13396_ (.A1(_04401_),
    .A2(net255),
    .B1(rst),
    .Y(_06334_));
 sky130_fd_sc_hd__o221a_1 _13397_ (.A1(net303),
    .A2(net182),
    .B1(_00187_),
    .B2(net160),
    .C1(_06334_),
    .X(_00073_));
 sky130_fd_sc_hd__o221a_1 _13398_ (.A1(net303),
    .A2(net248),
    .B1(net182),
    .B2(net362),
    .C1(net278),
    .X(_06335_));
 sky130_fd_sc_hd__o21a_1 _13399_ (.A1(_00223_),
    .A2(net160),
    .B1(net387),
    .X(_00074_));
 sky130_fd_sc_hd__o221a_1 _13400_ (.A1(net362),
    .A2(net248),
    .B1(net182),
    .B2(net317),
    .C1(net278),
    .X(_06336_));
 sky130_fd_sc_hd__o21a_1 _13401_ (.A1(net155),
    .A2(net160),
    .B1(net363),
    .X(_00075_));
 sky130_fd_sc_hd__o221a_1 _13402_ (.A1(net317),
    .A2(net248),
    .B1(net182),
    .B2(\div_shifter[10] ),
    .C1(net278),
    .X(_06337_));
 sky130_fd_sc_hd__o21a_1 _13403_ (.A1(_00492_),
    .A2(net160),
    .B1(net318),
    .X(_00076_));
 sky130_fd_sc_hd__o221a_1 _13404_ (.A1(net455),
    .A2(net248),
    .B1(net182),
    .B2(net418),
    .C1(net278),
    .X(_06338_));
 sky130_fd_sc_hd__o21a_1 _13405_ (.A1(net145),
    .A2(net161),
    .B1(net456),
    .X(_00077_));
 sky130_fd_sc_hd__o221a_1 _13406_ (.A1(net418),
    .A2(net248),
    .B1(net182),
    .B2(\div_shifter[12] ),
    .C1(net278),
    .X(_06340_));
 sky130_fd_sc_hd__o21a_1 _13407_ (.A1(_00456_),
    .A2(net160),
    .B1(net419),
    .X(_00078_));
 sky130_fd_sc_hd__o221a_1 _13408_ (.A1(\div_shifter[12] ),
    .A2(net248),
    .B1(net182),
    .B2(net390),
    .C1(net278),
    .X(_06341_));
 sky130_fd_sc_hd__o21a_1 _13409_ (.A1(net108),
    .A2(net160),
    .B1(net391),
    .X(_00079_));
 sky130_fd_sc_hd__o221a_1 _13410_ (.A1(net390),
    .A2(net248),
    .B1(net182),
    .B2(net430),
    .C1(net278),
    .X(_06342_));
 sky130_fd_sc_hd__o21a_1 _13411_ (.A1(_00436_),
    .A2(net160),
    .B1(net431),
    .X(_00080_));
 sky130_fd_sc_hd__o221a_1 _13412_ (.A1(net430),
    .A2(net248),
    .B1(net182),
    .B2(net405),
    .C1(net279),
    .X(_06343_));
 sky130_fd_sc_hd__o21a_1 _13413_ (.A1(net117),
    .A2(net160),
    .B1(net435),
    .X(_00081_));
 sky130_fd_sc_hd__o221a_1 _13414_ (.A1(net405),
    .A2(net248),
    .B1(net182),
    .B2(net320),
    .C1(net278),
    .X(_06344_));
 sky130_fd_sc_hd__o21a_1 _13415_ (.A1(_00383_),
    .A2(net160),
    .B1(net406),
    .X(_00082_));
 sky130_fd_sc_hd__o221a_1 _13416_ (.A1(net320),
    .A2(net248),
    .B1(net182),
    .B2(\div_shifter[17] ),
    .C1(net278),
    .X(_06346_));
 sky130_fd_sc_hd__o21a_1 _13417_ (.A1(net87),
    .A2(net160),
    .B1(net321),
    .X(_00083_));
 sky130_fd_sc_hd__o221a_1 _13418_ (.A1(\div_shifter[17] ),
    .A2(net249),
    .B1(net183),
    .B2(net449),
    .C1(net278),
    .X(_06347_));
 sky130_fd_sc_hd__o21a_1 _13419_ (.A1(_00363_),
    .A2(net160),
    .B1(net450),
    .X(_00084_));
 sky130_fd_sc_hd__o221a_1 _13420_ (.A1(\div_shifter[18] ),
    .A2(net249),
    .B1(net182),
    .B2(net411),
    .C1(net279),
    .X(_06348_));
 sky130_fd_sc_hd__o21a_1 _13421_ (.A1(net89),
    .A2(net161),
    .B1(net412),
    .X(_00085_));
 sky130_fd_sc_hd__o221a_1 _13422_ (.A1(net411),
    .A2(net249),
    .B1(net183),
    .B2(net357),
    .C1(net279),
    .X(_06349_));
 sky130_fd_sc_hd__o21a_1 _13423_ (.A1(_00404_),
    .A2(net161),
    .B1(net437),
    .X(_00086_));
 sky130_fd_sc_hd__o221a_1 _13424_ (.A1(net357),
    .A2(net249),
    .B1(net183),
    .B2(\div_shifter[21] ),
    .C1(net279),
    .X(_06350_));
 sky130_fd_sc_hd__o21a_1 _13425_ (.A1(net97),
    .A2(net161),
    .B1(net358),
    .X(_00087_));
 sky130_fd_sc_hd__o221a_1 _13426_ (.A1(\div_shifter[21] ),
    .A2(net249),
    .B1(net183),
    .B2(net444),
    .C1(net279),
    .X(_06352_));
 sky130_fd_sc_hd__o21a_1 _13427_ (.A1(_00278_),
    .A2(net161),
    .B1(net445),
    .X(_00088_));
 sky130_fd_sc_hd__o221a_1 _13428_ (.A1(\div_shifter[22] ),
    .A2(_04412_),
    .B1(net183),
    .B2(net368),
    .C1(net279),
    .X(_06353_));
 sky130_fd_sc_hd__o21a_1 _13429_ (.A1(net98),
    .A2(net162),
    .B1(net369),
    .X(_00089_));
 sky130_fd_sc_hd__o221a_1 _13430_ (.A1(net368),
    .A2(_04412_),
    .B1(net183),
    .B2(net428),
    .C1(net279),
    .X(_06354_));
 sky130_fd_sc_hd__o21a_1 _13431_ (.A1(_00331_),
    .A2(net162),
    .B1(net429),
    .X(_00090_));
 sky130_fd_sc_hd__o221a_1 _13432_ (.A1(\div_shifter[24] ),
    .A2(net249),
    .B1(net183),
    .B2(net393),
    .C1(net281),
    .X(_06355_));
 sky130_fd_sc_hd__o21a_1 _13433_ (.A1(net92),
    .A2(net162),
    .B1(net394),
    .X(_00091_));
 sky130_fd_sc_hd__o221a_1 _13434_ (.A1(net393),
    .A2(net249),
    .B1(net183),
    .B2(net351),
    .C1(net281),
    .X(_06356_));
 sky130_fd_sc_hd__o21a_1 _13435_ (.A1(_00313_),
    .A2(net162),
    .B1(net408),
    .X(_00092_));
 sky130_fd_sc_hd__o221a_1 _13436_ (.A1(net351),
    .A2(net249),
    .B1(net183),
    .B2(net323),
    .C1(net281),
    .X(_06358_));
 sky130_fd_sc_hd__o21a_1 _13437_ (.A1(net93),
    .A2(net162),
    .B1(net352),
    .X(_00093_));
 sky130_fd_sc_hd__o221a_1 _13438_ (.A1(net323),
    .A2(net249),
    .B1(net183),
    .B2(\div_shifter[28] ),
    .C1(net281),
    .X(_06359_));
 sky130_fd_sc_hd__o21a_1 _13439_ (.A1(_00558_),
    .A2(net162),
    .B1(net324),
    .X(_00094_));
 sky130_fd_sc_hd__o221a_1 _13440_ (.A1(net379),
    .A2(net249),
    .B1(net183),
    .B2(net330),
    .C1(net281),
    .X(_06360_));
 sky130_fd_sc_hd__o21a_1 _13441_ (.A1(_00787_),
    .A2(net162),
    .B1(net380),
    .X(_00095_));
 sky130_fd_sc_hd__o221a_1 _13442_ (.A1(net330),
    .A2(net249),
    .B1(net183),
    .B2(\div_shifter[30] ),
    .C1(net282),
    .X(_06361_));
 sky130_fd_sc_hd__o21a_1 _13443_ (.A1(_02078_),
    .A2(net161),
    .B1(net331),
    .X(_00096_));
 sky130_fd_sc_hd__o221a_1 _13444_ (.A1(net421),
    .A2(net249),
    .B1(net183),
    .B2(\div_shifter[31] ),
    .C1(net282),
    .X(_06362_));
 sky130_fd_sc_hd__o21a_1 _13445_ (.A1(net61),
    .A2(net161),
    .B1(net422),
    .X(_00097_));
 sky130_fd_sc_hd__nand3_1 _13446_ (.A(\div_shifter[31] ),
    .B(net311),
    .C(net2),
    .Y(_06364_));
 sky130_fd_sc_hd__a21o_1 _13447_ (.A1(net311),
    .A2(net2),
    .B1(\div_shifter[31] ),
    .X(_06365_));
 sky130_fd_sc_hd__a32o_1 _13448_ (.A1(net251),
    .A2(_06364_),
    .A3(_06365_),
    .B1(net185),
    .B2(net543),
    .X(_06366_));
 sky130_fd_sc_hd__and2_1 _13449_ (.A(net276),
    .B(net544),
    .X(_00098_));
 sky130_fd_sc_hd__and2_1 _13450_ (.A(net560),
    .B(net185),
    .X(_06367_));
 sky130_fd_sc_hd__xnor2_1 _13451_ (.A(_06247_),
    .B(_06248_),
    .Y(_06368_));
 sky130_fd_sc_hd__nand2_1 _13452_ (.A(net2),
    .B(_06368_),
    .Y(_06369_));
 sky130_fd_sc_hd__o211a_1 _13453_ (.A1(net543),
    .A2(net2),
    .B1(_06369_),
    .C1(net251),
    .X(_06370_));
 sky130_fd_sc_hd__o21a_1 _13454_ (.A1(_06367_),
    .A2(_06370_),
    .B1(net273),
    .X(_00099_));
 sky130_fd_sc_hd__nand2b_1 _13455_ (.A_N(_06244_),
    .B(_06245_),
    .Y(_06371_));
 sky130_fd_sc_hd__xnor2_1 _13456_ (.A(_06249_),
    .B(_06371_),
    .Y(_06373_));
 sky130_fd_sc_hd__mux2_1 _13457_ (.A0(net560),
    .A1(_06373_),
    .S(net1),
    .X(_06374_));
 sky130_fd_sc_hd__a22o_1 _13458_ (.A1(net583),
    .A2(net185),
    .B1(_06374_),
    .B2(net251),
    .X(_06375_));
 sky130_fd_sc_hd__and2_1 _13459_ (.A(net273),
    .B(net584),
    .X(_00100_));
 sky130_fd_sc_hd__nand2b_1 _13460_ (.A_N(_06242_),
    .B(_06243_),
    .Y(_06376_));
 sky130_fd_sc_hd__xnor2_1 _13461_ (.A(_06250_),
    .B(_06376_),
    .Y(_06377_));
 sky130_fd_sc_hd__mux2_1 _13462_ (.A0(\div_shifter[34] ),
    .A1(_06377_),
    .S(net1),
    .X(_06378_));
 sky130_fd_sc_hd__a22o_1 _13463_ (.A1(net562),
    .A2(net185),
    .B1(_06378_),
    .B2(net251),
    .X(_06379_));
 sky130_fd_sc_hd__and2_1 _13464_ (.A(net276),
    .B(net563),
    .X(_00101_));
 sky130_fd_sc_hd__xnor2_1 _13465_ (.A(_06241_),
    .B(_06252_),
    .Y(_06380_));
 sky130_fd_sc_hd__mux2_1 _13466_ (.A0(net562),
    .A1(_06380_),
    .S(net1),
    .X(_06382_));
 sky130_fd_sc_hd__a22o_1 _13467_ (.A1(net581),
    .A2(net186),
    .B1(_06382_),
    .B2(net252),
    .X(_06383_));
 sky130_fd_sc_hd__and2_1 _13468_ (.A(net276),
    .B(net582),
    .X(_00102_));
 sky130_fd_sc_hd__xnor2_1 _13469_ (.A(_06237_),
    .B(_06253_),
    .Y(_06384_));
 sky130_fd_sc_hd__mux2_1 _13470_ (.A0(net581),
    .A1(_06384_),
    .S(net2),
    .X(_06385_));
 sky130_fd_sc_hd__a22o_1 _13471_ (.A1(net592),
    .A2(net187),
    .B1(_06385_),
    .B2(net253),
    .X(_06386_));
 sky130_fd_sc_hd__and2_1 _13472_ (.A(net276),
    .B(_06386_),
    .X(_00103_));
 sky130_fd_sc_hd__nand2b_1 _13473_ (.A_N(_06233_),
    .B(_06234_),
    .Y(_06387_));
 sky130_fd_sc_hd__xnor2_1 _13474_ (.A(_06254_),
    .B(_06387_),
    .Y(_06388_));
 sky130_fd_sc_hd__mux2_1 _13475_ (.A0(\div_shifter[37] ),
    .A1(_06388_),
    .S(net2),
    .X(_06389_));
 sky130_fd_sc_hd__a22o_1 _13476_ (.A1(net585),
    .A2(net187),
    .B1(_06389_),
    .B2(net253),
    .X(_06391_));
 sky130_fd_sc_hd__and2_1 _13477_ (.A(net277),
    .B(net586),
    .X(_00104_));
 sky130_fd_sc_hd__nand2b_1 _13478_ (.A_N(_06231_),
    .B(_06232_),
    .Y(_06392_));
 sky130_fd_sc_hd__xnor2_1 _13479_ (.A(_06255_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__mux2_1 _13480_ (.A0(\div_shifter[38] ),
    .A1(_06393_),
    .S(net2),
    .X(_06394_));
 sky130_fd_sc_hd__a22o_1 _13481_ (.A1(net574),
    .A2(net187),
    .B1(_06394_),
    .B2(net253),
    .X(_06395_));
 sky130_fd_sc_hd__and2_1 _13482_ (.A(net277),
    .B(net575),
    .X(_00105_));
 sky130_fd_sc_hd__nand2b_1 _13483_ (.A_N(_06228_),
    .B(_06230_),
    .Y(_06396_));
 sky130_fd_sc_hd__xnor2_1 _13484_ (.A(_06256_),
    .B(_06396_),
    .Y(_06397_));
 sky130_fd_sc_hd__mux2_1 _13485_ (.A0(net574),
    .A1(_06397_),
    .S(net532),
    .X(_06398_));
 sky130_fd_sc_hd__a22o_1 _13486_ (.A1(net593),
    .A2(net186),
    .B1(_06398_),
    .B2(net252),
    .X(_06400_));
 sky130_fd_sc_hd__and2_1 _13487_ (.A(net275),
    .B(_06400_),
    .X(_00106_));
 sky130_fd_sc_hd__nand2b_1 _13488_ (.A_N(_06226_),
    .B(_06227_),
    .Y(_06401_));
 sky130_fd_sc_hd__xnor2_1 _13489_ (.A(_06257_),
    .B(_06401_),
    .Y(_06402_));
 sky130_fd_sc_hd__mux2_1 _13490_ (.A0(\div_shifter[40] ),
    .A1(_06402_),
    .S(net1),
    .X(_06403_));
 sky130_fd_sc_hd__a22o_1 _13491_ (.A1(net551),
    .A2(net186),
    .B1(_06403_),
    .B2(net252),
    .X(_06404_));
 sky130_fd_sc_hd__and2_1 _13492_ (.A(net274),
    .B(net552),
    .X(_00107_));
 sky130_fd_sc_hd__nand2b_1 _13493_ (.A_N(_06224_),
    .B(_06225_),
    .Y(_06405_));
 sky130_fd_sc_hd__xnor2_1 _13494_ (.A(_06258_),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__mux2_1 _13495_ (.A0(net551),
    .A1(_06406_),
    .S(net532),
    .X(_06407_));
 sky130_fd_sc_hd__a22o_1 _13496_ (.A1(net578),
    .A2(net186),
    .B1(_06407_),
    .B2(net252),
    .X(_06409_));
 sky130_fd_sc_hd__and2_1 _13497_ (.A(net274),
    .B(net579),
    .X(_00108_));
 sky130_fd_sc_hd__nand2b_1 _13498_ (.A_N(_06222_),
    .B(_06223_),
    .Y(_06410_));
 sky130_fd_sc_hd__xnor2_1 _13499_ (.A(_06259_),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__mux2_1 _13500_ (.A0(net578),
    .A1(_06411_),
    .S(net1),
    .X(_06412_));
 sky130_fd_sc_hd__a22o_1 _13501_ (.A1(net589),
    .A2(net184),
    .B1(_06412_),
    .B2(net250),
    .X(_06413_));
 sky130_fd_sc_hd__and2_1 _13502_ (.A(net274),
    .B(_06413_),
    .X(_00109_));
 sky130_fd_sc_hd__nand2b_1 _13503_ (.A_N(_06220_),
    .B(_06221_),
    .Y(_06414_));
 sky130_fd_sc_hd__xnor2_1 _13504_ (.A(_06260_),
    .B(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__mux2_1 _13505_ (.A0(\div_shifter[43] ),
    .A1(_06415_),
    .S(net1),
    .X(_06416_));
 sky130_fd_sc_hd__a22o_1 _13506_ (.A1(net569),
    .A2(net184),
    .B1(_06416_),
    .B2(net250),
    .X(_06418_));
 sky130_fd_sc_hd__and2_1 _13507_ (.A(net274),
    .B(net570),
    .X(_00110_));
 sky130_fd_sc_hd__nand2b_1 _13508_ (.A_N(_06217_),
    .B(_06219_),
    .Y(_06419_));
 sky130_fd_sc_hd__xnor2_1 _13509_ (.A(_06261_),
    .B(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__mux2_1 _13510_ (.A0(net569),
    .A1(_06420_),
    .S(net1),
    .X(_06421_));
 sky130_fd_sc_hd__a22o_1 _13511_ (.A1(net587),
    .A2(net186),
    .B1(_06421_),
    .B2(net252),
    .X(_06422_));
 sky130_fd_sc_hd__and2_1 _13512_ (.A(net274),
    .B(net588),
    .X(_00111_));
 sky130_fd_sc_hd__nand2b_1 _13513_ (.A_N(_06215_),
    .B(_06216_),
    .Y(_06423_));
 sky130_fd_sc_hd__xnor2_1 _13514_ (.A(_06263_),
    .B(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__mux2_1 _13515_ (.A0(\div_shifter[45] ),
    .A1(_06424_),
    .S(net1),
    .X(_06425_));
 sky130_fd_sc_hd__a22o_1 _13516_ (.A1(net549),
    .A2(net186),
    .B1(_06425_),
    .B2(net252),
    .X(_06427_));
 sky130_fd_sc_hd__and2_1 _13517_ (.A(net274),
    .B(net550),
    .X(_00112_));
 sky130_fd_sc_hd__nand2b_1 _13518_ (.A_N(_06213_),
    .B(_06214_),
    .Y(_06428_));
 sky130_fd_sc_hd__xnor2_1 _13519_ (.A(_06264_),
    .B(_06428_),
    .Y(_06429_));
 sky130_fd_sc_hd__mux2_1 _13520_ (.A0(net549),
    .A1(_06429_),
    .S(net1),
    .X(_06430_));
 sky130_fd_sc_hd__a22o_1 _13521_ (.A1(net594),
    .A2(net186),
    .B1(_06430_),
    .B2(net252),
    .X(_06431_));
 sky130_fd_sc_hd__and2_1 _13522_ (.A(net275),
    .B(_06431_),
    .X(_00113_));
 sky130_fd_sc_hd__xnor2_1 _13523_ (.A(_06212_),
    .B(_06265_),
    .Y(_06432_));
 sky130_fd_sc_hd__mux2_1 _13524_ (.A0(\div_shifter[47] ),
    .A1(_06432_),
    .S(net1),
    .X(_06433_));
 sky130_fd_sc_hd__a22o_1 _13525_ (.A1(net590),
    .A2(net186),
    .B1(_06433_),
    .B2(net252),
    .X(_06434_));
 sky130_fd_sc_hd__and2_1 _13526_ (.A(net275),
    .B(net591),
    .X(_00114_));
 sky130_fd_sc_hd__xor2_1 _13527_ (.A(_06209_),
    .B(_06266_),
    .X(_06436_));
 sky130_fd_sc_hd__mux2_1 _13528_ (.A0(\div_shifter[48] ),
    .A1(_06436_),
    .S(net1),
    .X(_06437_));
 sky130_fd_sc_hd__a22o_1 _13529_ (.A1(net555),
    .A2(net186),
    .B1(_06437_),
    .B2(net252),
    .X(_06438_));
 sky130_fd_sc_hd__and2_1 _13530_ (.A(net275),
    .B(net556),
    .X(_00115_));
 sky130_fd_sc_hd__xnor2_1 _13531_ (.A(_06205_),
    .B(_06267_),
    .Y(_06439_));
 sky130_fd_sc_hd__mux2_1 _13532_ (.A0(net555),
    .A1(_06439_),
    .S(net1),
    .X(_06440_));
 sky130_fd_sc_hd__a22o_1 _13533_ (.A1(net557),
    .A2(net186),
    .B1(_06440_),
    .B2(net252),
    .X(_06441_));
 sky130_fd_sc_hd__and2_1 _13534_ (.A(net275),
    .B(net558),
    .X(_00116_));
 sky130_fd_sc_hd__nand2b_1 _13535_ (.A_N(_06201_),
    .B(_06202_),
    .Y(_06442_));
 sky130_fd_sc_hd__xnor2_1 _13536_ (.A(_06268_),
    .B(_06442_),
    .Y(_06444_));
 sky130_fd_sc_hd__mux2_1 _13537_ (.A0(net557),
    .A1(_06444_),
    .S(net1),
    .X(_06445_));
 sky130_fd_sc_hd__a22o_1 _13538_ (.A1(net559),
    .A2(net186),
    .B1(_06445_),
    .B2(net252),
    .X(_06446_));
 sky130_fd_sc_hd__and2_1 _13539_ (.A(net275),
    .B(_06446_),
    .X(_00117_));
 sky130_fd_sc_hd__xnor2_1 _13540_ (.A(_06200_),
    .B(_06269_),
    .Y(_06447_));
 sky130_fd_sc_hd__mux2_1 _13541_ (.A0(net559),
    .A1(_06447_),
    .S(net1),
    .X(_06448_));
 sky130_fd_sc_hd__a22o_1 _13542_ (.A1(net573),
    .A2(net186),
    .B1(_06448_),
    .B2(net252),
    .X(_06449_));
 sky130_fd_sc_hd__and2_1 _13543_ (.A(net274),
    .B(_06449_),
    .X(_00118_));
 sky130_fd_sc_hd__xor2_1 _13544_ (.A(_06197_),
    .B(_06270_),
    .X(_06450_));
 sky130_fd_sc_hd__mux2_1 _13545_ (.A0(\div_shifter[52] ),
    .A1(_06450_),
    .S(net1),
    .X(_06451_));
 sky130_fd_sc_hd__a22o_1 _13546_ (.A1(net564),
    .A2(net186),
    .B1(_06451_),
    .B2(net253),
    .X(_06453_));
 sky130_fd_sc_hd__and2_1 _13547_ (.A(net276),
    .B(net565),
    .X(_00119_));
 sky130_fd_sc_hd__xnor2_1 _13548_ (.A(_06193_),
    .B(_06271_),
    .Y(_06454_));
 sky130_fd_sc_hd__mux2_1 _13549_ (.A0(\div_shifter[53] ),
    .A1(_06454_),
    .S(net532),
    .X(_06455_));
 sky130_fd_sc_hd__a22o_1 _13550_ (.A1(net553),
    .A2(net187),
    .B1(_06455_),
    .B2(net253),
    .X(_06456_));
 sky130_fd_sc_hd__and2_1 _13551_ (.A(net277),
    .B(net554),
    .X(_00120_));
 sky130_fd_sc_hd__nand2b_1 _13552_ (.A_N(_06189_),
    .B(_06190_),
    .Y(_06457_));
 sky130_fd_sc_hd__xnor2_1 _13553_ (.A(_06272_),
    .B(_06457_),
    .Y(_06458_));
 sky130_fd_sc_hd__mux2_1 _13554_ (.A0(net553),
    .A1(_06458_),
    .S(net2),
    .X(_06459_));
 sky130_fd_sc_hd__a22o_1 _13555_ (.A1(net580),
    .A2(net186),
    .B1(_06459_),
    .B2(net253),
    .X(_06460_));
 sky130_fd_sc_hd__and2_1 _13556_ (.A(net277),
    .B(_06460_),
    .X(_00121_));
 sky130_fd_sc_hd__xnor2_1 _13557_ (.A(_06188_),
    .B(_06274_),
    .Y(_06462_));
 sky130_fd_sc_hd__mux2_1 _13558_ (.A0(\div_shifter[55] ),
    .A1(_06462_),
    .S(net2),
    .X(_06463_));
 sky130_fd_sc_hd__a22o_1 _13559_ (.A1(net567),
    .A2(net188),
    .B1(_06463_),
    .B2(net253),
    .X(_06464_));
 sky130_fd_sc_hd__and2_1 _13560_ (.A(net277),
    .B(net568),
    .X(_00122_));
 sky130_fd_sc_hd__xor2_1 _13561_ (.A(_06184_),
    .B(_06275_),
    .X(_06465_));
 sky130_fd_sc_hd__mux2_1 _13562_ (.A0(net567),
    .A1(_06465_),
    .S(net2),
    .X(_06466_));
 sky130_fd_sc_hd__a22o_1 _13563_ (.A1(net576),
    .A2(net188),
    .B1(_06466_),
    .B2(net253),
    .X(_06467_));
 sky130_fd_sc_hd__and2_1 _13564_ (.A(net277),
    .B(net577),
    .X(_00123_));
 sky130_fd_sc_hd__xnor2_1 _13565_ (.A(_06181_),
    .B(_06276_),
    .Y(_06468_));
 sky130_fd_sc_hd__mux2_1 _13566_ (.A0(\div_shifter[57] ),
    .A1(_06468_),
    .S(net2),
    .X(_06470_));
 sky130_fd_sc_hd__a22o_1 _13567_ (.A1(net571),
    .A2(net188),
    .B1(_06470_),
    .B2(net254),
    .X(_06471_));
 sky130_fd_sc_hd__and2_1 _13568_ (.A(net281),
    .B(net572),
    .X(_00124_));
 sky130_fd_sc_hd__nand2b_1 _13569_ (.A_N(_06177_),
    .B(_06178_),
    .Y(_06472_));
 sky130_fd_sc_hd__xnor2_1 _13570_ (.A(_06277_),
    .B(_06472_),
    .Y(_06473_));
 sky130_fd_sc_hd__mux2_1 _13571_ (.A0(\div_shifter[58] ),
    .A1(_06473_),
    .S(net2),
    .X(_06474_));
 sky130_fd_sc_hd__a22o_1 _13572_ (.A1(net547),
    .A2(net188),
    .B1(_06474_),
    .B2(net254),
    .X(_06475_));
 sky130_fd_sc_hd__and2_1 _13573_ (.A(net280),
    .B(net548),
    .X(_00125_));
 sky130_fd_sc_hd__and2b_1 _13574_ (.A_N(_06176_),
    .B(_06278_),
    .X(_06476_));
 sky130_fd_sc_hd__nor2_1 _13575_ (.A(_06279_),
    .B(_06476_),
    .Y(_06477_));
 sky130_fd_sc_hd__mux2_1 _13576_ (.A0(\div_shifter[59] ),
    .A1(_06477_),
    .S(net2),
    .X(_06479_));
 sky130_fd_sc_hd__a22o_1 _13577_ (.A1(net545),
    .A2(net188),
    .B1(_06479_),
    .B2(net254),
    .X(_06480_));
 sky130_fd_sc_hd__and2_1 _13578_ (.A(net280),
    .B(net546),
    .X(_00126_));
 sky130_fd_sc_hd__nor3_1 _13579_ (.A(_06172_),
    .B(_06173_),
    .C(_06279_),
    .Y(_06481_));
 sky130_fd_sc_hd__nor2_1 _13580_ (.A(_06280_),
    .B(_06481_),
    .Y(_06482_));
 sky130_fd_sc_hd__mux2_1 _13581_ (.A0(net545),
    .A1(_06482_),
    .S(net2),
    .X(_06483_));
 sky130_fd_sc_hd__a22o_1 _13582_ (.A1(net566),
    .A2(net188),
    .B1(_06483_),
    .B2(net254),
    .X(_06484_));
 sky130_fd_sc_hd__and2_1 _13583_ (.A(net280),
    .B(_06484_),
    .X(_00127_));
 sky130_fd_sc_hd__and2_1 _13584_ (.A(net531),
    .B(net188),
    .X(_06485_));
 sky130_fd_sc_hd__xnor2_1 _13585_ (.A(_06169_),
    .B(_06281_),
    .Y(_06486_));
 sky130_fd_sc_hd__nand2_1 _13586_ (.A(net2),
    .B(_06486_),
    .Y(_06488_));
 sky130_fd_sc_hd__o211a_1 _13587_ (.A1(net566),
    .A2(net2),
    .B1(_06488_),
    .C1(net254),
    .X(_06489_));
 sky130_fd_sc_hd__o21a_1 _13588_ (.A1(_06485_),
    .A2(_06489_),
    .B1(net281),
    .X(_00128_));
 sky130_fd_sc_hd__xor2_1 _13589_ (.A(\divi2_l[31] ),
    .B(_06282_),
    .X(_06490_));
 sky130_fd_sc_hd__a32o_1 _13590_ (.A1(\div_shifter[62] ),
    .A2(net254),
    .A3(_06490_),
    .B1(net188),
    .B2(net438),
    .X(_06491_));
 sky130_fd_sc_hd__and2_1 _13591_ (.A(net277),
    .B(net439),
    .X(_00129_));
 sky130_fd_sc_hd__a21o_1 _13592_ (.A1(net489),
    .A2(net254),
    .B1(net166),
    .X(_06492_));
 sky130_fd_sc_hd__or2_1 _13593_ (.A(net489),
    .B(net254),
    .X(_06493_));
 sky130_fd_sc_hd__and3b_1 _13594_ (.A_N(_06492_),
    .B(_06493_),
    .C(net280),
    .X(_00130_));
 sky130_fd_sc_hd__a21oi_1 _13595_ (.A1(net489),
    .A2(net254),
    .B1(net301),
    .Y(_06494_));
 sky130_fd_sc_hd__a211oi_1 _13596_ (.A1(net301),
    .A2(_06492_),
    .B1(_06494_),
    .C1(rst),
    .Y(_00131_));
 sky130_fd_sc_hd__and2_1 _13597_ (.A(net254),
    .B(_06122_),
    .X(_06496_));
 sky130_fd_sc_hd__and3b_1 _13598_ (.A_N(_06496_),
    .B(net467),
    .C(net162),
    .X(_06497_));
 sky130_fd_sc_hd__and4b_1 _13599_ (.A_N(net467),
    .B(net301),
    .C(net516),
    .D(net254),
    .X(_06498_));
 sky130_fd_sc_hd__o21a_1 _13600_ (.A1(net468),
    .A2(_06498_),
    .B1(net280),
    .X(_00132_));
 sky130_fd_sc_hd__o21ai_1 _13601_ (.A1(net166),
    .A2(_06496_),
    .B1(net313),
    .Y(_06499_));
 sky130_fd_sc_hd__o211a_1 _13602_ (.A1(net313),
    .A2(_06496_),
    .B1(_06499_),
    .C1(net280),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_1 _13603_ (.A1(net441),
    .A2(net188),
    .B1(_06123_),
    .B2(net254),
    .X(_06500_));
 sky130_fd_sc_hd__a21o_1 _13604_ (.A1(net313),
    .A2(_06122_),
    .B1(net441),
    .X(_06501_));
 sky130_fd_sc_hd__and3_1 _13605_ (.A(net280),
    .B(_06500_),
    .C(net442),
    .X(_00134_));
 sky130_fd_sc_hd__o21a_1 _13606_ (.A1(net457),
    .A2(_06124_),
    .B1(net281),
    .X(_00135_));
 sky130_fd_sc_hd__dfxtp_1 _13607_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00000_),
    .Q(busy_l));
 sky130_fd_sc_hd__dfxtp_1 _13608_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00001_),
    .Q(divi1_sign));
 sky130_fd_sc_hd__dfxtp_1 _13609_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net312),
    .Q(\divi2_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13610_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net310),
    .Q(\divi2_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13611_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net308),
    .Q(\divi2_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13612_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net306),
    .Q(\divi2_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13613_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00006_),
    .Q(\divi2_l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13614_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net378),
    .Q(\divi2_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13615_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00008_),
    .Q(\divi2_l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13616_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net373),
    .Q(\divi2_l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13617_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00010_),
    .Q(\divi2_l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13618_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00011_),
    .Q(\divi2_l[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13619_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00012_),
    .Q(\divi2_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13620_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00013_),
    .Q(\divi2_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13621_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00014_),
    .Q(\divi2_l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13622_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00015_),
    .Q(\divi2_l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13623_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00016_),
    .Q(\divi2_l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13624_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00017_),
    .Q(\divi2_l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13625_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00018_),
    .Q(\divi2_l[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13626_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00019_),
    .Q(\divi2_l[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13627_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00020_),
    .Q(\divi2_l[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13628_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00021_),
    .Q(\divi2_l[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13629_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00022_),
    .Q(\divi2_l[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13630_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net385),
    .Q(\divi2_l[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13631_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net348),
    .Q(\divi2_l[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13632_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00025_),
    .Q(\divi2_l[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13633_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00026_),
    .Q(\divi2_l[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13634_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net339),
    .Q(\divi2_l[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13635_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00028_),
    .Q(\divi2_l[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13636_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00029_),
    .Q(\divi2_l[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13637_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00030_),
    .Q(\divi2_l[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13638_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00031_),
    .Q(\divi2_l[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13639_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00032_),
    .Q(\divi2_l[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13640_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00033_),
    .Q(\divi2_l[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13641_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00034_),
    .Q(\div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13642_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net488),
    .Q(\div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13643_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00036_),
    .Q(\div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13644_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net526),
    .Q(\div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13645_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00038_),
    .Q(\div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13646_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net482),
    .Q(\div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13647_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00040_),
    .Q(\div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13648_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00041_),
    .Q(\div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13649_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00042_),
    .Q(\div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13650_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net463),
    .Q(\div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13651_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net540),
    .Q(\div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13652_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net509),
    .Q(\div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13653_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00046_),
    .Q(\div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13654_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00047_),
    .Q(\div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13655_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00048_),
    .Q(\div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13656_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00049_),
    .Q(\div_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13657_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00050_),
    .Q(\div_res[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13658_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net500),
    .Q(\div_res[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13659_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00052_),
    .Q(\div_res[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13660_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net485),
    .Q(\div_res[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13661_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net477),
    .Q(\div_res[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13662_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00055_),
    .Q(\div_res[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13663_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net474),
    .Q(\div_res[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13664_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00057_),
    .Q(\div_res[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13665_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00058_),
    .Q(\div_res[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13666_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00059_),
    .Q(\div_res[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13667_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00060_),
    .Q(\div_res[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13668_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net466),
    .Q(\div_res[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13669_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net519),
    .Q(\div_res[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13670_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net497),
    .Q(\div_res[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13671_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00064_),
    .Q(\div_res[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13672_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net454),
    .Q(\div_res[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13673_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00066_),
    .Q(\div_shifter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13674_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net300),
    .Q(\div_shifter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13675_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00068_),
    .Q(\div_shifter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13676_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00069_),
    .Q(\div_shifter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13677_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00070_),
    .Q(\div_shifter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13678_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net398),
    .Q(\div_shifter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13679_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00072_),
    .Q(\div_shifter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13680_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net304),
    .Q(\div_shifter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13681_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00074_),
    .Q(\div_shifter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13682_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00075_),
    .Q(\div_shifter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13683_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net319),
    .Q(\div_shifter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13684_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00077_),
    .Q(\div_shifter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13685_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net420),
    .Q(\div_shifter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13686_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net392),
    .Q(\div_shifter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13687_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00080_),
    .Q(\div_shifter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13688_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00081_),
    .Q(\div_shifter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13689_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00082_),
    .Q(\div_shifter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13690_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net322),
    .Q(\div_shifter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13691_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net451),
    .Q(\div_shifter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13692_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net413),
    .Q(\div_shifter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13693_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00086_),
    .Q(\div_shifter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13694_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net359),
    .Q(\div_shifter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13695_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net446),
    .Q(\div_shifter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13696_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net370),
    .Q(\div_shifter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13697_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00090_),
    .Q(\div_shifter[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13698_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net395),
    .Q(\div_shifter[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13699_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00092_),
    .Q(\div_shifter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13700_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00093_),
    .Q(\div_shifter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13701_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net325),
    .Q(\div_shifter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13702_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00095_),
    .Q(\div_shifter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13703_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net332),
    .Q(\div_shifter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13704_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net423),
    .Q(\div_shifter[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13705_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00098_),
    .Q(\div_shifter[32] ));
 sky130_fd_sc_hd__dfxtp_2 _13706_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net561),
    .Q(\div_shifter[33] ));
 sky130_fd_sc_hd__dfxtp_2 _13707_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00100_),
    .Q(\div_shifter[34] ));
 sky130_fd_sc_hd__dfxtp_1 _13708_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00101_),
    .Q(\div_shifter[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13709_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00102_),
    .Q(\div_shifter[36] ));
 sky130_fd_sc_hd__dfxtp_2 _13710_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00103_),
    .Q(\div_shifter[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13711_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00104_),
    .Q(\div_shifter[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13712_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00105_),
    .Q(\div_shifter[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13713_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00106_),
    .Q(\div_shifter[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13714_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00107_),
    .Q(\div_shifter[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13715_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00108_),
    .Q(\div_shifter[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13716_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00109_),
    .Q(\div_shifter[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13717_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00110_),
    .Q(\div_shifter[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13718_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00111_),
    .Q(\div_shifter[45] ));
 sky130_fd_sc_hd__dfxtp_1 _13719_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00112_),
    .Q(\div_shifter[46] ));
 sky130_fd_sc_hd__dfxtp_2 _13720_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00113_),
    .Q(\div_shifter[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13721_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00114_),
    .Q(\div_shifter[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13722_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00115_),
    .Q(\div_shifter[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13723_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00116_),
    .Q(\div_shifter[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13724_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00117_),
    .Q(\div_shifter[51] ));
 sky130_fd_sc_hd__dfxtp_1 _13725_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00118_),
    .Q(\div_shifter[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13726_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00119_),
    .Q(\div_shifter[53] ));
 sky130_fd_sc_hd__dfxtp_1 _13727_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00120_),
    .Q(\div_shifter[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13728_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00121_),
    .Q(\div_shifter[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13729_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00122_),
    .Q(\div_shifter[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13730_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00123_),
    .Q(\div_shifter[57] ));
 sky130_fd_sc_hd__dfxtp_1 _13731_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00124_),
    .Q(\div_shifter[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13732_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00125_),
    .Q(\div_shifter[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13733_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00126_),
    .Q(\div_shifter[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13734_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00127_),
    .Q(\div_shifter[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13735_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00128_),
    .Q(\div_shifter[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13736_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net440),
    .Q(\div_shifter[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13737_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00130_),
    .Q(\div_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13738_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net302),
    .Q(\div_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13739_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net469),
    .Q(\div_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13740_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net314),
    .Q(\div_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13741_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net443),
    .Q(\div_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13742_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net458),
    .Q(div_complete));
 sky130_fd_sc_hd__buf_12 _13743_ (.A(instruction[5]),
    .X(loadstore_size[0]));
 sky130_fd_sc_hd__buf_12 _13744_ (.A(net297),
    .X(loadstore_size[1]));
 sky130_fd_sc_hd__buf_12 _13745_ (.A(instruction[8]),
    .X(pred_idx[0]));
 sky130_fd_sc_hd__buf_12 _13746_ (.A(instruction[9]),
    .X(pred_idx[1]));
 sky130_fd_sc_hd__buf_12 _13747_ (.A(instruction[10]),
    .X(pred_idx[2]));
 sky130_fd_sc_hd__buf_12 _13748_ (.A(net298),
    .X(sign_extend));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__buf_6 fanout1 (.A(_06286_),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_8 fanout10 (.A(_02066_),
    .X(net10));
 sky130_fd_sc_hd__buf_8 fanout100 (.A(_00230_),
    .X(net100));
 sky130_fd_sc_hd__buf_8 fanout103 (.A(_00219_),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_8 fanout104 (.A(_00196_),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(_00196_),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(_00477_),
    .X(net106));
 sky130_fd_sc_hd__buf_12 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__buf_8 fanout109 (.A(_00430_),
    .X(net109));
 sky130_fd_sc_hd__buf_6 fanout110 (.A(_00415_),
    .X(net110));
 sky130_fd_sc_hd__buf_6 fanout111 (.A(_00414_),
    .X(net111));
 sky130_fd_sc_hd__buf_8 fanout113 (.A(_00411_),
    .X(net113));
 sky130_fd_sc_hd__buf_8 fanout115 (.A(_00391_),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_16 fanout116 (.A(net118),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_16 fanout117 (.A(net118),
    .X(net117));
 sky130_fd_sc_hd__buf_8 fanout118 (.A(_00380_),
    .X(net118));
 sky130_fd_sc_hd__buf_6 fanout119 (.A(_00376_),
    .X(net119));
 sky130_fd_sc_hd__buf_6 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(_00376_),
    .X(net120));
 sky130_fd_sc_hd__buf_6 fanout123 (.A(_00371_),
    .X(net123));
 sky130_fd_sc_hd__buf_6 fanout124 (.A(_00286_),
    .X(net124));
 sky130_fd_sc_hd__buf_6 fanout125 (.A(_00267_),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(_00231_),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(_00231_),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_8 fanout128 (.A(_00228_),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(_00228_),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_8 fanout13 (.A(_00798_),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(_00205_),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_8 fanout131 (.A(_00205_),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_8 fanout132 (.A(_00157_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_8 fanout133 (.A(_06701_),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(_06681_),
    .X(net135));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(net144),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__buf_4 fanout138 (.A(net144),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net141),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_8 fanout14 (.A(_00337_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 fanout141 (.A(net144),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 fanout144 (.A(_06680_),
    .X(net144));
 sky130_fd_sc_hd__buf_8 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_12 fanout146 (.A(net147),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_16 fanout147 (.A(_00452_),
    .X(net147));
 sky130_fd_sc_hd__buf_6 fanout149 (.A(_00339_),
    .X(net149));
 sky130_fd_sc_hd__buf_4 fanout15 (.A(_00337_),
    .X(net15));
 sky130_fd_sc_hd__buf_6 fanout150 (.A(_00327_),
    .X(net150));
 sky130_fd_sc_hd__buf_8 fanout151 (.A(_00326_),
    .X(net151));
 sky130_fd_sc_hd__buf_6 fanout152 (.A(_00320_),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_16 fanout154 (.A(net156),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_8 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_12 fanout156 (.A(_00215_),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_8 fanout157 (.A(_00160_),
    .X(net157));
 sky130_fd_sc_hd__buf_6 fanout158 (.A(_06727_),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_8 fanout159 (.A(net163),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_8 fanout16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__buf_4 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 fanout163 (.A(_06126_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_4 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(_06125_),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(_02424_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_8 fanout168 (.A(_02355_),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_4 fanout169 (.A(_02355_),
    .X(net169));
 sky130_fd_sc_hd__buf_8 fanout17 (.A(_00562_),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(net172),
    .X(net170));
 sky130_fd_sc_hd__buf_4 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(_02354_),
    .X(net172));
 sky130_fd_sc_hd__buf_12 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_16 fanout175 (.A(_00187_),
    .X(net175));
 sky130_fd_sc_hd__buf_6 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__buf_8 fanout178 (.A(_06704_),
    .X(net178));
 sky130_fd_sc_hd__buf_12 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout18 (.A(_00413_),
    .X(net18));
 sky130_fd_sc_hd__buf_8 fanout180 (.A(_06690_),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_16 fanout181 (.A(_06689_),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__buf_4 fanout183 (.A(_06662_),
    .X(net183));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(net187),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_8 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__buf_2 fanout187 (.A(_06661_),
    .X(net187));
 sky130_fd_sc_hd__buf_4 fanout188 (.A(_06661_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_8 fanout189 (.A(_02444_),
    .X(net189));
 sky130_fd_sc_hd__buf_8 fanout19 (.A(_00413_),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(_02444_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(_02442_),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(_02439_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_8 fanout194 (.A(_02436_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(_02428_),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(_02428_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_16 fanout197 (.A(_06737_),
    .X(net197));
 sky130_fd_sc_hd__buf_8 fanout198 (.A(_06737_),
    .X(net198));
 sky130_fd_sc_hd__buf_12 fanout199 (.A(_06736_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_8 fanout2 (.A(_06286_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_8 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_12 fanout200 (.A(_06694_),
    .X(net200));
 sky130_fd_sc_hd__buf_12 fanout201 (.A(_06693_),
    .X(net201));
 sky130_fd_sc_hd__buf_6 fanout202 (.A(_06693_),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_8 fanout204 (.A(_06678_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 fanout205 (.A(_06666_),
    .X(net205));
 sky130_fd_sc_hd__buf_6 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(_06577_),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_8 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(net212),
    .X(net209));
 sky130_fd_sc_hd__buf_8 fanout21 (.A(_00408_),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_8 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_4 fanout212 (.A(_06576_),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_8 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 fanout214 (.A(_06568_),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_8 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(_06561_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 fanout217 (.A(_06560_),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(_06554_),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_8 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_8 fanout220 (.A(_06547_),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_8 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(_06546_),
    .X(net222));
 sky130_fd_sc_hd__buf_4 fanout223 (.A(_06537_),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(_06537_),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_4 fanout226 (.A(_04895_),
    .X(net226));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_2 fanout228 (.A(_02624_),
    .X(net228));
 sky130_fd_sc_hd__buf_4 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_8 fanout23 (.A(_00394_),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_8 fanout230 (.A(_02624_),
    .X(net230));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_8 fanout232 (.A(_02445_),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(_02433_),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_8 fanout234 (.A(_02426_),
    .X(net234));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(_02349_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 fanout236 (.A(_00139_),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_8 fanout237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_8 fanout238 (.A(net241),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_8 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_8 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__buf_8 fanout240 (.A(net241),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_4 fanout241 (.A(_06653_),
    .X(net241));
 sky130_fd_sc_hd__buf_8 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_8 fanout243 (.A(_06652_),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__buf_4 fanout245 (.A(_06536_),
    .X(net245));
 sky130_fd_sc_hd__buf_8 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__buf_6 fanout247 (.A(_04873_),
    .X(net247));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(_04412_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_8 fanout25 (.A(_00388_),
    .X(net25));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net251),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net255),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(net255),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_4 fanout253 (.A(net255),
    .X(net253));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net407),
    .X(net255));
 sky130_fd_sc_hd__buf_4 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_4 fanout257 (.A(_02431_),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_8 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__buf_6 fanout259 (.A(_06683_),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_8 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_8 fanout260 (.A(_06682_),
    .X(net260));
 sky130_fd_sc_hd__buf_4 fanout261 (.A(_06682_),
    .X(net261));
 sky130_fd_sc_hd__buf_8 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__buf_4 fanout263 (.A(_04797_),
    .X(net263));
 sky130_fd_sc_hd__buf_8 fanout264 (.A(_04797_),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_8 fanout265 (.A(_04797_),
    .X(net265));
 sky130_fd_sc_hd__buf_4 fanout266 (.A(_04786_),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_8 fanout267 (.A(_04764_),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__buf_6 fanout269 (.A(_04764_),
    .X(net269));
 sky130_fd_sc_hd__buf_8 fanout27 (.A(_00373_),
    .X(net27));
 sky130_fd_sc_hd__buf_8 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(_04753_),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 fanout273 (.A(net282),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net282),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_4 fanout275 (.A(net282),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net282),
    .X(net276));
 sky130_fd_sc_hd__buf_2 fanout277 (.A(net282),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__buf_2 fanout279 (.A(net282),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_8 fanout28 (.A(_00367_),
    .X(net28));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_4 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(_04630_),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_8 fanout283 (.A(_04609_),
    .X(net283));
 sky130_fd_sc_hd__buf_2 fanout284 (.A(_04609_),
    .X(net284));
 sky130_fd_sc_hd__buf_6 fanout285 (.A(_04456_),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 fanout286 (.A(_04456_),
    .X(net286));
 sky130_fd_sc_hd__buf_6 fanout287 (.A(reg1_val[7]),
    .X(net287));
 sky130_fd_sc_hd__buf_8 fanout288 (.A(reg1_val[30]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_8 fanout289 (.A(reg1_val[1]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_8 fanout29 (.A(_00367_),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_8 fanout290 (.A(reg1_val[11]),
    .X(net290));
 sky130_fd_sc_hd__buf_8 fanout291 (.A(reg1_val[0]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_8 fanout292 (.A(reg1_val[0]),
    .X(net292));
 sky130_fd_sc_hd__buf_4 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_4 fanout294 (.A(net296),
    .X(net294));
 sky130_fd_sc_hd__buf_4 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_4 fanout296 (.A(instruction[7]),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_8 fanout297 (.A(instruction[6]),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_8 fanout298 (.A(instruction[4]),
    .X(net298));
 sky130_fd_sc_hd__buf_6 fanout3 (.A(net4),
    .X(net3));
 sky130_fd_sc_hd__buf_6 fanout30 (.A(_00341_),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout31 (.A(_00341_),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_8 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_6 fanout33 (.A(_00321_),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_8 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_8 fanout35 (.A(_00317_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_8 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_8 fanout37 (.A(_00288_),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_8 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_8 fanout39 (.A(_00282_),
    .X(net39));
 sky130_fd_sc_hd__buf_8 fanout4 (.A(_02188_),
    .X(net4));
 sky130_fd_sc_hd__buf_6 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 fanout41 (.A(_00209_),
    .X(net41));
 sky130_fd_sc_hd__buf_8 fanout42 (.A(_00202_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_8 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_4 fanout44 (.A(_00176_),
    .X(net44));
 sky130_fd_sc_hd__buf_6 fanout45 (.A(_00162_),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(_00162_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_8 fanout47 (.A(_00149_),
    .X(net47));
 sky130_fd_sc_hd__buf_4 fanout48 (.A(_00149_),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_8 fanout49 (.A(_00143_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 fanout5 (.A(_02176_),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(_00143_),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_8 fanout51 (.A(_00137_),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(_00137_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_8 fanout53 (.A(_06731_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(_06731_),
    .X(net54));
 sky130_fd_sc_hd__buf_6 fanout56 (.A(_06724_),
    .X(net56));
 sky130_fd_sc_hd__buf_4 fanout57 (.A(_06724_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_8 fanout58 (.A(net60),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_8 fanout59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout6 (.A(_02175_),
    .X(net6));
 sky130_fd_sc_hd__buf_8 fanout60 (.A(_02186_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 fanout61 (.A(net63),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_8 fanout63 (.A(_02185_),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_16 fanout64 (.A(net65),
    .X(net64));
 sky130_fd_sc_hd__buf_12 fanout65 (.A(_00788_),
    .X(net65));
 sky130_fd_sc_hd__buf_6 fanout66 (.A(net67),
    .X(net66));
 sky130_fd_sc_hd__buf_6 fanout67 (.A(_00497_),
    .X(net67));
 sky130_fd_sc_hd__buf_6 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__buf_6 fanout69 (.A(_00496_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_8 fanout7 (.A(_02175_),
    .X(net7));
 sky130_fd_sc_hd__buf_8 fanout70 (.A(_00468_),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_16 fanout71 (.A(_00467_),
    .X(net71));
 sky130_fd_sc_hd__buf_8 fanout72 (.A(_00466_),
    .X(net72));
 sky130_fd_sc_hd__buf_8 fanout74 (.A(_00463_),
    .X(net74));
 sky130_fd_sc_hd__buf_8 fanout75 (.A(_00460_),
    .X(net75));
 sky130_fd_sc_hd__buf_6 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_8 fanout77 (.A(_00447_),
    .X(net77));
 sky130_fd_sc_hd__buf_6 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_8 fanout8 (.A(net9),
    .X(net8));
 sky130_fd_sc_hd__buf_8 fanout80 (.A(_00444_),
    .X(net80));
 sky130_fd_sc_hd__buf_8 fanout82 (.A(_00442_),
    .X(net82));
 sky130_fd_sc_hd__buf_6 fanout83 (.A(net84),
    .X(net83));
 sky130_fd_sc_hd__buf_8 fanout84 (.A(_00440_),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_8 fanout85 (.A(_00398_),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_16 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_16 fanout87 (.A(_00358_),
    .X(net87));
 sky130_fd_sc_hd__buf_12 fanout88 (.A(net90),
    .X(net88));
 sky130_fd_sc_hd__buf_8 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_6 fanout9 (.A(_02080_),
    .X(net9));
 sky130_fd_sc_hd__buf_6 fanout90 (.A(_00353_),
    .X(net90));
 sky130_fd_sc_hd__buf_12 fanout91 (.A(_00309_),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_16 fanout92 (.A(_00308_),
    .X(net92));
 sky130_fd_sc_hd__buf_8 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_8 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_16 fanout95 (.A(_00301_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_16 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__buf_12 fanout97 (.A(_00273_),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_16 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__buf_12 fanout99 (.A(_00262_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\div_shifter[1] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_00004_),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_00071_),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\div_shifter[3] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_06329_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\divi2_l[23] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_06156_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\divi2_l[10] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_06140_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net434),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_06344_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(busy_l),
    .X(net407));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold11 (.A(\divi2_l[1] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_06356_),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\divi2_l[9] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_06139_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\div_shifter[19] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_06348_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_00085_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\divi2_l[19] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_06151_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\divi2_l[24] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_06157_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_00003_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\div_shifter[11] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_06340_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_00078_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\div_shifter[30] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_06362_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_00097_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\divi2_l[16] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_06148_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\div_shifter[4] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_06330_),
    .X(net427));
 sky130_fd_sc_hd__buf_1 hold13 (.A(\divi2_l[0] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\div_shifter[24] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_06354_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\div_shifter[14] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_06342_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\divi2_l[20] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_06152_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\div_shifter[15] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_06343_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\div_shifter[20] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_06349_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00002_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\div_shifter[63] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_06491_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_00129_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\div_counter[4] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_06501_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_00134_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\div_shifter[22] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_06352_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_00088_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\div_shifter[0] ),
    .X(net447));
 sky130_fd_sc_hd__buf_1 hold15 (.A(\div_counter[3] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_06325_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\div_shifter[18] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_06347_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_00084_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\div_res[31] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_06324_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_00065_),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\div_shifter[10] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_06338_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(div_complete),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_00133_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_00135_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\div_shifter[6] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_06332_),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\div_res[8] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_06298_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_00043_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\div_res[26] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_06319_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_00061_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\div_counter[2] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(divi1_sign),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_06497_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_00132_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\divi2_l[31] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_06166_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\div_res[21] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_06313_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_00056_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(net510),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_06311_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_00054_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_06127_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\div_res[7] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_06296_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\div_res[5] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_06293_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_00039_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(net501),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_06310_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_00053_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\div_res[0] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_06288_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\div_shifter[9] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_00035_),
    .X(net488));
 sky130_fd_sc_hd__buf_1 hold191 (.A(net516),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_06123_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\div_res[14] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_06304_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\div_res[15] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_06305_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\div_res[29] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_06322_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_00063_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_00067_),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_06337_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\div_res[17] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_06307_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_00051_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\div_res[18] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_06308_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net527),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_06314_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\div_res[25] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_06318_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\div_res[11] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_00076_),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_06300_),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_00045_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\div_res[20] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(_06312_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\div_res[12] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_06301_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\div_res[24] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_06317_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\div_counter[0] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\div_res[28] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\div_shifter[16] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_06320_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_00062_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net535),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_06294_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\div_res[30] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_06323_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\div_res[3] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_06290_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_00037_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\div_res[23] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_06346_),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_06316_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\div_res[16] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_06306_),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\div_shifter[62] ),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_2 hold234 (.A(_06286_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\div_res[13] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_06302_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\div_res[6] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\div_res[4] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(_06292_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_00083_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\div_res[9] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(_06299_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_00044_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\div_res[2] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_06289_),
    .X(net542));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold245 (.A(\div_shifter[32] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_06366_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\div_shifter[60] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_06480_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\div_shifter[59] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\div_shifter[27] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_06475_),
    .X(net548));
 sky130_fd_sc_hd__buf_1 hold251 (.A(net598),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_06427_),
    .X(net550));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold253 (.A(\div_shifter[41] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_06404_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\div_shifter[54] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_06456_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\div_shifter[49] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_06438_),
    .X(net556));
 sky130_fd_sc_hd__buf_1 hold259 (.A(\div_shifter[50] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_06359_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_06441_),
    .X(net558));
 sky130_fd_sc_hd__buf_1 hold261 (.A(net596),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\div_shifter[33] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_00099_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\div_shifter[35] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_06379_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\div_shifter[53] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_06453_),
    .X(net565));
 sky130_fd_sc_hd__buf_1 hold268 (.A(net597),
    .X(net566));
 sky130_fd_sc_hd__buf_1 hold269 (.A(\div_shifter[56] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_00094_),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_06464_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\div_shifter[44] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_06418_),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\div_shifter[58] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_06471_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\div_shifter[52] ),
    .X(net573));
 sky130_fd_sc_hd__buf_1 hold276 (.A(net599),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_06395_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\div_shifter[57] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(_06467_),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\divi2_l[28] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\div_shifter[42] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_06409_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\div_shifter[55] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\div_shifter[36] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_06383_),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\div_shifter[34] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_06375_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\div_shifter[38] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_06391_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\div_shifter[45] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_06162_),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_06422_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\div_shifter[43] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\div_shifter[48] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(_06434_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\div_shifter[37] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\div_shifter[40] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\div_shifter[47] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\div_res[13] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\div_shifter[51] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\div_shifter[61] ),
    .X(net597));
 sky130_fd_sc_hd__buf_1 hold3 (.A(\div_counter[1] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\divi2_l[29] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\div_shifter[46] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\div_shifter[39] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_06163_),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\div_shifter[29] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_06361_),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_00096_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\divi2_l[6] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_06136_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\divi2_l[18] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_06150_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\divi2_l[25] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_00131_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_06158_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_00027_),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\divi2_l[27] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_06161_),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\divi2_l[30] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_06164_),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\divi2_l[26] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_06160_),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\divi2_l[22] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_06155_),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\div_shifter[7] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_00024_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\divi2_l[12] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_06143_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\div_shifter[26] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_06358_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\divi2_l[17] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_06149_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\divi2_l[13] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_06144_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net436),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_00073_),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_06350_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_00087_),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\divi2_l[11] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_06142_),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net386),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_06336_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\divi2_l[14] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_06145_),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\divi2_l[8] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_06138_),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\divi2_l[3] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\div_shifter[23] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_06353_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_00089_),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\divi2_l[7] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_06137_),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_00009_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\div_shifter[2] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_06328_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\divi2_l[5] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_06134_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_00005_),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_00007_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\div_shifter[28] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_06360_),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\divi2_l[4] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_06133_),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\divi2_l[21] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_06154_),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_00023_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\div_shifter[8] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_06335_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\divi2_l[2] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\divi2_l[15] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_06146_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\div_shifter[13] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_06341_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_00079_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\div_shifter[25] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_06355_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_00091_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\div_shifter[5] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_06331_),
    .X(net397));
 sky130_fd_sc_hd__buf_6 max_cap102 (.A(_00220_),
    .X(net102));
 sky130_fd_sc_hd__buf_6 max_cap107 (.A(_00476_),
    .X(net107));
 sky130_fd_sc_hd__buf_4 max_cap11 (.A(_02065_),
    .X(net11));
 sky130_fd_sc_hd__buf_6 max_cap112 (.A(_00412_),
    .X(net112));
 sky130_fd_sc_hd__buf_6 max_cap114 (.A(_00392_),
    .X(net114));
 sky130_fd_sc_hd__buf_4 max_cap121 (.A(_00375_),
    .X(net121));
 sky130_fd_sc_hd__buf_6 max_cap148 (.A(_00340_),
    .X(net148));
 sky130_fd_sc_hd__buf_6 max_cap153 (.A(_00319_),
    .X(net153));
 sky130_fd_sc_hd__buf_2 max_cap173 (.A(_00247_),
    .X(net173));
 sky130_fd_sc_hd__buf_1 max_cap176 (.A(_06711_),
    .X(net176));
 sky130_fd_sc_hd__buf_4 max_cap55 (.A(_06730_),
    .X(net55));
 sky130_fd_sc_hd__buf_6 max_cap73 (.A(_00464_),
    .X(net73));
 sky130_fd_sc_hd__buf_6 max_cap78 (.A(_00446_),
    .X(net78));
 sky130_fd_sc_hd__buf_6 max_cap81 (.A(_00443_),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_8 wire101 (.A(_00229_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 wire122 (.A(_00372_),
    .X(net122));
endmodule

