VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multiplexer
  CLASS BLOCK ;
  FOREIGN multiplexer ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 1000.000 ;
  PIN custom_settings[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END custom_settings[0]
  PIN custom_settings[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END custom_settings[10]
  PIN custom_settings[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 186.360 4.000 186.960 ;
    END
  END custom_settings[11]
  PIN custom_settings[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END custom_settings[12]
  PIN custom_settings[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END custom_settings[13]
  PIN custom_settings[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 4.000 195.120 ;
    END
  END custom_settings[14]
  PIN custom_settings[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END custom_settings[15]
  PIN custom_settings[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END custom_settings[16]
  PIN custom_settings[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END custom_settings[17]
  PIN custom_settings[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END custom_settings[18]
  PIN custom_settings[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END custom_settings[19]
  PIN custom_settings[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END custom_settings[1]
  PIN custom_settings[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END custom_settings[20]
  PIN custom_settings[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END custom_settings[21]
  PIN custom_settings[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END custom_settings[22]
  PIN custom_settings[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END custom_settings[23]
  PIN custom_settings[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END custom_settings[24]
  PIN custom_settings[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END custom_settings[25]
  PIN custom_settings[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END custom_settings[26]
  PIN custom_settings[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END custom_settings[27]
  PIN custom_settings[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END custom_settings[28]
  PIN custom_settings[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END custom_settings[29]
  PIN custom_settings[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END custom_settings[2]
  PIN custom_settings[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END custom_settings[30]
  PIN custom_settings[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.760 4.000 241.360 ;
    END
  END custom_settings[31]
  PIN custom_settings[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END custom_settings[3]
  PIN custom_settings[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END custom_settings[4]
  PIN custom_settings[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END custom_settings[5]
  PIN custom_settings[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END custom_settings[6]
  PIN custom_settings[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END custom_settings[7]
  PIN custom_settings[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END custom_settings[8]
  PIN custom_settings[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END custom_settings[9]
  PIN io_in_0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 3.770 996.000 4.050 1000.000 ;
    END
  END io_in_0
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 4.000 282.160 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 314.200 4.000 314.800 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END io_oeb[9]
  PIN io_oeb_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END io_oeb_scrapcpu[0]
  PIN io_oeb_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END io_oeb_scrapcpu[10]
  PIN io_oeb_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END io_oeb_scrapcpu[11]
  PIN io_oeb_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END io_oeb_scrapcpu[12]
  PIN io_oeb_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END io_oeb_scrapcpu[13]
  PIN io_oeb_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END io_oeb_scrapcpu[14]
  PIN io_oeb_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END io_oeb_scrapcpu[15]
  PIN io_oeb_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END io_oeb_scrapcpu[16]
  PIN io_oeb_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END io_oeb_scrapcpu[17]
  PIN io_oeb_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END io_oeb_scrapcpu[18]
  PIN io_oeb_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END io_oeb_scrapcpu[19]
  PIN io_oeb_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 553.560 4.000 554.160 ;
    END
  END io_oeb_scrapcpu[1]
  PIN io_oeb_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END io_oeb_scrapcpu[20]
  PIN io_oeb_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END io_oeb_scrapcpu[21]
  PIN io_oeb_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END io_oeb_scrapcpu[22]
  PIN io_oeb_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END io_oeb_scrapcpu[23]
  PIN io_oeb_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END io_oeb_scrapcpu[24]
  PIN io_oeb_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END io_oeb_scrapcpu[25]
  PIN io_oeb_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END io_oeb_scrapcpu[26]
  PIN io_oeb_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.280 4.000 624.880 ;
    END
  END io_oeb_scrapcpu[27]
  PIN io_oeb_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END io_oeb_scrapcpu[28]
  PIN io_oeb_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END io_oeb_scrapcpu[29]
  PIN io_oeb_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END io_oeb_scrapcpu[2]
  PIN io_oeb_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END io_oeb_scrapcpu[30]
  PIN io_oeb_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.160 4.000 635.760 ;
    END
  END io_oeb_scrapcpu[31]
  PIN io_oeb_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END io_oeb_scrapcpu[32]
  PIN io_oeb_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 640.600 4.000 641.200 ;
    END
  END io_oeb_scrapcpu[33]
  PIN io_oeb_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END io_oeb_scrapcpu[34]
  PIN io_oeb_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END io_oeb_scrapcpu[35]
  PIN io_oeb_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END io_oeb_scrapcpu[3]
  PIN io_oeb_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END io_oeb_scrapcpu[4]
  PIN io_oeb_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END io_oeb_scrapcpu[5]
  PIN io_oeb_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END io_oeb_scrapcpu[6]
  PIN io_oeb_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END io_oeb_scrapcpu[7]
  PIN io_oeb_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END io_oeb_scrapcpu[8]
  PIN io_oeb_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END io_oeb_scrapcpu[9]
  PIN io_oeb_vliw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 746.680 4.000 747.280 ;
    END
  END io_oeb_vliw[0]
  PIN io_oeb_vliw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.880 4.000 774.480 ;
    END
  END io_oeb_vliw[10]
  PIN io_oeb_vliw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END io_oeb_vliw[11]
  PIN io_oeb_vliw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END io_oeb_vliw[12]
  PIN io_oeb_vliw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END io_oeb_vliw[13]
  PIN io_oeb_vliw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END io_oeb_vliw[14]
  PIN io_oeb_vliw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 787.480 4.000 788.080 ;
    END
  END io_oeb_vliw[15]
  PIN io_oeb_vliw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 790.200 4.000 790.800 ;
    END
  END io_oeb_vliw[16]
  PIN io_oeb_vliw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END io_oeb_vliw[17]
  PIN io_oeb_vliw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END io_oeb_vliw[18]
  PIN io_oeb_vliw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 798.360 4.000 798.960 ;
    END
  END io_oeb_vliw[19]
  PIN io_oeb_vliw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END io_oeb_vliw[1]
  PIN io_oeb_vliw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END io_oeb_vliw[20]
  PIN io_oeb_vliw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.800 4.000 804.400 ;
    END
  END io_oeb_vliw[21]
  PIN io_oeb_vliw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 806.520 4.000 807.120 ;
    END
  END io_oeb_vliw[22]
  PIN io_oeb_vliw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END io_oeb_vliw[23]
  PIN io_oeb_vliw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 4.000 812.560 ;
    END
  END io_oeb_vliw[24]
  PIN io_oeb_vliw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 814.680 4.000 815.280 ;
    END
  END io_oeb_vliw[25]
  PIN io_oeb_vliw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END io_oeb_vliw[26]
  PIN io_oeb_vliw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 820.120 4.000 820.720 ;
    END
  END io_oeb_vliw[27]
  PIN io_oeb_vliw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END io_oeb_vliw[28]
  PIN io_oeb_vliw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END io_oeb_vliw[29]
  PIN io_oeb_vliw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END io_oeb_vliw[2]
  PIN io_oeb_vliw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 828.280 4.000 828.880 ;
    END
  END io_oeb_vliw[30]
  PIN io_oeb_vliw[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 831.000 4.000 831.600 ;
    END
  END io_oeb_vliw[31]
  PIN io_oeb_vliw[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.720 4.000 834.320 ;
    END
  END io_oeb_vliw[32]
  PIN io_oeb_vliw[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END io_oeb_vliw[33]
  PIN io_oeb_vliw[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END io_oeb_vliw[34]
  PIN io_oeb_vliw[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.880 4.000 842.480 ;
    END
  END io_oeb_vliw[35]
  PIN io_oeb_vliw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END io_oeb_vliw[3]
  PIN io_oeb_vliw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END io_oeb_vliw[4]
  PIN io_oeb_vliw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END io_oeb_vliw[5]
  PIN io_oeb_vliw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END io_oeb_vliw[6]
  PIN io_oeb_vliw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END io_oeb_vliw[7]
  PIN io_oeb_vliw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END io_oeb_vliw[8]
  PIN io_oeb_vliw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.160 4.000 771.760 ;
    END
  END io_oeb_vliw[9]
  PIN io_oeb_z80[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END io_oeb_z80[0]
  PIN io_oeb_z80[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END io_oeb_z80[10]
  PIN io_oeb_z80[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END io_oeb_z80[11]
  PIN io_oeb_z80[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END io_oeb_z80[12]
  PIN io_oeb_z80[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END io_oeb_z80[13]
  PIN io_oeb_z80[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END io_oeb_z80[14]
  PIN io_oeb_z80[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END io_oeb_z80[15]
  PIN io_oeb_z80[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.280 4.000 692.880 ;
    END
  END io_oeb_z80[16]
  PIN io_oeb_z80[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END io_oeb_z80[17]
  PIN io_oeb_z80[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END io_oeb_z80[18]
  PIN io_oeb_z80[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END io_oeb_z80[19]
  PIN io_oeb_z80[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END io_oeb_z80[1]
  PIN io_oeb_z80[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END io_oeb_z80[20]
  PIN io_oeb_z80[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END io_oeb_z80[21]
  PIN io_oeb_z80[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END io_oeb_z80[22]
  PIN io_oeb_z80[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END io_oeb_z80[23]
  PIN io_oeb_z80[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END io_oeb_z80[24]
  PIN io_oeb_z80[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END io_oeb_z80[25]
  PIN io_oeb_z80[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END io_oeb_z80[26]
  PIN io_oeb_z80[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END io_oeb_z80[27]
  PIN io_oeb_z80[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END io_oeb_z80[28]
  PIN io_oeb_z80[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END io_oeb_z80[29]
  PIN io_oeb_z80[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END io_oeb_z80[2]
  PIN io_oeb_z80[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 730.360 4.000 730.960 ;
    END
  END io_oeb_z80[30]
  PIN io_oeb_z80[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END io_oeb_z80[31]
  PIN io_oeb_z80[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END io_oeb_z80[32]
  PIN io_oeb_z80[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 738.520 4.000 739.120 ;
    END
  END io_oeb_z80[33]
  PIN io_oeb_z80[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END io_oeb_z80[34]
  PIN io_oeb_z80[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END io_oeb_z80[35]
  PIN io_oeb_z80[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END io_oeb_z80[3]
  PIN io_oeb_z80[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END io_oeb_z80[4]
  PIN io_oeb_z80[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END io_oeb_z80[5]
  PIN io_oeb_z80[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END io_oeb_z80[6]
  PIN io_oeb_z80[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END io_oeb_z80[7]
  PIN io_oeb_z80[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END io_oeb_z80[8]
  PIN io_oeb_z80[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END io_oeb_z80[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 5.480 200.000 6.080 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 73.480 200.000 74.080 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 80.280 200.000 80.880 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 87.080 200.000 87.680 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 93.880 200.000 94.480 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 100.680 200.000 101.280 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 107.480 200.000 108.080 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 114.280 200.000 114.880 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 121.080 200.000 121.680 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 127.880 200.000 128.480 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 134.680 200.000 135.280 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 12.280 200.000 12.880 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 141.480 200.000 142.080 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 148.280 200.000 148.880 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 155.080 200.000 155.680 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 161.880 200.000 162.480 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 168.680 200.000 169.280 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 175.480 200.000 176.080 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 182.280 200.000 182.880 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 189.080 200.000 189.680 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 195.880 200.000 196.480 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 202.680 200.000 203.280 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 19.080 200.000 19.680 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 209.480 200.000 210.080 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 216.280 200.000 216.880 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 223.080 200.000 223.680 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 229.880 200.000 230.480 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 236.680 200.000 237.280 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 243.480 200.000 244.080 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 250.280 200.000 250.880 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 257.080 200.000 257.680 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 25.880 200.000 26.480 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 32.680 200.000 33.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 39.480 200.000 40.080 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 46.280 200.000 46.880 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 53.080 200.000 53.680 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 59.880 200.000 60.480 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 66.680 200.000 67.280 ;
    END
  END io_out[9]
  PIN io_out_scrapcpu[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END io_out_scrapcpu[0]
  PIN io_out_scrapcpu[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END io_out_scrapcpu[10]
  PIN io_out_scrapcpu[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END io_out_scrapcpu[11]
  PIN io_out_scrapcpu[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.200 4.000 382.800 ;
    END
  END io_out_scrapcpu[12]
  PIN io_out_scrapcpu[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END io_out_scrapcpu[13]
  PIN io_out_scrapcpu[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END io_out_scrapcpu[14]
  PIN io_out_scrapcpu[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END io_out_scrapcpu[15]
  PIN io_out_scrapcpu[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END io_out_scrapcpu[16]
  PIN io_out_scrapcpu[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END io_out_scrapcpu[17]
  PIN io_out_scrapcpu[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END io_out_scrapcpu[18]
  PIN io_out_scrapcpu[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END io_out_scrapcpu[19]
  PIN io_out_scrapcpu[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END io_out_scrapcpu[1]
  PIN io_out_scrapcpu[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END io_out_scrapcpu[20]
  PIN io_out_scrapcpu[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END io_out_scrapcpu[21]
  PIN io_out_scrapcpu[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END io_out_scrapcpu[22]
  PIN io_out_scrapcpu[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END io_out_scrapcpu[23]
  PIN io_out_scrapcpu[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END io_out_scrapcpu[24]
  PIN io_out_scrapcpu[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END io_out_scrapcpu[25]
  PIN io_out_scrapcpu[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.280 4.000 420.880 ;
    END
  END io_out_scrapcpu[26]
  PIN io_out_scrapcpu[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END io_out_scrapcpu[27]
  PIN io_out_scrapcpu[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END io_out_scrapcpu[28]
  PIN io_out_scrapcpu[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END io_out_scrapcpu[29]
  PIN io_out_scrapcpu[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.000 4.000 355.600 ;
    END
  END io_out_scrapcpu[2]
  PIN io_out_scrapcpu[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END io_out_scrapcpu[30]
  PIN io_out_scrapcpu[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END io_out_scrapcpu[31]
  PIN io_out_scrapcpu[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END io_out_scrapcpu[32]
  PIN io_out_scrapcpu[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END io_out_scrapcpu[33]
  PIN io_out_scrapcpu[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END io_out_scrapcpu[34]
  PIN io_out_scrapcpu[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END io_out_scrapcpu[35]
  PIN io_out_scrapcpu[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END io_out_scrapcpu[3]
  PIN io_out_scrapcpu[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END io_out_scrapcpu[4]
  PIN io_out_scrapcpu[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END io_out_scrapcpu[5]
  PIN io_out_scrapcpu[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END io_out_scrapcpu[6]
  PIN io_out_scrapcpu[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END io_out_scrapcpu[7]
  PIN io_out_scrapcpu[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END io_out_scrapcpu[8]
  PIN io_out_scrapcpu[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END io_out_scrapcpu[9]
  PIN io_out_vliw[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 18.950 996.000 19.230 1000.000 ;
    END
  END io_out_vliw[0]
  PIN io_out_vliw[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 69.550 996.000 69.830 1000.000 ;
    END
  END io_out_vliw[10]
  PIN io_out_vliw[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 74.610 996.000 74.890 1000.000 ;
    END
  END io_out_vliw[11]
  PIN io_out_vliw[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 79.670 996.000 79.950 1000.000 ;
    END
  END io_out_vliw[12]
  PIN io_out_vliw[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 84.730 996.000 85.010 1000.000 ;
    END
  END io_out_vliw[13]
  PIN io_out_vliw[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 89.790 996.000 90.070 1000.000 ;
    END
  END io_out_vliw[14]
  PIN io_out_vliw[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 94.850 996.000 95.130 1000.000 ;
    END
  END io_out_vliw[15]
  PIN io_out_vliw[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 996.000 100.190 1000.000 ;
    END
  END io_out_vliw[16]
  PIN io_out_vliw[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 104.970 996.000 105.250 1000.000 ;
    END
  END io_out_vliw[17]
  PIN io_out_vliw[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 110.030 996.000 110.310 1000.000 ;
    END
  END io_out_vliw[18]
  PIN io_out_vliw[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 115.090 996.000 115.370 1000.000 ;
    END
  END io_out_vliw[19]
  PIN io_out_vliw[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 24.010 996.000 24.290 1000.000 ;
    END
  END io_out_vliw[1]
  PIN io_out_vliw[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 996.000 120.430 1000.000 ;
    END
  END io_out_vliw[20]
  PIN io_out_vliw[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 125.210 996.000 125.490 1000.000 ;
    END
  END io_out_vliw[21]
  PIN io_out_vliw[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 130.270 996.000 130.550 1000.000 ;
    END
  END io_out_vliw[22]
  PIN io_out_vliw[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 135.330 996.000 135.610 1000.000 ;
    END
  END io_out_vliw[23]
  PIN io_out_vliw[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 140.390 996.000 140.670 1000.000 ;
    END
  END io_out_vliw[24]
  PIN io_out_vliw[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 145.450 996.000 145.730 1000.000 ;
    END
  END io_out_vliw[25]
  PIN io_out_vliw[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 150.510 996.000 150.790 1000.000 ;
    END
  END io_out_vliw[26]
  PIN io_out_vliw[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 155.570 996.000 155.850 1000.000 ;
    END
  END io_out_vliw[27]
  PIN io_out_vliw[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 160.630 996.000 160.910 1000.000 ;
    END
  END io_out_vliw[28]
  PIN io_out_vliw[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 165.690 996.000 165.970 1000.000 ;
    END
  END io_out_vliw[29]
  PIN io_out_vliw[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 996.000 29.350 1000.000 ;
    END
  END io_out_vliw[2]
  PIN io_out_vliw[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 170.750 996.000 171.030 1000.000 ;
    END
  END io_out_vliw[30]
  PIN io_out_vliw[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 175.810 996.000 176.090 1000.000 ;
    END
  END io_out_vliw[31]
  PIN io_out_vliw[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 180.870 996.000 181.150 1000.000 ;
    END
  END io_out_vliw[32]
  PIN io_out_vliw[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 185.930 996.000 186.210 1000.000 ;
    END
  END io_out_vliw[33]
  PIN io_out_vliw[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 190.990 996.000 191.270 1000.000 ;
    END
  END io_out_vliw[34]
  PIN io_out_vliw[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 196.050 996.000 196.330 1000.000 ;
    END
  END io_out_vliw[35]
  PIN io_out_vliw[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 34.130 996.000 34.410 1000.000 ;
    END
  END io_out_vliw[3]
  PIN io_out_vliw[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 39.190 996.000 39.470 1000.000 ;
    END
  END io_out_vliw[4]
  PIN io_out_vliw[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 44.250 996.000 44.530 1000.000 ;
    END
  END io_out_vliw[5]
  PIN io_out_vliw[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 49.310 996.000 49.590 1000.000 ;
    END
  END io_out_vliw[6]
  PIN io_out_vliw[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 54.370 996.000 54.650 1000.000 ;
    END
  END io_out_vliw[7]
  PIN io_out_vliw[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 59.430 996.000 59.710 1000.000 ;
    END
  END io_out_vliw[8]
  PIN io_out_vliw[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 996.000 64.770 1000.000 ;
    END
  END io_out_vliw[9]
  PIN io_out_z80[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 753.480 200.000 754.080 ;
    END
  END io_out_z80[0]
  PIN io_out_z80[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 821.480 200.000 822.080 ;
    END
  END io_out_z80[10]
  PIN io_out_z80[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 828.280 200.000 828.880 ;
    END
  END io_out_z80[11]
  PIN io_out_z80[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 835.080 200.000 835.680 ;
    END
  END io_out_z80[12]
  PIN io_out_z80[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 841.880 200.000 842.480 ;
    END
  END io_out_z80[13]
  PIN io_out_z80[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 848.680 200.000 849.280 ;
    END
  END io_out_z80[14]
  PIN io_out_z80[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 855.480 200.000 856.080 ;
    END
  END io_out_z80[15]
  PIN io_out_z80[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 862.280 200.000 862.880 ;
    END
  END io_out_z80[16]
  PIN io_out_z80[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 869.080 200.000 869.680 ;
    END
  END io_out_z80[17]
  PIN io_out_z80[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 875.880 200.000 876.480 ;
    END
  END io_out_z80[18]
  PIN io_out_z80[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 882.680 200.000 883.280 ;
    END
  END io_out_z80[19]
  PIN io_out_z80[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 760.280 200.000 760.880 ;
    END
  END io_out_z80[1]
  PIN io_out_z80[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 889.480 200.000 890.080 ;
    END
  END io_out_z80[20]
  PIN io_out_z80[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 896.280 200.000 896.880 ;
    END
  END io_out_z80[21]
  PIN io_out_z80[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 903.080 200.000 903.680 ;
    END
  END io_out_z80[22]
  PIN io_out_z80[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 909.880 200.000 910.480 ;
    END
  END io_out_z80[23]
  PIN io_out_z80[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 916.680 200.000 917.280 ;
    END
  END io_out_z80[24]
  PIN io_out_z80[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 923.480 200.000 924.080 ;
    END
  END io_out_z80[25]
  PIN io_out_z80[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 930.280 200.000 930.880 ;
    END
  END io_out_z80[26]
  PIN io_out_z80[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 937.080 200.000 937.680 ;
    END
  END io_out_z80[27]
  PIN io_out_z80[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 943.880 200.000 944.480 ;
    END
  END io_out_z80[28]
  PIN io_out_z80[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 950.680 200.000 951.280 ;
    END
  END io_out_z80[29]
  PIN io_out_z80[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 767.080 200.000 767.680 ;
    END
  END io_out_z80[2]
  PIN io_out_z80[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 957.480 200.000 958.080 ;
    END
  END io_out_z80[30]
  PIN io_out_z80[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 964.280 200.000 964.880 ;
    END
  END io_out_z80[31]
  PIN io_out_z80[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 971.080 200.000 971.680 ;
    END
  END io_out_z80[32]
  PIN io_out_z80[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 977.880 200.000 978.480 ;
    END
  END io_out_z80[33]
  PIN io_out_z80[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 984.680 200.000 985.280 ;
    END
  END io_out_z80[34]
  PIN io_out_z80[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 991.480 200.000 992.080 ;
    END
  END io_out_z80[35]
  PIN io_out_z80[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 773.880 200.000 774.480 ;
    END
  END io_out_z80[3]
  PIN io_out_z80[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 780.680 200.000 781.280 ;
    END
  END io_out_z80[4]
  PIN io_out_z80[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 787.480 200.000 788.080 ;
    END
  END io_out_z80[5]
  PIN io_out_z80[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 794.280 200.000 794.880 ;
    END
  END io_out_z80[6]
  PIN io_out_z80[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 801.080 200.000 801.680 ;
    END
  END io_out_z80[7]
  PIN io_out_z80[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 807.880 200.000 808.480 ;
    END
  END io_out_z80[8]
  PIN io_out_z80[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 196.000 814.680 200.000 815.280 ;
    END
  END io_out_z80[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 481.480 200.000 482.080 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 549.480 200.000 550.080 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 556.280 200.000 556.880 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 563.080 200.000 563.680 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 569.880 200.000 570.480 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 576.680 200.000 577.280 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 583.480 200.000 584.080 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 590.280 200.000 590.880 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 597.080 200.000 597.680 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 603.880 200.000 604.480 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 610.680 200.000 611.280 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 488.280 200.000 488.880 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 617.480 200.000 618.080 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 624.280 200.000 624.880 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 631.080 200.000 631.680 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 637.880 200.000 638.480 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 644.680 200.000 645.280 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 651.480 200.000 652.080 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 658.280 200.000 658.880 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 665.080 200.000 665.680 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 671.880 200.000 672.480 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 678.680 200.000 679.280 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 495.080 200.000 495.680 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 685.480 200.000 686.080 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 692.280 200.000 692.880 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 699.080 200.000 699.680 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 705.880 200.000 706.480 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 712.680 200.000 713.280 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 719.480 200.000 720.080 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 726.280 200.000 726.880 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 733.080 200.000 733.680 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 739.880 200.000 740.480 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 746.680 200.000 747.280 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 501.880 200.000 502.480 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 508.680 200.000 509.280 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 515.480 200.000 516.080 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 522.280 200.000 522.880 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 529.080 200.000 529.680 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 535.880 200.000 536.480 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 542.680 200.000 543.280 ;
    END
  END la_data_out[9]
  PIN rst_scrapcpu
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END rst_scrapcpu
  PIN rst_vliw
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 8.830 996.000 9.110 1000.000 ;
    END
  END rst_vliw
  PIN rst_z80
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 13.890 996.000 14.170 1000.000 ;
    END
  END rst_z80
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.470 0.000 162.750 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 18.950 0.000 19.230 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 0.000 192.650 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.920 4.000 453.520 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.120 4.000 480.720 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 504.600 4.000 505.200 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 534.520 4.000 535.120 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 263.880 200.000 264.480 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 331.880 200.000 332.480 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 338.680 200.000 339.280 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 345.480 200.000 346.080 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 352.280 200.000 352.880 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 359.080 200.000 359.680 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 365.880 200.000 366.480 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 372.680 200.000 373.280 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 379.480 200.000 380.080 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 386.280 200.000 386.880 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 393.080 200.000 393.680 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 270.680 200.000 271.280 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 399.880 200.000 400.480 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 406.680 200.000 407.280 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 413.480 200.000 414.080 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 420.280 200.000 420.880 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 427.080 200.000 427.680 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 433.880 200.000 434.480 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 440.680 200.000 441.280 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 447.480 200.000 448.080 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 454.280 200.000 454.880 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 461.080 200.000 461.680 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 277.480 200.000 278.080 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 467.880 200.000 468.480 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 474.680 200.000 475.280 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 284.280 200.000 284.880 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 291.080 200.000 291.680 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 297.880 200.000 298.480 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 304.680 200.000 305.280 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 311.480 200.000 312.080 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 318.280 200.000 318.880 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 325.080 200.000 325.680 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 545.400 4.000 546.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 987.445 ;
      LAYER met1 ;
        RECT 0.070 10.640 199.570 987.600 ;
      LAYER met2 ;
        RECT 0.100 995.720 3.490 996.610 ;
        RECT 4.330 995.720 8.550 996.610 ;
        RECT 9.390 995.720 13.610 996.610 ;
        RECT 14.450 995.720 18.670 996.610 ;
        RECT 19.510 995.720 23.730 996.610 ;
        RECT 24.570 995.720 28.790 996.610 ;
        RECT 29.630 995.720 33.850 996.610 ;
        RECT 34.690 995.720 38.910 996.610 ;
        RECT 39.750 995.720 43.970 996.610 ;
        RECT 44.810 995.720 49.030 996.610 ;
        RECT 49.870 995.720 54.090 996.610 ;
        RECT 54.930 995.720 59.150 996.610 ;
        RECT 59.990 995.720 64.210 996.610 ;
        RECT 65.050 995.720 69.270 996.610 ;
        RECT 70.110 995.720 74.330 996.610 ;
        RECT 75.170 995.720 79.390 996.610 ;
        RECT 80.230 995.720 84.450 996.610 ;
        RECT 85.290 995.720 89.510 996.610 ;
        RECT 90.350 995.720 94.570 996.610 ;
        RECT 95.410 995.720 99.630 996.610 ;
        RECT 100.470 995.720 104.690 996.610 ;
        RECT 105.530 995.720 109.750 996.610 ;
        RECT 110.590 995.720 114.810 996.610 ;
        RECT 115.650 995.720 119.870 996.610 ;
        RECT 120.710 995.720 124.930 996.610 ;
        RECT 125.770 995.720 129.990 996.610 ;
        RECT 130.830 995.720 135.050 996.610 ;
        RECT 135.890 995.720 140.110 996.610 ;
        RECT 140.950 995.720 145.170 996.610 ;
        RECT 146.010 995.720 150.230 996.610 ;
        RECT 151.070 995.720 155.290 996.610 ;
        RECT 156.130 995.720 160.350 996.610 ;
        RECT 161.190 995.720 165.410 996.610 ;
        RECT 166.250 995.720 170.470 996.610 ;
        RECT 171.310 995.720 175.530 996.610 ;
        RECT 176.370 995.720 180.590 996.610 ;
        RECT 181.430 995.720 185.650 996.610 ;
        RECT 186.490 995.720 190.710 996.610 ;
        RECT 191.550 995.720 195.770 996.610 ;
        RECT 196.610 995.720 199.940 996.610 ;
        RECT 0.100 4.280 199.940 995.720 ;
        RECT 0.100 4.000 6.710 4.280 ;
        RECT 7.550 4.000 12.690 4.280 ;
        RECT 13.530 4.000 18.670 4.280 ;
        RECT 19.510 4.000 24.650 4.280 ;
        RECT 25.490 4.000 30.630 4.280 ;
        RECT 31.470 4.000 36.610 4.280 ;
        RECT 37.450 4.000 42.590 4.280 ;
        RECT 43.430 4.000 48.570 4.280 ;
        RECT 49.410 4.000 54.550 4.280 ;
        RECT 55.390 4.000 60.530 4.280 ;
        RECT 61.370 4.000 66.510 4.280 ;
        RECT 67.350 4.000 72.490 4.280 ;
        RECT 73.330 4.000 78.470 4.280 ;
        RECT 79.310 4.000 84.450 4.280 ;
        RECT 85.290 4.000 90.430 4.280 ;
        RECT 91.270 4.000 96.410 4.280 ;
        RECT 97.250 4.000 102.390 4.280 ;
        RECT 103.230 4.000 108.370 4.280 ;
        RECT 109.210 4.000 114.350 4.280 ;
        RECT 115.190 4.000 120.330 4.280 ;
        RECT 121.170 4.000 126.310 4.280 ;
        RECT 127.150 4.000 132.290 4.280 ;
        RECT 133.130 4.000 138.270 4.280 ;
        RECT 139.110 4.000 144.250 4.280 ;
        RECT 145.090 4.000 150.230 4.280 ;
        RECT 151.070 4.000 156.210 4.280 ;
        RECT 157.050 4.000 162.190 4.280 ;
        RECT 163.030 4.000 168.170 4.280 ;
        RECT 169.010 4.000 174.150 4.280 ;
        RECT 174.990 4.000 180.130 4.280 ;
        RECT 180.970 4.000 186.110 4.280 ;
        RECT 186.950 4.000 192.090 4.280 ;
        RECT 192.930 4.000 199.940 4.280 ;
      LAYER met3 ;
        RECT 1.905 991.080 195.600 991.945 ;
        RECT 1.905 985.680 196.000 991.080 ;
        RECT 1.905 984.280 195.600 985.680 ;
        RECT 1.905 978.880 196.000 984.280 ;
        RECT 1.905 977.480 195.600 978.880 ;
        RECT 1.905 972.080 196.000 977.480 ;
        RECT 1.905 970.680 195.600 972.080 ;
        RECT 1.905 965.280 196.000 970.680 ;
        RECT 1.905 963.880 195.600 965.280 ;
        RECT 1.905 958.480 196.000 963.880 ;
        RECT 1.905 957.080 195.600 958.480 ;
        RECT 1.905 951.680 196.000 957.080 ;
        RECT 1.905 950.280 195.600 951.680 ;
        RECT 1.905 944.880 196.000 950.280 ;
        RECT 1.905 943.480 195.600 944.880 ;
        RECT 1.905 938.080 196.000 943.480 ;
        RECT 1.905 936.680 195.600 938.080 ;
        RECT 1.905 931.280 196.000 936.680 ;
        RECT 1.905 929.880 195.600 931.280 ;
        RECT 1.905 924.480 196.000 929.880 ;
        RECT 1.905 923.080 195.600 924.480 ;
        RECT 1.905 917.680 196.000 923.080 ;
        RECT 1.905 916.280 195.600 917.680 ;
        RECT 1.905 910.880 196.000 916.280 ;
        RECT 1.905 909.480 195.600 910.880 ;
        RECT 1.905 904.080 196.000 909.480 ;
        RECT 1.905 902.680 195.600 904.080 ;
        RECT 1.905 897.280 196.000 902.680 ;
        RECT 1.905 895.880 195.600 897.280 ;
        RECT 1.905 890.480 196.000 895.880 ;
        RECT 1.905 889.080 195.600 890.480 ;
        RECT 1.905 883.680 196.000 889.080 ;
        RECT 1.905 882.280 195.600 883.680 ;
        RECT 1.905 876.880 196.000 882.280 ;
        RECT 1.905 875.480 195.600 876.880 ;
        RECT 1.905 870.080 196.000 875.480 ;
        RECT 1.905 868.680 195.600 870.080 ;
        RECT 1.905 863.280 196.000 868.680 ;
        RECT 1.905 861.880 195.600 863.280 ;
        RECT 1.905 856.480 196.000 861.880 ;
        RECT 1.905 855.080 195.600 856.480 ;
        RECT 1.905 849.680 196.000 855.080 ;
        RECT 1.905 848.280 195.600 849.680 ;
        RECT 1.905 842.880 196.000 848.280 ;
        RECT 4.400 841.480 195.600 842.880 ;
        RECT 1.905 840.160 196.000 841.480 ;
        RECT 4.400 838.760 196.000 840.160 ;
        RECT 1.905 837.440 196.000 838.760 ;
        RECT 4.400 836.080 196.000 837.440 ;
        RECT 4.400 836.040 195.600 836.080 ;
        RECT 1.905 834.720 195.600 836.040 ;
        RECT 4.400 834.680 195.600 834.720 ;
        RECT 4.400 833.320 196.000 834.680 ;
        RECT 1.905 832.000 196.000 833.320 ;
        RECT 4.400 830.600 196.000 832.000 ;
        RECT 1.905 829.280 196.000 830.600 ;
        RECT 4.400 827.880 195.600 829.280 ;
        RECT 1.905 826.560 196.000 827.880 ;
        RECT 4.400 825.160 196.000 826.560 ;
        RECT 1.905 823.840 196.000 825.160 ;
        RECT 4.400 822.480 196.000 823.840 ;
        RECT 4.400 822.440 195.600 822.480 ;
        RECT 1.905 821.120 195.600 822.440 ;
        RECT 4.400 821.080 195.600 821.120 ;
        RECT 4.400 819.720 196.000 821.080 ;
        RECT 1.905 818.400 196.000 819.720 ;
        RECT 4.400 817.000 196.000 818.400 ;
        RECT 1.905 815.680 196.000 817.000 ;
        RECT 4.400 814.280 195.600 815.680 ;
        RECT 1.905 812.960 196.000 814.280 ;
        RECT 4.400 811.560 196.000 812.960 ;
        RECT 1.905 810.240 196.000 811.560 ;
        RECT 4.400 808.880 196.000 810.240 ;
        RECT 4.400 808.840 195.600 808.880 ;
        RECT 1.905 807.520 195.600 808.840 ;
        RECT 4.400 807.480 195.600 807.520 ;
        RECT 4.400 806.120 196.000 807.480 ;
        RECT 1.905 804.800 196.000 806.120 ;
        RECT 4.400 803.400 196.000 804.800 ;
        RECT 1.905 802.080 196.000 803.400 ;
        RECT 4.400 800.680 195.600 802.080 ;
        RECT 1.905 799.360 196.000 800.680 ;
        RECT 4.400 797.960 196.000 799.360 ;
        RECT 1.905 796.640 196.000 797.960 ;
        RECT 4.400 795.280 196.000 796.640 ;
        RECT 4.400 795.240 195.600 795.280 ;
        RECT 1.905 793.920 195.600 795.240 ;
        RECT 4.400 793.880 195.600 793.920 ;
        RECT 4.400 792.520 196.000 793.880 ;
        RECT 1.905 791.200 196.000 792.520 ;
        RECT 4.400 789.800 196.000 791.200 ;
        RECT 1.905 788.480 196.000 789.800 ;
        RECT 4.400 787.080 195.600 788.480 ;
        RECT 1.905 785.760 196.000 787.080 ;
        RECT 4.400 784.360 196.000 785.760 ;
        RECT 1.905 783.040 196.000 784.360 ;
        RECT 4.400 781.680 196.000 783.040 ;
        RECT 4.400 781.640 195.600 781.680 ;
        RECT 1.905 780.320 195.600 781.640 ;
        RECT 4.400 780.280 195.600 780.320 ;
        RECT 4.400 778.920 196.000 780.280 ;
        RECT 1.905 777.600 196.000 778.920 ;
        RECT 4.400 776.200 196.000 777.600 ;
        RECT 1.905 774.880 196.000 776.200 ;
        RECT 4.400 773.480 195.600 774.880 ;
        RECT 1.905 772.160 196.000 773.480 ;
        RECT 4.400 770.760 196.000 772.160 ;
        RECT 1.905 769.440 196.000 770.760 ;
        RECT 4.400 768.080 196.000 769.440 ;
        RECT 4.400 768.040 195.600 768.080 ;
        RECT 1.905 766.720 195.600 768.040 ;
        RECT 4.400 766.680 195.600 766.720 ;
        RECT 4.400 765.320 196.000 766.680 ;
        RECT 1.905 764.000 196.000 765.320 ;
        RECT 4.400 762.600 196.000 764.000 ;
        RECT 1.905 761.280 196.000 762.600 ;
        RECT 4.400 759.880 195.600 761.280 ;
        RECT 1.905 758.560 196.000 759.880 ;
        RECT 4.400 757.160 196.000 758.560 ;
        RECT 1.905 755.840 196.000 757.160 ;
        RECT 4.400 754.480 196.000 755.840 ;
        RECT 4.400 754.440 195.600 754.480 ;
        RECT 1.905 753.120 195.600 754.440 ;
        RECT 4.400 753.080 195.600 753.120 ;
        RECT 4.400 751.720 196.000 753.080 ;
        RECT 1.905 750.400 196.000 751.720 ;
        RECT 4.400 749.000 196.000 750.400 ;
        RECT 1.905 747.680 196.000 749.000 ;
        RECT 4.400 746.280 195.600 747.680 ;
        RECT 1.905 744.960 196.000 746.280 ;
        RECT 4.400 743.560 196.000 744.960 ;
        RECT 1.905 742.240 196.000 743.560 ;
        RECT 4.400 740.880 196.000 742.240 ;
        RECT 4.400 740.840 195.600 740.880 ;
        RECT 1.905 739.520 195.600 740.840 ;
        RECT 4.400 739.480 195.600 739.520 ;
        RECT 4.400 738.120 196.000 739.480 ;
        RECT 1.905 736.800 196.000 738.120 ;
        RECT 4.400 735.400 196.000 736.800 ;
        RECT 1.905 734.080 196.000 735.400 ;
        RECT 4.400 732.680 195.600 734.080 ;
        RECT 1.905 731.360 196.000 732.680 ;
        RECT 4.400 729.960 196.000 731.360 ;
        RECT 1.905 728.640 196.000 729.960 ;
        RECT 4.400 727.280 196.000 728.640 ;
        RECT 4.400 727.240 195.600 727.280 ;
        RECT 1.905 725.920 195.600 727.240 ;
        RECT 4.400 725.880 195.600 725.920 ;
        RECT 4.400 724.520 196.000 725.880 ;
        RECT 1.905 723.200 196.000 724.520 ;
        RECT 4.400 721.800 196.000 723.200 ;
        RECT 1.905 720.480 196.000 721.800 ;
        RECT 4.400 719.080 195.600 720.480 ;
        RECT 1.905 717.760 196.000 719.080 ;
        RECT 4.400 716.360 196.000 717.760 ;
        RECT 1.905 715.040 196.000 716.360 ;
        RECT 4.400 713.680 196.000 715.040 ;
        RECT 4.400 713.640 195.600 713.680 ;
        RECT 1.905 712.320 195.600 713.640 ;
        RECT 4.400 712.280 195.600 712.320 ;
        RECT 4.400 710.920 196.000 712.280 ;
        RECT 1.905 709.600 196.000 710.920 ;
        RECT 4.400 708.200 196.000 709.600 ;
        RECT 1.905 706.880 196.000 708.200 ;
        RECT 4.400 705.480 195.600 706.880 ;
        RECT 1.905 704.160 196.000 705.480 ;
        RECT 4.400 702.760 196.000 704.160 ;
        RECT 1.905 701.440 196.000 702.760 ;
        RECT 4.400 700.080 196.000 701.440 ;
        RECT 4.400 700.040 195.600 700.080 ;
        RECT 1.905 698.720 195.600 700.040 ;
        RECT 4.400 698.680 195.600 698.720 ;
        RECT 4.400 697.320 196.000 698.680 ;
        RECT 1.905 696.000 196.000 697.320 ;
        RECT 4.400 694.600 196.000 696.000 ;
        RECT 1.905 693.280 196.000 694.600 ;
        RECT 4.400 691.880 195.600 693.280 ;
        RECT 1.905 690.560 196.000 691.880 ;
        RECT 4.400 689.160 196.000 690.560 ;
        RECT 1.905 687.840 196.000 689.160 ;
        RECT 4.400 686.480 196.000 687.840 ;
        RECT 4.400 686.440 195.600 686.480 ;
        RECT 1.905 685.120 195.600 686.440 ;
        RECT 4.400 685.080 195.600 685.120 ;
        RECT 4.400 683.720 196.000 685.080 ;
        RECT 1.905 682.400 196.000 683.720 ;
        RECT 4.400 681.000 196.000 682.400 ;
        RECT 1.905 679.680 196.000 681.000 ;
        RECT 4.400 678.280 195.600 679.680 ;
        RECT 1.905 676.960 196.000 678.280 ;
        RECT 4.400 675.560 196.000 676.960 ;
        RECT 1.905 674.240 196.000 675.560 ;
        RECT 4.400 672.880 196.000 674.240 ;
        RECT 4.400 672.840 195.600 672.880 ;
        RECT 1.905 671.520 195.600 672.840 ;
        RECT 4.400 671.480 195.600 671.520 ;
        RECT 4.400 670.120 196.000 671.480 ;
        RECT 1.905 668.800 196.000 670.120 ;
        RECT 4.400 667.400 196.000 668.800 ;
        RECT 1.905 666.080 196.000 667.400 ;
        RECT 4.400 664.680 195.600 666.080 ;
        RECT 1.905 663.360 196.000 664.680 ;
        RECT 4.400 661.960 196.000 663.360 ;
        RECT 1.905 660.640 196.000 661.960 ;
        RECT 4.400 659.280 196.000 660.640 ;
        RECT 4.400 659.240 195.600 659.280 ;
        RECT 1.905 657.920 195.600 659.240 ;
        RECT 4.400 657.880 195.600 657.920 ;
        RECT 4.400 656.520 196.000 657.880 ;
        RECT 1.905 655.200 196.000 656.520 ;
        RECT 4.400 653.800 196.000 655.200 ;
        RECT 1.905 652.480 196.000 653.800 ;
        RECT 4.400 651.080 195.600 652.480 ;
        RECT 1.905 649.760 196.000 651.080 ;
        RECT 4.400 648.360 196.000 649.760 ;
        RECT 1.905 647.040 196.000 648.360 ;
        RECT 4.400 645.680 196.000 647.040 ;
        RECT 4.400 645.640 195.600 645.680 ;
        RECT 1.905 644.320 195.600 645.640 ;
        RECT 4.400 644.280 195.600 644.320 ;
        RECT 4.400 642.920 196.000 644.280 ;
        RECT 1.905 641.600 196.000 642.920 ;
        RECT 4.400 640.200 196.000 641.600 ;
        RECT 1.905 638.880 196.000 640.200 ;
        RECT 4.400 637.480 195.600 638.880 ;
        RECT 1.905 636.160 196.000 637.480 ;
        RECT 4.400 634.760 196.000 636.160 ;
        RECT 1.905 633.440 196.000 634.760 ;
        RECT 4.400 632.080 196.000 633.440 ;
        RECT 4.400 632.040 195.600 632.080 ;
        RECT 1.905 630.720 195.600 632.040 ;
        RECT 4.400 630.680 195.600 630.720 ;
        RECT 4.400 629.320 196.000 630.680 ;
        RECT 1.905 628.000 196.000 629.320 ;
        RECT 4.400 626.600 196.000 628.000 ;
        RECT 1.905 625.280 196.000 626.600 ;
        RECT 4.400 623.880 195.600 625.280 ;
        RECT 1.905 622.560 196.000 623.880 ;
        RECT 4.400 621.160 196.000 622.560 ;
        RECT 1.905 619.840 196.000 621.160 ;
        RECT 4.400 618.480 196.000 619.840 ;
        RECT 4.400 618.440 195.600 618.480 ;
        RECT 1.905 617.120 195.600 618.440 ;
        RECT 4.400 617.080 195.600 617.120 ;
        RECT 4.400 615.720 196.000 617.080 ;
        RECT 1.905 614.400 196.000 615.720 ;
        RECT 4.400 613.000 196.000 614.400 ;
        RECT 1.905 611.680 196.000 613.000 ;
        RECT 4.400 610.280 195.600 611.680 ;
        RECT 1.905 608.960 196.000 610.280 ;
        RECT 4.400 607.560 196.000 608.960 ;
        RECT 1.905 606.240 196.000 607.560 ;
        RECT 4.400 604.880 196.000 606.240 ;
        RECT 4.400 604.840 195.600 604.880 ;
        RECT 1.905 603.520 195.600 604.840 ;
        RECT 4.400 603.480 195.600 603.520 ;
        RECT 4.400 602.120 196.000 603.480 ;
        RECT 1.905 600.800 196.000 602.120 ;
        RECT 4.400 599.400 196.000 600.800 ;
        RECT 1.905 598.080 196.000 599.400 ;
        RECT 4.400 596.680 195.600 598.080 ;
        RECT 1.905 595.360 196.000 596.680 ;
        RECT 4.400 593.960 196.000 595.360 ;
        RECT 1.905 592.640 196.000 593.960 ;
        RECT 4.400 591.280 196.000 592.640 ;
        RECT 4.400 591.240 195.600 591.280 ;
        RECT 1.905 589.920 195.600 591.240 ;
        RECT 4.400 589.880 195.600 589.920 ;
        RECT 4.400 588.520 196.000 589.880 ;
        RECT 1.905 587.200 196.000 588.520 ;
        RECT 4.400 585.800 196.000 587.200 ;
        RECT 1.905 584.480 196.000 585.800 ;
        RECT 4.400 583.080 195.600 584.480 ;
        RECT 1.905 581.760 196.000 583.080 ;
        RECT 4.400 580.360 196.000 581.760 ;
        RECT 1.905 579.040 196.000 580.360 ;
        RECT 4.400 577.680 196.000 579.040 ;
        RECT 4.400 577.640 195.600 577.680 ;
        RECT 1.905 576.320 195.600 577.640 ;
        RECT 4.400 576.280 195.600 576.320 ;
        RECT 4.400 574.920 196.000 576.280 ;
        RECT 1.905 573.600 196.000 574.920 ;
        RECT 4.400 572.200 196.000 573.600 ;
        RECT 1.905 570.880 196.000 572.200 ;
        RECT 4.400 569.480 195.600 570.880 ;
        RECT 1.905 568.160 196.000 569.480 ;
        RECT 4.400 566.760 196.000 568.160 ;
        RECT 1.905 565.440 196.000 566.760 ;
        RECT 4.400 564.080 196.000 565.440 ;
        RECT 4.400 564.040 195.600 564.080 ;
        RECT 1.905 562.720 195.600 564.040 ;
        RECT 4.400 562.680 195.600 562.720 ;
        RECT 4.400 561.320 196.000 562.680 ;
        RECT 1.905 560.000 196.000 561.320 ;
        RECT 4.400 558.600 196.000 560.000 ;
        RECT 1.905 557.280 196.000 558.600 ;
        RECT 4.400 555.880 195.600 557.280 ;
        RECT 1.905 554.560 196.000 555.880 ;
        RECT 4.400 553.160 196.000 554.560 ;
        RECT 1.905 551.840 196.000 553.160 ;
        RECT 4.400 550.480 196.000 551.840 ;
        RECT 4.400 550.440 195.600 550.480 ;
        RECT 1.905 549.120 195.600 550.440 ;
        RECT 4.400 549.080 195.600 549.120 ;
        RECT 4.400 547.720 196.000 549.080 ;
        RECT 1.905 546.400 196.000 547.720 ;
        RECT 4.400 545.000 196.000 546.400 ;
        RECT 1.905 543.680 196.000 545.000 ;
        RECT 4.400 542.280 195.600 543.680 ;
        RECT 1.905 540.960 196.000 542.280 ;
        RECT 4.400 539.560 196.000 540.960 ;
        RECT 1.905 538.240 196.000 539.560 ;
        RECT 4.400 536.880 196.000 538.240 ;
        RECT 4.400 536.840 195.600 536.880 ;
        RECT 1.905 535.520 195.600 536.840 ;
        RECT 4.400 535.480 195.600 535.520 ;
        RECT 4.400 534.120 196.000 535.480 ;
        RECT 1.905 532.800 196.000 534.120 ;
        RECT 4.400 531.400 196.000 532.800 ;
        RECT 1.905 530.080 196.000 531.400 ;
        RECT 4.400 528.680 195.600 530.080 ;
        RECT 1.905 527.360 196.000 528.680 ;
        RECT 4.400 525.960 196.000 527.360 ;
        RECT 1.905 524.640 196.000 525.960 ;
        RECT 4.400 523.280 196.000 524.640 ;
        RECT 4.400 523.240 195.600 523.280 ;
        RECT 1.905 521.920 195.600 523.240 ;
        RECT 4.400 521.880 195.600 521.920 ;
        RECT 4.400 520.520 196.000 521.880 ;
        RECT 1.905 519.200 196.000 520.520 ;
        RECT 4.400 517.800 196.000 519.200 ;
        RECT 1.905 516.480 196.000 517.800 ;
        RECT 4.400 515.080 195.600 516.480 ;
        RECT 1.905 513.760 196.000 515.080 ;
        RECT 4.400 512.360 196.000 513.760 ;
        RECT 1.905 511.040 196.000 512.360 ;
        RECT 4.400 509.680 196.000 511.040 ;
        RECT 4.400 509.640 195.600 509.680 ;
        RECT 1.905 508.320 195.600 509.640 ;
        RECT 4.400 508.280 195.600 508.320 ;
        RECT 4.400 506.920 196.000 508.280 ;
        RECT 1.905 505.600 196.000 506.920 ;
        RECT 4.400 504.200 196.000 505.600 ;
        RECT 1.905 502.880 196.000 504.200 ;
        RECT 4.400 501.480 195.600 502.880 ;
        RECT 1.905 500.160 196.000 501.480 ;
        RECT 4.400 498.760 196.000 500.160 ;
        RECT 1.905 497.440 196.000 498.760 ;
        RECT 4.400 496.080 196.000 497.440 ;
        RECT 4.400 496.040 195.600 496.080 ;
        RECT 1.905 494.720 195.600 496.040 ;
        RECT 4.400 494.680 195.600 494.720 ;
        RECT 4.400 493.320 196.000 494.680 ;
        RECT 1.905 492.000 196.000 493.320 ;
        RECT 4.400 490.600 196.000 492.000 ;
        RECT 1.905 489.280 196.000 490.600 ;
        RECT 4.400 487.880 195.600 489.280 ;
        RECT 1.905 486.560 196.000 487.880 ;
        RECT 4.400 485.160 196.000 486.560 ;
        RECT 1.905 483.840 196.000 485.160 ;
        RECT 4.400 482.480 196.000 483.840 ;
        RECT 4.400 482.440 195.600 482.480 ;
        RECT 1.905 481.120 195.600 482.440 ;
        RECT 4.400 481.080 195.600 481.120 ;
        RECT 4.400 479.720 196.000 481.080 ;
        RECT 1.905 478.400 196.000 479.720 ;
        RECT 4.400 477.000 196.000 478.400 ;
        RECT 1.905 475.680 196.000 477.000 ;
        RECT 4.400 474.280 195.600 475.680 ;
        RECT 1.905 472.960 196.000 474.280 ;
        RECT 4.400 471.560 196.000 472.960 ;
        RECT 1.905 470.240 196.000 471.560 ;
        RECT 4.400 468.880 196.000 470.240 ;
        RECT 4.400 468.840 195.600 468.880 ;
        RECT 1.905 467.520 195.600 468.840 ;
        RECT 4.400 467.480 195.600 467.520 ;
        RECT 4.400 466.120 196.000 467.480 ;
        RECT 1.905 464.800 196.000 466.120 ;
        RECT 4.400 463.400 196.000 464.800 ;
        RECT 1.905 462.080 196.000 463.400 ;
        RECT 4.400 460.680 195.600 462.080 ;
        RECT 1.905 459.360 196.000 460.680 ;
        RECT 4.400 457.960 196.000 459.360 ;
        RECT 1.905 456.640 196.000 457.960 ;
        RECT 4.400 455.280 196.000 456.640 ;
        RECT 4.400 455.240 195.600 455.280 ;
        RECT 1.905 453.920 195.600 455.240 ;
        RECT 4.400 453.880 195.600 453.920 ;
        RECT 4.400 452.520 196.000 453.880 ;
        RECT 1.905 451.200 196.000 452.520 ;
        RECT 4.400 449.800 196.000 451.200 ;
        RECT 1.905 448.480 196.000 449.800 ;
        RECT 4.400 447.080 195.600 448.480 ;
        RECT 1.905 445.760 196.000 447.080 ;
        RECT 4.400 444.360 196.000 445.760 ;
        RECT 1.905 443.040 196.000 444.360 ;
        RECT 4.400 441.680 196.000 443.040 ;
        RECT 4.400 441.640 195.600 441.680 ;
        RECT 1.905 440.320 195.600 441.640 ;
        RECT 4.400 440.280 195.600 440.320 ;
        RECT 4.400 438.920 196.000 440.280 ;
        RECT 1.905 437.600 196.000 438.920 ;
        RECT 4.400 436.200 196.000 437.600 ;
        RECT 1.905 434.880 196.000 436.200 ;
        RECT 4.400 433.480 195.600 434.880 ;
        RECT 1.905 432.160 196.000 433.480 ;
        RECT 4.400 430.760 196.000 432.160 ;
        RECT 1.905 429.440 196.000 430.760 ;
        RECT 4.400 428.080 196.000 429.440 ;
        RECT 4.400 428.040 195.600 428.080 ;
        RECT 1.905 426.720 195.600 428.040 ;
        RECT 4.400 426.680 195.600 426.720 ;
        RECT 4.400 425.320 196.000 426.680 ;
        RECT 1.905 424.000 196.000 425.320 ;
        RECT 4.400 422.600 196.000 424.000 ;
        RECT 1.905 421.280 196.000 422.600 ;
        RECT 4.400 419.880 195.600 421.280 ;
        RECT 1.905 418.560 196.000 419.880 ;
        RECT 4.400 417.160 196.000 418.560 ;
        RECT 1.905 415.840 196.000 417.160 ;
        RECT 4.400 414.480 196.000 415.840 ;
        RECT 4.400 414.440 195.600 414.480 ;
        RECT 1.905 413.120 195.600 414.440 ;
        RECT 4.400 413.080 195.600 413.120 ;
        RECT 4.400 411.720 196.000 413.080 ;
        RECT 1.905 410.400 196.000 411.720 ;
        RECT 4.400 409.000 196.000 410.400 ;
        RECT 1.905 407.680 196.000 409.000 ;
        RECT 4.400 406.280 195.600 407.680 ;
        RECT 1.905 404.960 196.000 406.280 ;
        RECT 4.400 403.560 196.000 404.960 ;
        RECT 1.905 402.240 196.000 403.560 ;
        RECT 4.400 400.880 196.000 402.240 ;
        RECT 4.400 400.840 195.600 400.880 ;
        RECT 1.905 399.520 195.600 400.840 ;
        RECT 4.400 399.480 195.600 399.520 ;
        RECT 4.400 398.120 196.000 399.480 ;
        RECT 1.905 396.800 196.000 398.120 ;
        RECT 4.400 395.400 196.000 396.800 ;
        RECT 1.905 394.080 196.000 395.400 ;
        RECT 4.400 392.680 195.600 394.080 ;
        RECT 1.905 391.360 196.000 392.680 ;
        RECT 4.400 389.960 196.000 391.360 ;
        RECT 1.905 388.640 196.000 389.960 ;
        RECT 4.400 387.280 196.000 388.640 ;
        RECT 4.400 387.240 195.600 387.280 ;
        RECT 1.905 385.920 195.600 387.240 ;
        RECT 4.400 385.880 195.600 385.920 ;
        RECT 4.400 384.520 196.000 385.880 ;
        RECT 1.905 383.200 196.000 384.520 ;
        RECT 4.400 381.800 196.000 383.200 ;
        RECT 1.905 380.480 196.000 381.800 ;
        RECT 4.400 379.080 195.600 380.480 ;
        RECT 1.905 377.760 196.000 379.080 ;
        RECT 4.400 376.360 196.000 377.760 ;
        RECT 1.905 375.040 196.000 376.360 ;
        RECT 4.400 373.680 196.000 375.040 ;
        RECT 4.400 373.640 195.600 373.680 ;
        RECT 1.905 372.320 195.600 373.640 ;
        RECT 4.400 372.280 195.600 372.320 ;
        RECT 4.400 370.920 196.000 372.280 ;
        RECT 1.905 369.600 196.000 370.920 ;
        RECT 4.400 368.200 196.000 369.600 ;
        RECT 1.905 366.880 196.000 368.200 ;
        RECT 4.400 365.480 195.600 366.880 ;
        RECT 1.905 364.160 196.000 365.480 ;
        RECT 4.400 362.760 196.000 364.160 ;
        RECT 1.905 361.440 196.000 362.760 ;
        RECT 4.400 360.080 196.000 361.440 ;
        RECT 4.400 360.040 195.600 360.080 ;
        RECT 1.905 358.720 195.600 360.040 ;
        RECT 4.400 358.680 195.600 358.720 ;
        RECT 4.400 357.320 196.000 358.680 ;
        RECT 1.905 356.000 196.000 357.320 ;
        RECT 4.400 354.600 196.000 356.000 ;
        RECT 1.905 353.280 196.000 354.600 ;
        RECT 4.400 351.880 195.600 353.280 ;
        RECT 1.905 350.560 196.000 351.880 ;
        RECT 4.400 349.160 196.000 350.560 ;
        RECT 1.905 347.840 196.000 349.160 ;
        RECT 4.400 346.480 196.000 347.840 ;
        RECT 4.400 346.440 195.600 346.480 ;
        RECT 1.905 345.120 195.600 346.440 ;
        RECT 4.400 345.080 195.600 345.120 ;
        RECT 4.400 343.720 196.000 345.080 ;
        RECT 1.905 342.400 196.000 343.720 ;
        RECT 4.400 341.000 196.000 342.400 ;
        RECT 1.905 339.680 196.000 341.000 ;
        RECT 4.400 338.280 195.600 339.680 ;
        RECT 1.905 336.960 196.000 338.280 ;
        RECT 4.400 335.560 196.000 336.960 ;
        RECT 1.905 334.240 196.000 335.560 ;
        RECT 4.400 332.880 196.000 334.240 ;
        RECT 4.400 332.840 195.600 332.880 ;
        RECT 1.905 331.520 195.600 332.840 ;
        RECT 4.400 331.480 195.600 331.520 ;
        RECT 4.400 330.120 196.000 331.480 ;
        RECT 1.905 328.800 196.000 330.120 ;
        RECT 4.400 327.400 196.000 328.800 ;
        RECT 1.905 326.080 196.000 327.400 ;
        RECT 4.400 324.680 195.600 326.080 ;
        RECT 1.905 323.360 196.000 324.680 ;
        RECT 4.400 321.960 196.000 323.360 ;
        RECT 1.905 320.640 196.000 321.960 ;
        RECT 4.400 319.280 196.000 320.640 ;
        RECT 4.400 319.240 195.600 319.280 ;
        RECT 1.905 317.920 195.600 319.240 ;
        RECT 4.400 317.880 195.600 317.920 ;
        RECT 4.400 316.520 196.000 317.880 ;
        RECT 1.905 315.200 196.000 316.520 ;
        RECT 4.400 313.800 196.000 315.200 ;
        RECT 1.905 312.480 196.000 313.800 ;
        RECT 4.400 311.080 195.600 312.480 ;
        RECT 1.905 309.760 196.000 311.080 ;
        RECT 4.400 308.360 196.000 309.760 ;
        RECT 1.905 307.040 196.000 308.360 ;
        RECT 4.400 305.680 196.000 307.040 ;
        RECT 4.400 305.640 195.600 305.680 ;
        RECT 1.905 304.320 195.600 305.640 ;
        RECT 4.400 304.280 195.600 304.320 ;
        RECT 4.400 302.920 196.000 304.280 ;
        RECT 1.905 301.600 196.000 302.920 ;
        RECT 4.400 300.200 196.000 301.600 ;
        RECT 1.905 298.880 196.000 300.200 ;
        RECT 4.400 297.480 195.600 298.880 ;
        RECT 1.905 296.160 196.000 297.480 ;
        RECT 4.400 294.760 196.000 296.160 ;
        RECT 1.905 293.440 196.000 294.760 ;
        RECT 4.400 292.080 196.000 293.440 ;
        RECT 4.400 292.040 195.600 292.080 ;
        RECT 1.905 290.720 195.600 292.040 ;
        RECT 4.400 290.680 195.600 290.720 ;
        RECT 4.400 289.320 196.000 290.680 ;
        RECT 1.905 288.000 196.000 289.320 ;
        RECT 4.400 286.600 196.000 288.000 ;
        RECT 1.905 285.280 196.000 286.600 ;
        RECT 4.400 283.880 195.600 285.280 ;
        RECT 1.905 282.560 196.000 283.880 ;
        RECT 4.400 281.160 196.000 282.560 ;
        RECT 1.905 279.840 196.000 281.160 ;
        RECT 4.400 278.480 196.000 279.840 ;
        RECT 4.400 278.440 195.600 278.480 ;
        RECT 1.905 277.120 195.600 278.440 ;
        RECT 4.400 277.080 195.600 277.120 ;
        RECT 4.400 275.720 196.000 277.080 ;
        RECT 1.905 274.400 196.000 275.720 ;
        RECT 4.400 273.000 196.000 274.400 ;
        RECT 1.905 271.680 196.000 273.000 ;
        RECT 4.400 270.280 195.600 271.680 ;
        RECT 1.905 268.960 196.000 270.280 ;
        RECT 4.400 267.560 196.000 268.960 ;
        RECT 1.905 266.240 196.000 267.560 ;
        RECT 4.400 264.880 196.000 266.240 ;
        RECT 4.400 264.840 195.600 264.880 ;
        RECT 1.905 263.520 195.600 264.840 ;
        RECT 4.400 263.480 195.600 263.520 ;
        RECT 4.400 262.120 196.000 263.480 ;
        RECT 1.905 260.800 196.000 262.120 ;
        RECT 4.400 259.400 196.000 260.800 ;
        RECT 1.905 258.080 196.000 259.400 ;
        RECT 4.400 256.680 195.600 258.080 ;
        RECT 1.905 255.360 196.000 256.680 ;
        RECT 4.400 253.960 196.000 255.360 ;
        RECT 1.905 252.640 196.000 253.960 ;
        RECT 4.400 251.280 196.000 252.640 ;
        RECT 4.400 251.240 195.600 251.280 ;
        RECT 1.905 249.920 195.600 251.240 ;
        RECT 4.400 249.880 195.600 249.920 ;
        RECT 4.400 248.520 196.000 249.880 ;
        RECT 1.905 247.200 196.000 248.520 ;
        RECT 4.400 245.800 196.000 247.200 ;
        RECT 1.905 244.480 196.000 245.800 ;
        RECT 4.400 243.080 195.600 244.480 ;
        RECT 1.905 241.760 196.000 243.080 ;
        RECT 4.400 240.360 196.000 241.760 ;
        RECT 1.905 239.040 196.000 240.360 ;
        RECT 4.400 237.680 196.000 239.040 ;
        RECT 4.400 237.640 195.600 237.680 ;
        RECT 1.905 236.320 195.600 237.640 ;
        RECT 4.400 236.280 195.600 236.320 ;
        RECT 4.400 234.920 196.000 236.280 ;
        RECT 1.905 233.600 196.000 234.920 ;
        RECT 4.400 232.200 196.000 233.600 ;
        RECT 1.905 230.880 196.000 232.200 ;
        RECT 4.400 229.480 195.600 230.880 ;
        RECT 1.905 228.160 196.000 229.480 ;
        RECT 4.400 226.760 196.000 228.160 ;
        RECT 1.905 225.440 196.000 226.760 ;
        RECT 4.400 224.080 196.000 225.440 ;
        RECT 4.400 224.040 195.600 224.080 ;
        RECT 1.905 222.720 195.600 224.040 ;
        RECT 4.400 222.680 195.600 222.720 ;
        RECT 4.400 221.320 196.000 222.680 ;
        RECT 1.905 220.000 196.000 221.320 ;
        RECT 4.400 218.600 196.000 220.000 ;
        RECT 1.905 217.280 196.000 218.600 ;
        RECT 4.400 215.880 195.600 217.280 ;
        RECT 1.905 214.560 196.000 215.880 ;
        RECT 4.400 213.160 196.000 214.560 ;
        RECT 1.905 211.840 196.000 213.160 ;
        RECT 4.400 210.480 196.000 211.840 ;
        RECT 4.400 210.440 195.600 210.480 ;
        RECT 1.905 209.120 195.600 210.440 ;
        RECT 4.400 209.080 195.600 209.120 ;
        RECT 4.400 207.720 196.000 209.080 ;
        RECT 1.905 206.400 196.000 207.720 ;
        RECT 4.400 205.000 196.000 206.400 ;
        RECT 1.905 203.680 196.000 205.000 ;
        RECT 4.400 202.280 195.600 203.680 ;
        RECT 1.905 200.960 196.000 202.280 ;
        RECT 4.400 199.560 196.000 200.960 ;
        RECT 1.905 198.240 196.000 199.560 ;
        RECT 4.400 196.880 196.000 198.240 ;
        RECT 4.400 196.840 195.600 196.880 ;
        RECT 1.905 195.520 195.600 196.840 ;
        RECT 4.400 195.480 195.600 195.520 ;
        RECT 4.400 194.120 196.000 195.480 ;
        RECT 1.905 192.800 196.000 194.120 ;
        RECT 4.400 191.400 196.000 192.800 ;
        RECT 1.905 190.080 196.000 191.400 ;
        RECT 4.400 188.680 195.600 190.080 ;
        RECT 1.905 187.360 196.000 188.680 ;
        RECT 4.400 185.960 196.000 187.360 ;
        RECT 1.905 184.640 196.000 185.960 ;
        RECT 4.400 183.280 196.000 184.640 ;
        RECT 4.400 183.240 195.600 183.280 ;
        RECT 1.905 181.920 195.600 183.240 ;
        RECT 4.400 181.880 195.600 181.920 ;
        RECT 4.400 180.520 196.000 181.880 ;
        RECT 1.905 179.200 196.000 180.520 ;
        RECT 4.400 177.800 196.000 179.200 ;
        RECT 1.905 176.480 196.000 177.800 ;
        RECT 4.400 175.080 195.600 176.480 ;
        RECT 1.905 173.760 196.000 175.080 ;
        RECT 4.400 172.360 196.000 173.760 ;
        RECT 1.905 171.040 196.000 172.360 ;
        RECT 4.400 169.680 196.000 171.040 ;
        RECT 4.400 169.640 195.600 169.680 ;
        RECT 1.905 168.320 195.600 169.640 ;
        RECT 4.400 168.280 195.600 168.320 ;
        RECT 4.400 166.920 196.000 168.280 ;
        RECT 1.905 165.600 196.000 166.920 ;
        RECT 4.400 164.200 196.000 165.600 ;
        RECT 1.905 162.880 196.000 164.200 ;
        RECT 4.400 161.480 195.600 162.880 ;
        RECT 1.905 160.160 196.000 161.480 ;
        RECT 4.400 158.760 196.000 160.160 ;
        RECT 1.905 157.440 196.000 158.760 ;
        RECT 4.400 156.080 196.000 157.440 ;
        RECT 4.400 156.040 195.600 156.080 ;
        RECT 1.905 154.680 195.600 156.040 ;
        RECT 1.905 149.280 196.000 154.680 ;
        RECT 1.905 147.880 195.600 149.280 ;
        RECT 1.905 142.480 196.000 147.880 ;
        RECT 1.905 141.080 195.600 142.480 ;
        RECT 1.905 135.680 196.000 141.080 ;
        RECT 1.905 134.280 195.600 135.680 ;
        RECT 1.905 128.880 196.000 134.280 ;
        RECT 1.905 127.480 195.600 128.880 ;
        RECT 1.905 122.080 196.000 127.480 ;
        RECT 1.905 120.680 195.600 122.080 ;
        RECT 1.905 115.280 196.000 120.680 ;
        RECT 1.905 113.880 195.600 115.280 ;
        RECT 1.905 108.480 196.000 113.880 ;
        RECT 1.905 107.080 195.600 108.480 ;
        RECT 1.905 101.680 196.000 107.080 ;
        RECT 1.905 100.280 195.600 101.680 ;
        RECT 1.905 94.880 196.000 100.280 ;
        RECT 1.905 93.480 195.600 94.880 ;
        RECT 1.905 88.080 196.000 93.480 ;
        RECT 1.905 86.680 195.600 88.080 ;
        RECT 1.905 81.280 196.000 86.680 ;
        RECT 1.905 79.880 195.600 81.280 ;
        RECT 1.905 74.480 196.000 79.880 ;
        RECT 1.905 73.080 195.600 74.480 ;
        RECT 1.905 67.680 196.000 73.080 ;
        RECT 1.905 66.280 195.600 67.680 ;
        RECT 1.905 60.880 196.000 66.280 ;
        RECT 1.905 59.480 195.600 60.880 ;
        RECT 1.905 54.080 196.000 59.480 ;
        RECT 1.905 52.680 195.600 54.080 ;
        RECT 1.905 47.280 196.000 52.680 ;
        RECT 1.905 45.880 195.600 47.280 ;
        RECT 1.905 40.480 196.000 45.880 ;
        RECT 1.905 39.080 195.600 40.480 ;
        RECT 1.905 33.680 196.000 39.080 ;
        RECT 1.905 32.280 195.600 33.680 ;
        RECT 1.905 26.880 196.000 32.280 ;
        RECT 1.905 25.480 195.600 26.880 ;
        RECT 1.905 20.080 196.000 25.480 ;
        RECT 1.905 18.680 195.600 20.080 ;
        RECT 1.905 13.280 196.000 18.680 ;
        RECT 1.905 11.880 195.600 13.280 ;
        RECT 1.905 6.480 196.000 11.880 ;
        RECT 1.905 5.615 195.600 6.480 ;
      LAYER met4 ;
        RECT 3.055 17.175 20.640 800.865 ;
        RECT 23.040 17.175 97.440 800.865 ;
        RECT 99.840 17.175 174.240 800.865 ;
        RECT 176.640 17.175 185.545 800.865 ;
  END
END multiplexer
END LIBRARY

