magic
tech sky130B
magscale 1 2
timestamp 1717368054
<< metal1 >>
rect 300118 700340 300124 700392
rect 300176 700380 300182 700392
rect 322198 700380 322204 700392
rect 300176 700352 322204 700380
rect 300176 700340 300182 700352
rect 322198 700340 322204 700352
rect 322256 700340 322262 700392
rect 527174 700340 527180 700392
rect 527232 700380 527238 700392
rect 543918 700380 543924 700392
rect 527232 700352 543924 700380
rect 527232 700340 527238 700352
rect 543918 700340 543924 700352
rect 543976 700340 543982 700392
rect 170306 700272 170312 700324
rect 170364 700312 170370 700324
rect 324958 700312 324964 700324
rect 170364 700284 324964 700312
rect 170364 700272 170370 700284
rect 324958 700272 324964 700284
rect 325016 700272 325022 700324
rect 332502 700272 332508 700324
rect 332560 700312 332566 700324
rect 340138 700312 340144 700324
rect 332560 700284 340144 700312
rect 332560 700272 332566 700284
rect 340138 700272 340144 700284
rect 340196 700272 340202 700324
rect 509142 700272 509148 700324
rect 509200 700312 509206 700324
rect 559650 700312 559656 700324
rect 509200 700284 559656 700312
rect 509200 700272 509206 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 40494 699660 40500 699712
rect 40552 699700 40558 699712
rect 41414 699700 41420 699712
rect 40552 699672 41420 699700
rect 40552 699660 40558 699672
rect 41414 699660 41420 699672
rect 41472 699700 41478 699712
rect 86218 699700 86224 699712
rect 41472 699672 86224 699700
rect 41472 699660 41478 699672
rect 86218 699660 86224 699672
rect 86276 699660 86282 699712
rect 478506 699660 478512 699712
rect 478564 699700 478570 699712
rect 479518 699700 479524 699712
rect 478564 699672 479524 699700
rect 478564 699660 478570 699672
rect 479518 699660 479524 699672
rect 479576 699660 479582 699712
rect 255958 687896 255964 687948
rect 256016 687936 256022 687948
rect 267642 687936 267648 687948
rect 256016 687908 267648 687936
rect 256016 687896 256022 687908
rect 267642 687896 267648 687908
rect 267700 687896 267706 687948
rect 283834 687148 283840 687200
rect 283892 687188 283898 687200
rect 286318 687188 286324 687200
rect 283892 687160 286324 687188
rect 283892 687148 283898 687160
rect 286318 687148 286324 687160
rect 286376 687148 286382 687200
rect 348786 686468 348792 686520
rect 348844 686508 348850 686520
rect 358078 686508 358084 686520
rect 348844 686480 358084 686508
rect 348844 686468 348850 686480
rect 358078 686468 358084 686480
rect 358136 686468 358142 686520
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 26142 683176 26148 683188
rect 3476 683148 26148 683176
rect 3476 683136 3482 683148
rect 26142 683136 26148 683148
rect 26200 683176 26206 683188
rect 87598 683176 87604 683188
rect 26200 683148 87604 683176
rect 26200 683136 26206 683148
rect 87598 683136 87604 683148
rect 87656 683136 87662 683188
rect 358078 680348 358084 680400
rect 358136 680388 358142 680400
rect 360838 680388 360844 680400
rect 358136 680360 360844 680388
rect 358136 680348 358142 680360
rect 360838 680348 360844 680360
rect 360896 680348 360902 680400
rect 340138 677492 340144 677544
rect 340196 677532 340202 677544
rect 345658 677532 345664 677544
rect 340196 677504 345664 677532
rect 340196 677492 340202 677504
rect 345658 677492 345664 677504
rect 345716 677492 345722 677544
rect 250438 674772 250444 674824
rect 250496 674812 250502 674824
rect 255958 674812 255964 674824
rect 250496 674784 255964 674812
rect 250496 674772 250502 674784
rect 255958 674772 255964 674784
rect 256016 674772 256022 674824
rect 360838 672052 360844 672104
rect 360896 672092 360902 672104
rect 366358 672092 366364 672104
rect 360896 672064 366364 672092
rect 360896 672052 360902 672064
rect 366358 672052 366364 672064
rect 366416 672052 366422 672104
rect 242434 661716 242440 661768
rect 242492 661756 242498 661768
rect 250438 661756 250444 661768
rect 242492 661728 250444 661756
rect 242492 661716 242498 661728
rect 250438 661716 250444 661728
rect 250496 661716 250502 661768
rect 345658 660288 345664 660340
rect 345716 660328 345722 660340
rect 355962 660328 355968 660340
rect 345716 660300 355968 660328
rect 345716 660288 345722 660300
rect 355962 660288 355968 660300
rect 356020 660288 356026 660340
rect 45462 658248 45468 658300
rect 45520 658288 45526 658300
rect 105446 658288 105452 658300
rect 45520 658260 105452 658288
rect 45520 658248 45526 658260
rect 105446 658248 105452 658260
rect 105504 658288 105510 658300
rect 106182 658288 106188 658300
rect 105504 658260 106188 658288
rect 105504 658248 105510 658260
rect 106182 658248 106188 658260
rect 106240 658248 106246 658300
rect 489730 657976 489736 658028
rect 489788 658016 489794 658028
rect 501782 658016 501788 658028
rect 489788 657988 501788 658016
rect 489788 657976 489794 657988
rect 501782 657976 501788 657988
rect 501840 657976 501846 658028
rect 486970 657840 486976 657892
rect 487028 657880 487034 657892
rect 496262 657880 496268 657892
rect 487028 657852 496268 657880
rect 487028 657840 487034 657852
rect 496262 657840 496268 657852
rect 496320 657840 496326 657892
rect 364978 657772 364984 657824
rect 365036 657812 365042 657824
rect 491018 657812 491024 657824
rect 365036 657784 491024 657812
rect 365036 657772 365042 657784
rect 491018 657772 491024 657784
rect 491076 657772 491082 657824
rect 322198 657704 322204 657756
rect 322256 657744 322262 657756
rect 490466 657744 490472 657756
rect 322256 657716 490472 657744
rect 322256 657704 322262 657716
rect 490466 657704 490472 657716
rect 490524 657744 490530 657756
rect 491202 657744 491208 657756
rect 490524 657716 491208 657744
rect 490524 657704 490530 657716
rect 491202 657704 491208 657716
rect 491260 657704 491266 657756
rect 494698 657704 494704 657756
rect 494756 657744 494762 657756
rect 510062 657744 510068 657756
rect 494756 657716 510068 657744
rect 494756 657704 494762 657716
rect 510062 657704 510068 657716
rect 510120 657704 510126 657756
rect 286318 657636 286324 657688
rect 286376 657676 286382 657688
rect 294598 657676 294604 657688
rect 286376 657648 294604 657676
rect 286376 657636 286382 657648
rect 294598 657636 294604 657648
rect 294656 657636 294662 657688
rect 324958 657636 324964 657688
rect 325016 657676 325022 657688
rect 516134 657676 516140 657688
rect 325016 657648 516140 657676
rect 325016 657636 325022 657648
rect 516134 657636 516140 657648
rect 516192 657636 516198 657688
rect 106182 657568 106188 657620
rect 106240 657608 106246 657620
rect 518342 657608 518348 657620
rect 106240 657580 518348 657608
rect 106240 657568 106246 657580
rect 518342 657568 518348 657580
rect 518400 657568 518406 657620
rect 86218 657500 86224 657552
rect 86276 657540 86282 657552
rect 519722 657540 519728 657552
rect 86276 657512 519728 657540
rect 86276 657500 86282 657512
rect 519722 657500 519728 657512
rect 519780 657500 519786 657552
rect 144178 657432 144184 657484
rect 144236 657472 144242 657484
rect 525242 657472 525248 657484
rect 144236 657444 525248 657472
rect 144236 657432 144242 657444
rect 525242 657432 525248 657444
rect 525300 657432 525306 657484
rect 532142 657432 532148 657484
rect 532200 657472 532206 657484
rect 546586 657472 546592 657484
rect 532200 657444 546592 657472
rect 532200 657432 532206 657444
rect 546586 657432 546592 657444
rect 546644 657432 546650 657484
rect 488442 657364 488448 657416
rect 488500 657404 488506 657416
rect 493502 657404 493508 657416
rect 488500 657376 493508 657404
rect 488500 657364 488506 657376
rect 493502 657364 493508 657376
rect 493560 657364 493566 657416
rect 509142 657364 509148 657416
rect 509200 657404 509206 657416
rect 540974 657404 540980 657416
rect 509200 657376 540980 657404
rect 509200 657364 509206 657376
rect 540974 657364 540980 657376
rect 541032 657364 541038 657416
rect 58618 657296 58624 657348
rect 58676 657336 58682 657348
rect 522482 657336 522488 657348
rect 58676 657308 522488 657336
rect 58676 657296 58682 657308
rect 522482 657296 522488 657308
rect 522540 657296 522546 657348
rect 526622 657296 526628 657348
rect 526680 657336 526686 657348
rect 544102 657336 544108 657348
rect 526680 657308 544108 657336
rect 526680 657296 526686 657308
rect 544102 657296 544108 657308
rect 544160 657296 544166 657348
rect 488258 657228 488264 657280
rect 488316 657268 488322 657280
rect 503162 657268 503168 657280
rect 488316 657240 503168 657268
rect 488316 657228 488322 657240
rect 503162 657228 503168 657240
rect 503220 657228 503226 657280
rect 530762 657228 530768 657280
rect 530820 657268 530826 657280
rect 544194 657268 544200 657280
rect 530820 657240 544200 657268
rect 530820 657228 530826 657240
rect 544194 657228 544200 657240
rect 544252 657228 544258 657280
rect 490558 657160 490564 657212
rect 490616 657200 490622 657212
rect 491110 657200 491116 657212
rect 490616 657172 491116 657200
rect 490616 657160 490622 657172
rect 491110 657160 491116 657172
rect 491168 657200 491174 657212
rect 511442 657200 511448 657212
rect 491168 657172 511448 657200
rect 491168 657160 491174 657172
rect 511442 657160 511448 657172
rect 511500 657160 511506 657212
rect 528002 657160 528008 657212
rect 528060 657200 528066 657212
rect 544010 657200 544016 657212
rect 528060 657172 544016 657200
rect 528060 657160 528066 657172
rect 544010 657160 544016 657172
rect 544068 657160 544074 657212
rect 491202 657092 491208 657144
rect 491260 657132 491266 657144
rect 514202 657132 514208 657144
rect 491260 657104 514208 657132
rect 491260 657092 491266 657104
rect 514202 657092 514208 657104
rect 514260 657092 514266 657144
rect 529382 657092 529388 657144
rect 529440 657132 529446 657144
rect 545390 657132 545396 657144
rect 529440 657104 545396 657132
rect 529440 657092 529446 657104
rect 545390 657092 545396 657104
rect 545448 657092 545454 657144
rect 485682 657024 485688 657076
rect 485740 657064 485746 657076
rect 494882 657064 494888 657076
rect 485740 657036 494888 657064
rect 485740 657024 485746 657036
rect 494882 657024 494888 657036
rect 494940 657024 494946 657076
rect 512822 657064 512828 657076
rect 499546 657036 512828 657064
rect 490374 656956 490380 657008
rect 490432 656996 490438 657008
rect 491018 656996 491024 657008
rect 490432 656968 491024 656996
rect 490432 656956 490438 656968
rect 491018 656956 491024 656968
rect 491076 656996 491082 657008
rect 499546 656996 499574 657036
rect 512822 657024 512828 657036
rect 512880 657024 512886 657076
rect 534902 657024 534908 657076
rect 534960 657064 534966 657076
rect 547966 657064 547972 657076
rect 534960 657036 547972 657064
rect 534960 657024 534966 657036
rect 547966 657024 547972 657036
rect 548024 657024 548030 657076
rect 491076 656968 499574 656996
rect 491076 656956 491082 656968
rect 533522 656956 533528 657008
rect 533580 656996 533586 657008
rect 545482 656996 545488 657008
rect 533580 656968 545488 656996
rect 533580 656956 533586 656968
rect 545482 656956 545488 656968
rect 545540 656956 545546 657008
rect 516134 656888 516140 656940
rect 516192 656928 516198 656940
rect 516962 656928 516968 656940
rect 516192 656900 516968 656928
rect 516192 656888 516198 656900
rect 516962 656888 516968 656900
rect 517020 656928 517026 656940
rect 540330 656928 540336 656940
rect 517020 656900 540336 656928
rect 517020 656888 517026 656900
rect 540330 656888 540336 656900
rect 540388 656888 540394 656940
rect 366358 656820 366364 656872
rect 366416 656860 366422 656872
rect 371878 656860 371884 656872
rect 366416 656832 371884 656860
rect 366416 656820 366422 656832
rect 371878 656820 371884 656832
rect 371936 656820 371942 656872
rect 505922 655596 505928 655648
rect 505980 655636 505986 655648
rect 540422 655636 540428 655648
rect 505980 655608 540428 655636
rect 505980 655596 505986 655608
rect 540422 655596 540428 655608
rect 540480 655596 540486 655648
rect 504542 655528 504548 655580
rect 504600 655568 504606 655580
rect 543734 655568 543740 655580
rect 504600 655540 543740 655568
rect 504600 655528 504606 655540
rect 543734 655528 543740 655540
rect 543792 655528 543798 655580
rect 239398 655460 239404 655512
rect 239456 655500 239462 655512
rect 242434 655500 242440 655512
rect 239456 655472 242440 655500
rect 239456 655460 239462 655472
rect 242434 655460 242440 655472
rect 242492 655460 242498 655512
rect 355962 654780 355968 654832
rect 356020 654820 356026 654832
rect 366358 654820 366364 654832
rect 356020 654792 366364 654820
rect 356020 654780 356026 654792
rect 366358 654780 366364 654792
rect 366416 654780 366422 654832
rect 486878 654576 486884 654628
rect 486936 654616 486942 654628
rect 498654 654616 498660 654628
rect 486936 654588 498660 654616
rect 486936 654576 486942 654588
rect 498654 654576 498660 654588
rect 498712 654576 498718 654628
rect 156598 654508 156604 654560
rect 156656 654548 156662 654560
rect 523494 654548 523500 654560
rect 156656 654520 523500 654548
rect 156656 654508 156662 654520
rect 523494 654508 523500 654520
rect 523552 654508 523558 654560
rect 489638 654440 489644 654492
rect 489696 654480 489702 654492
rect 491846 654480 491852 654492
rect 489696 654452 491852 654480
rect 489696 654440 489702 654452
rect 491846 654440 491852 654452
rect 491904 654440 491910 654492
rect 497366 654440 497372 654492
rect 497424 654440 497430 654492
rect 485590 654372 485596 654424
rect 485648 654412 485654 654424
rect 497384 654412 497412 654440
rect 485648 654384 497412 654412
rect 485648 654372 485654 654384
rect 488442 654236 488448 654288
rect 488500 654276 488506 654288
rect 490650 654276 490656 654288
rect 488500 654248 490656 654276
rect 488500 654236 488506 654248
rect 490650 654236 490656 654248
rect 490708 654236 490714 654288
rect 178034 654100 178040 654152
rect 178092 654140 178098 654152
rect 368382 654140 368388 654152
rect 178092 654112 368388 654140
rect 178092 654100 178098 654112
rect 368382 654100 368388 654112
rect 368440 654100 368446 654152
rect 371878 651992 371884 652044
rect 371936 652032 371942 652044
rect 377398 652032 377404 652044
rect 371936 652004 377404 652032
rect 371936 651992 371942 652004
rect 377398 651992 377404 652004
rect 377456 651992 377462 652044
rect 213822 651516 213828 651568
rect 213880 651556 213886 651568
rect 361942 651556 361948 651568
rect 213880 651528 361948 651556
rect 213880 651516 213886 651528
rect 361942 651516 361948 651528
rect 362000 651516 362006 651568
rect 233142 651448 233148 651500
rect 233200 651488 233206 651500
rect 464338 651488 464344 651500
rect 233200 651460 464344 651488
rect 233200 651448 233206 651460
rect 464338 651448 464344 651460
rect 464396 651448 464402 651500
rect 227714 651380 227720 651432
rect 227772 651420 227778 651432
rect 483658 651420 483664 651432
rect 227772 651392 483664 651420
rect 227772 651380 227778 651392
rect 483658 651380 483664 651392
rect 483716 651380 483722 651432
rect 231762 650292 231768 650344
rect 231820 650332 231826 650344
rect 374362 650332 374368 650344
rect 231820 650304 374368 650332
rect 231820 650292 231826 650304
rect 374362 650292 374368 650304
rect 374420 650292 374426 650344
rect 226334 650224 226340 650276
rect 226392 650264 226398 650276
rect 375650 650264 375656 650276
rect 226392 650236 375656 650264
rect 226392 650224 226398 650236
rect 375650 650224 375656 650236
rect 375708 650224 375714 650276
rect 214558 650156 214564 650208
rect 214616 650196 214622 650208
rect 374822 650196 374828 650208
rect 214616 650168 374828 650196
rect 214616 650156 214622 650168
rect 374822 650156 374828 650168
rect 374880 650156 374886 650208
rect 212442 650088 212448 650140
rect 212500 650128 212506 650140
rect 374546 650128 374552 650140
rect 212500 650100 374552 650128
rect 212500 650088 212506 650100
rect 374546 650088 374552 650100
rect 374604 650088 374610 650140
rect 186314 650020 186320 650072
rect 186372 650060 186378 650072
rect 374730 650060 374736 650072
rect 186372 650032 374736 650060
rect 186372 650020 186378 650032
rect 374730 650020 374736 650032
rect 374788 650020 374794 650072
rect 543550 650020 543556 650072
rect 543608 650060 543614 650072
rect 549254 650060 549260 650072
rect 543608 650032 549260 650060
rect 543608 650020 543614 650032
rect 549254 650020 549260 650032
rect 549312 650020 549318 650072
rect 205634 648796 205640 648848
rect 205692 648836 205698 648848
rect 467098 648836 467104 648848
rect 205692 648808 467104 648836
rect 205692 648796 205698 648808
rect 467098 648796 467104 648808
rect 467156 648796 467162 648848
rect 224218 648728 224224 648780
rect 224276 648768 224282 648780
rect 486418 648768 486424 648780
rect 224276 648740 486424 648768
rect 224276 648728 224282 648740
rect 486418 648728 486424 648740
rect 486476 648728 486482 648780
rect 199654 648660 199660 648712
rect 199712 648700 199718 648712
rect 469950 648700 469956 648712
rect 199712 648672 469956 648700
rect 199712 648660 199718 648672
rect 469950 648660 469956 648672
rect 470008 648660 470014 648712
rect 198734 648592 198740 648644
rect 198792 648632 198798 648644
rect 472618 648632 472624 648644
rect 198792 648604 472624 648632
rect 198792 648592 198798 648604
rect 472618 648592 472624 648604
rect 472676 648592 472682 648644
rect 234614 647504 234620 647556
rect 234672 647544 234678 647556
rect 354214 647544 354220 647556
rect 234672 647516 354220 647544
rect 234672 647504 234678 647516
rect 354214 647504 354220 647516
rect 354272 647504 354278 647556
rect 217502 647436 217508 647488
rect 217560 647476 217566 647488
rect 472894 647476 472900 647488
rect 217560 647448 472900 647476
rect 217560 647436 217566 647448
rect 472894 647436 472900 647448
rect 472952 647436 472958 647488
rect 203334 647368 203340 647420
rect 203392 647408 203398 647420
rect 471238 647408 471244 647420
rect 203392 647380 471244 647408
rect 203392 647368 203398 647380
rect 471238 647368 471244 647380
rect 471296 647368 471302 647420
rect 176562 647300 176568 647352
rect 176620 647340 176626 647352
rect 478138 647340 478144 647352
rect 176620 647312 478144 647340
rect 176620 647300 176626 647312
rect 478138 647300 478144 647312
rect 478196 647300 478202 647352
rect 54386 647232 54392 647284
rect 54444 647272 54450 647284
rect 372246 647272 372252 647284
rect 54444 647244 372252 647272
rect 54444 647232 54450 647244
rect 372246 647232 372252 647244
rect 372304 647232 372310 647284
rect 366358 647164 366364 647216
rect 366416 647204 366422 647216
rect 371878 647204 371884 647216
rect 366416 647176 371884 647204
rect 366416 647164 366422 647176
rect 371878 647164 371884 647176
rect 371936 647164 371942 647216
rect 294598 646484 294604 646536
rect 294656 646524 294662 646536
rect 304258 646524 304264 646536
rect 294656 646496 304264 646524
rect 294656 646484 294662 646496
rect 304258 646484 304264 646496
rect 304316 646484 304322 646536
rect 115842 646144 115848 646196
rect 115900 646184 115906 646196
rect 325878 646184 325884 646196
rect 115900 646156 325884 646184
rect 115900 646144 115906 646156
rect 325878 646144 325884 646156
rect 325936 646144 325942 646196
rect 240686 646076 240692 646128
rect 240744 646116 240750 646128
rect 462958 646116 462964 646128
rect 240744 646088 462964 646116
rect 240744 646076 240750 646088
rect 462958 646076 462964 646088
rect 463016 646076 463022 646128
rect 209774 646008 209780 646060
rect 209832 646048 209838 646060
rect 483750 646048 483756 646060
rect 209832 646020 483756 646048
rect 209832 646008 209838 646020
rect 483750 646008 483756 646020
rect 483808 646008 483814 646060
rect 204622 645940 204628 645992
rect 204680 645980 204686 645992
rect 482370 645980 482376 645992
rect 204680 645952 482376 645980
rect 204680 645940 204686 645952
rect 482370 645940 482376 645952
rect 482428 645940 482434 645992
rect 151078 645912 151084 645924
rect 149072 645884 151084 645912
rect 146202 645804 146208 645856
rect 146260 645844 146266 645856
rect 149072 645844 149100 645884
rect 151078 645872 151084 645884
rect 151136 645872 151142 645924
rect 176562 645872 176568 645924
rect 176620 645912 176626 645924
rect 479702 645912 479708 645924
rect 176620 645884 479708 645912
rect 176620 645872 176626 645884
rect 479702 645872 479708 645884
rect 479760 645872 479766 645924
rect 146260 645816 149100 645844
rect 146260 645804 146266 645816
rect 177298 644784 177304 644836
rect 177356 644824 177362 644836
rect 393222 644824 393228 644836
rect 177356 644796 393228 644824
rect 177356 644784 177362 644796
rect 393222 644784 393228 644796
rect 393280 644784 393286 644836
rect 218790 644716 218796 644768
rect 218848 644756 218854 644768
rect 464430 644756 464436 644768
rect 218848 644728 464436 644756
rect 218848 644716 218854 644728
rect 464430 644716 464436 644728
rect 464488 644716 464494 644768
rect 230382 644648 230388 644700
rect 230440 644688 230446 644700
rect 476758 644688 476764 644700
rect 230440 644660 476764 644688
rect 230440 644648 230446 644660
rect 476758 644648 476764 644660
rect 476816 644648 476822 644700
rect 138658 644580 138664 644632
rect 138716 644620 138722 644632
rect 390186 644620 390192 644632
rect 138716 644592 390192 644620
rect 138716 644580 138722 644592
rect 390186 644580 390192 644592
rect 390244 644580 390250 644632
rect 131114 644512 131120 644564
rect 131172 644552 131178 644564
rect 384114 644552 384120 644564
rect 131172 644524 384120 644552
rect 131172 644512 131178 644524
rect 384114 644512 384120 644524
rect 384172 644512 384178 644564
rect 91094 644444 91100 644496
rect 91152 644484 91158 644496
rect 351638 644484 351644 644496
rect 91152 644456 351644 644484
rect 91152 644444 91158 644456
rect 351638 644444 351644 644456
rect 351696 644444 351702 644496
rect 186958 643696 186964 643748
rect 187016 643736 187022 643748
rect 239398 643736 239404 643748
rect 187016 643708 239404 643736
rect 187016 643696 187022 643708
rect 239398 643696 239404 643708
rect 239456 643696 239462 643748
rect 176746 643492 176752 643544
rect 176804 643532 176810 643544
rect 389174 643532 389180 643544
rect 176804 643504 389180 643532
rect 176804 643492 176810 643504
rect 389174 643492 389180 643504
rect 389232 643492 389238 643544
rect 126882 643424 126888 643476
rect 126940 643464 126946 643476
rect 338758 643464 338764 643476
rect 126940 643436 338764 643464
rect 126940 643424 126946 643436
rect 338758 643424 338764 643436
rect 338816 643424 338822 643476
rect 176654 643356 176660 643408
rect 176712 643396 176718 643408
rect 419534 643396 419540 643408
rect 176712 643368 419540 643396
rect 176712 643356 176718 643368
rect 419534 643356 419540 643368
rect 419592 643356 419598 643408
rect 124122 643288 124128 643340
rect 124180 643328 124186 643340
rect 365806 643328 365812 643340
rect 124180 643300 365812 643328
rect 124180 643288 124186 643300
rect 365806 643288 365812 643300
rect 365864 643288 365870 643340
rect 377398 643288 377404 643340
rect 377456 643328 377462 643340
rect 380526 643328 380532 643340
rect 377456 643300 380532 643328
rect 377456 643288 377462 643300
rect 380526 643288 380532 643300
rect 380584 643288 380590 643340
rect 221734 643220 221740 643272
rect 221792 643260 221798 643272
rect 464522 643260 464528 643272
rect 221792 643232 464528 643260
rect 221792 643220 221798 643232
rect 464522 643220 464528 643232
rect 464580 643220 464586 643272
rect 225506 643152 225512 643204
rect 225564 643192 225570 643204
rect 483842 643192 483848 643204
rect 225564 643164 483848 643192
rect 225564 643152 225570 643164
rect 483842 643152 483848 643164
rect 483900 643152 483906 643204
rect 198458 643084 198464 643136
rect 198516 643124 198522 643136
rect 472710 643124 472716 643136
rect 198516 643096 472716 643124
rect 198516 643084 198522 643096
rect 472710 643084 472716 643096
rect 472768 643084 472774 643136
rect 294046 642404 294052 642456
rect 294104 642444 294110 642456
rect 340046 642444 340052 642456
rect 294104 642416 340052 642444
rect 294104 642404 294110 642416
rect 340046 642404 340052 642416
rect 340104 642404 340110 642456
rect 293954 642336 293960 642388
rect 294012 642376 294018 642388
rect 382090 642376 382096 642388
rect 294012 642348 382096 642376
rect 294012 642336 294018 642348
rect 382090 642336 382096 642348
rect 382148 642336 382154 642388
rect 178034 642268 178040 642320
rect 178092 642308 178098 642320
rect 346486 642308 346492 642320
rect 178092 642280 346492 642308
rect 178092 642268 178098 642280
rect 346486 642268 346492 642280
rect 346544 642268 346550 642320
rect 153930 642200 153936 642252
rect 153988 642240 153994 642252
rect 375558 642240 375564 642252
rect 153988 642212 375564 642240
rect 153988 642200 153994 642212
rect 375558 642200 375564 642212
rect 375616 642200 375622 642252
rect 216582 642132 216588 642184
rect 216640 642172 216646 642184
rect 464614 642172 464620 642184
rect 216640 642144 464620 642172
rect 216640 642132 216646 642144
rect 464614 642132 464620 642144
rect 464672 642132 464678 642184
rect 202414 642064 202420 642116
rect 202472 642104 202478 642116
rect 482554 642104 482560 642116
rect 202472 642076 482560 642104
rect 202472 642064 202478 642076
rect 482554 642064 482560 642076
rect 482612 642064 482618 642116
rect 177942 641996 177948 642048
rect 178000 642036 178006 642048
rect 458818 642036 458824 642048
rect 178000 642008 458824 642036
rect 178000 641996 178006 642008
rect 458818 641996 458824 642008
rect 458876 641996 458882 642048
rect 59262 641928 59268 641980
rect 59320 641968 59326 641980
rect 350350 641968 350356 641980
rect 59320 641940 350356 641968
rect 59320 641928 59326 641940
rect 350350 641928 350356 641940
rect 350408 641928 350414 641980
rect 144270 641860 144276 641912
rect 144328 641900 144334 641912
rect 146202 641900 146208 641912
rect 144328 641872 146208 641900
rect 144328 641860 144334 641872
rect 146202 641860 146208 641872
rect 146260 641860 146266 641912
rect 183094 641860 183100 641912
rect 183152 641900 183158 641912
rect 475470 641900 475476 641912
rect 183152 641872 475476 641900
rect 183152 641860 183158 641872
rect 475470 641860 475476 641872
rect 475528 641860 475534 641912
rect 59262 641792 59268 641844
rect 59320 641832 59326 641844
rect 352926 641832 352932 641844
rect 59320 641804 352932 641832
rect 59320 641792 59326 641804
rect 352926 641792 352932 641804
rect 352984 641792 352990 641844
rect 57882 641724 57888 641776
rect 57940 641764 57946 641776
rect 355502 641764 355508 641776
rect 57940 641736 355508 641764
rect 57940 641724 57946 641736
rect 355502 641724 355508 641736
rect 355560 641724 355566 641776
rect 380526 640976 380532 641028
rect 380584 641016 380590 641028
rect 387794 641016 387800 641028
rect 380584 640988 387800 641016
rect 380584 640976 380590 640988
rect 387794 640976 387800 640988
rect 387852 640976 387858 641028
rect 251082 640908 251088 640960
rect 251140 640948 251146 640960
rect 320726 640948 320732 640960
rect 251140 640920 320732 640948
rect 251140 640908 251146 640920
rect 320726 640908 320732 640920
rect 320784 640908 320790 640960
rect 249702 640840 249708 640892
rect 249760 640880 249766 640892
rect 322014 640880 322020 640892
rect 249760 640852 322020 640880
rect 249760 640840 249766 640852
rect 322014 640840 322020 640852
rect 322072 640840 322078 640892
rect 127618 640772 127624 640824
rect 127676 640812 127682 640824
rect 331030 640812 331036 640824
rect 127676 640784 331036 640812
rect 127676 640772 127682 640784
rect 331030 640772 331036 640784
rect 331088 640772 331094 640824
rect 222930 640704 222936 640756
rect 222988 640744 222994 640756
rect 465810 640744 465816 640756
rect 222988 640716 465816 640744
rect 222988 640704 222994 640716
rect 465810 640704 465816 640716
rect 465868 640704 465874 640756
rect 195882 640636 195888 640688
rect 195940 640676 195946 640688
rect 472802 640676 472808 640688
rect 195940 640648 472808 640676
rect 195940 640636 195946 640648
rect 472802 640636 472808 640648
rect 472860 640636 472866 640688
rect 59262 640568 59268 640620
rect 59320 640608 59326 640620
rect 337470 640608 337476 640620
rect 59320 640580 337476 640608
rect 59320 640568 59326 640580
rect 337470 640568 337476 640580
rect 337528 640568 337534 640620
rect 177574 640500 177580 640552
rect 177632 640540 177638 640552
rect 458910 640540 458916 640552
rect 177632 640512 458916 640540
rect 177632 640500 177638 640512
rect 458910 640500 458916 640512
rect 458968 640500 458974 640552
rect 56502 640432 56508 640484
rect 56560 640472 56566 640484
rect 349062 640472 349068 640484
rect 56560 640444 349068 640472
rect 56560 640432 56566 640444
rect 349062 640432 349068 640444
rect 349120 640432 349126 640484
rect 193122 640364 193128 640416
rect 193180 640404 193186 640416
rect 489362 640404 489368 640416
rect 193180 640376 489368 640404
rect 193180 640364 193186 640376
rect 489362 640364 489368 640376
rect 489420 640364 489426 640416
rect 148318 640296 148324 640348
rect 148376 640336 148382 640348
rect 149698 640336 149704 640348
rect 148376 640308 149704 640336
rect 148376 640296 148382 640308
rect 149698 640296 149704 640308
rect 149756 640296 149762 640348
rect 177942 640296 177948 640348
rect 178000 640336 178006 640348
rect 489178 640336 489184 640348
rect 178000 640308 489184 640336
rect 178000 640296 178006 640308
rect 489178 640296 489184 640308
rect 489236 640296 489242 640348
rect 109034 639548 109040 639600
rect 109092 639588 109098 639600
rect 309134 639588 309140 639600
rect 109092 639560 309140 639588
rect 109092 639548 109098 639560
rect 309134 639548 309140 639560
rect 309192 639548 309198 639600
rect 88978 639480 88984 639532
rect 89036 639520 89042 639532
rect 318150 639520 318156 639532
rect 89036 639492 318156 639520
rect 89036 639480 89042 639492
rect 318150 639480 318156 639492
rect 318208 639480 318214 639532
rect 220354 639412 220360 639464
rect 220412 639452 220418 639464
rect 471514 639452 471520 639464
rect 220412 639424 471520 639452
rect 220412 639412 220418 639424
rect 471514 639412 471520 639424
rect 471572 639412 471578 639464
rect 154482 639344 154488 639396
rect 154540 639384 154546 639396
rect 421558 639384 421564 639396
rect 154540 639356 421564 639384
rect 154540 639344 154546 639356
rect 421558 639344 421564 639356
rect 421616 639344 421622 639396
rect 88242 639276 88248 639328
rect 88300 639316 88306 639328
rect 385126 639316 385132 639328
rect 88300 639288 385132 639316
rect 88300 639276 88306 639288
rect 385126 639276 385132 639288
rect 385184 639276 385190 639328
rect 106182 639208 106188 639260
rect 106240 639248 106246 639260
rect 403342 639248 403348 639260
rect 106240 639220 403348 639248
rect 106240 639208 106246 639220
rect 403342 639208 403348 639220
rect 403400 639208 403406 639260
rect 107562 639140 107568 639192
rect 107620 639180 107626 639192
rect 405366 639180 405372 639192
rect 107620 639152 405372 639180
rect 107620 639140 107626 639152
rect 405366 639140 405372 639152
rect 405424 639140 405430 639192
rect 66162 639072 66168 639124
rect 66220 639112 66226 639124
rect 376846 639112 376852 639124
rect 66220 639084 376852 639112
rect 66220 639072 66226 639084
rect 376846 639072 376852 639084
rect 376904 639072 376910 639124
rect 88794 639004 88800 639056
rect 88852 639044 88858 639056
rect 403618 639044 403624 639056
rect 88852 639016 403624 639044
rect 88852 639004 88858 639016
rect 403618 639004 403624 639016
rect 403676 639004 403682 639056
rect 91002 638936 91008 638988
rect 91060 638976 91066 638988
rect 406378 638976 406384 638988
rect 91060 638948 406384 638976
rect 91060 638936 91066 638948
rect 406378 638936 406384 638948
rect 406436 638936 406442 638988
rect 234522 638324 234528 638376
rect 234580 638364 234586 638376
rect 291838 638364 291844 638376
rect 234580 638336 291844 638364
rect 234580 638324 234586 638336
rect 291838 638324 291844 638336
rect 291896 638324 291902 638376
rect 137278 638256 137284 638308
rect 137336 638296 137342 638308
rect 312998 638296 313004 638308
rect 137336 638268 313004 638296
rect 137336 638256 137342 638268
rect 312998 638256 313004 638268
rect 313056 638256 313062 638308
rect 227714 638188 227720 638240
rect 227772 638228 227778 638240
rect 414658 638228 414664 638240
rect 227772 638200 414664 638228
rect 227772 638188 227778 638200
rect 414658 638188 414664 638200
rect 414716 638188 414722 638240
rect 252462 638120 252468 638172
rect 252520 638160 252526 638172
rect 475654 638160 475660 638172
rect 252520 638132 475660 638160
rect 252520 638120 252526 638132
rect 475654 638120 475660 638132
rect 475712 638120 475718 638172
rect 86862 638052 86868 638104
rect 86920 638092 86926 638104
rect 319438 638092 319444 638104
rect 86920 638064 319444 638092
rect 86920 638052 86926 638064
rect 319438 638052 319444 638064
rect 319496 638052 319502 638104
rect 129734 637984 129740 638036
rect 129792 638024 129798 638036
rect 400858 638024 400864 638036
rect 129792 637996 400864 638024
rect 129792 637984 129798 637996
rect 400858 637984 400864 637996
rect 400916 637984 400922 638036
rect 118694 637916 118700 637968
rect 118752 637956 118758 637968
rect 397270 637956 397276 637968
rect 118752 637928 397276 637956
rect 118752 637916 118758 637928
rect 397270 637916 397276 637928
rect 397328 637916 397334 637968
rect 179046 637848 179052 637900
rect 179104 637888 179110 637900
rect 463234 637888 463240 637900
rect 179104 637860 463240 637888
rect 179104 637848 179110 637860
rect 463234 637848 463240 637860
rect 463292 637848 463298 637900
rect 81434 637780 81440 637832
rect 81492 637820 81498 637832
rect 367094 637820 367100 637832
rect 81492 637792 367100 637820
rect 81492 637780 81498 637792
rect 367094 637780 367100 637792
rect 367152 637780 367158 637832
rect 110414 637712 110420 637764
rect 110472 637752 110478 637764
rect 399294 637752 399300 637764
rect 110472 637724 399300 637752
rect 110472 637712 110478 637724
rect 399294 637712 399300 637724
rect 399352 637712 399358 637764
rect 102134 637644 102140 637696
rect 102192 637684 102198 637696
rect 400306 637684 400312 637696
rect 102192 637656 400312 637684
rect 102192 637644 102198 637656
rect 400306 637644 400312 637656
rect 400364 637644 400370 637696
rect 82814 637576 82820 637628
rect 82872 637616 82878 637628
rect 395338 637616 395344 637628
rect 82872 637588 395344 637616
rect 82872 637576 82878 637588
rect 395338 637576 395344 637588
rect 395396 637576 395402 637628
rect 73154 637508 73160 637560
rect 73212 637548 73218 637560
rect 176746 637548 176752 637560
rect 73212 637520 176752 637548
rect 73212 637508 73218 637520
rect 176746 637508 176752 637520
rect 176804 637508 176810 637560
rect 108298 637440 108304 637492
rect 108356 637480 108362 637492
rect 177298 637480 177304 637492
rect 108356 637452 177304 637480
rect 108356 637440 108362 637452
rect 177298 637440 177304 637452
rect 177356 637440 177362 637492
rect 117958 637372 117964 637424
rect 118016 637412 118022 637424
rect 176654 637412 176660 637424
rect 118016 637384 176660 637412
rect 118016 637372 118022 637384
rect 176654 637372 176660 637384
rect 176712 637372 176718 637424
rect 117222 637304 117228 637356
rect 117280 637344 117286 637356
rect 138658 637344 138664 637356
rect 117280 637316 138664 637344
rect 117280 637304 117286 637316
rect 138658 637304 138664 637316
rect 138716 637304 138722 637356
rect 128354 636964 128360 637016
rect 128412 637004 128418 637016
rect 292022 637004 292028 637016
rect 128412 636976 292028 637004
rect 128412 636964 128418 636976
rect 292022 636964 292028 636976
rect 292080 636964 292086 637016
rect 128446 636896 128452 636948
rect 128504 636936 128510 636948
rect 297450 636936 297456 636948
rect 128504 636908 297456 636936
rect 128504 636896 128510 636908
rect 297450 636896 297456 636908
rect 297508 636896 297514 636948
rect 125502 636828 125508 636880
rect 125560 636868 125566 636880
rect 297358 636868 297364 636880
rect 125560 636840 297364 636868
rect 125560 636828 125566 636840
rect 297358 636828 297364 636840
rect 297416 636828 297422 636880
rect 121454 636760 121460 636812
rect 121512 636800 121518 636812
rect 306558 636800 306564 636812
rect 121512 636772 306564 636800
rect 121512 636760 121518 636772
rect 306558 636760 306564 636772
rect 306616 636760 306622 636812
rect 245562 636692 245568 636744
rect 245620 636732 245626 636744
rect 456150 636732 456156 636744
rect 245620 636704 456156 636732
rect 245620 636692 245626 636704
rect 456150 636692 456156 636704
rect 456208 636692 456214 636744
rect 242802 636624 242808 636676
rect 242860 636664 242866 636676
rect 459002 636664 459008 636676
rect 242860 636636 459008 636664
rect 242860 636624 242866 636636
rect 459002 636624 459008 636636
rect 459060 636624 459066 636676
rect 235994 636556 236000 636608
rect 236052 636596 236058 636608
rect 456058 636596 456064 636608
rect 236052 636568 456064 636596
rect 236052 636556 236058 636568
rect 456058 636556 456064 636568
rect 456116 636556 456122 636608
rect 246942 636488 246948 636540
rect 247000 636528 247006 636540
rect 486510 636528 486516 636540
rect 247000 636500 486516 636528
rect 247000 636488 247006 636500
rect 486510 636488 486516 636500
rect 486568 636488 486574 636540
rect 240042 636420 240048 636472
rect 240100 636460 240106 636472
rect 489454 636460 489460 636472
rect 240100 636432 489460 636460
rect 240100 636420 240106 636432
rect 489454 636420 489460 636432
rect 489512 636420 489518 636472
rect 179322 636352 179328 636404
rect 179380 636392 179386 636404
rect 453298 636392 453304 636404
rect 179380 636364 453304 636392
rect 179380 636352 179386 636364
rect 453298 636352 453304 636364
rect 453356 636352 453362 636404
rect 191742 636284 191748 636336
rect 191800 636324 191806 636336
rect 472986 636324 472992 636336
rect 191800 636296 472992 636324
rect 191800 636284 191806 636296
rect 472986 636284 472992 636296
rect 473044 636284 473050 636336
rect 179966 636216 179972 636268
rect 180024 636256 180030 636268
rect 485130 636256 485136 636268
rect 180024 636228 485136 636256
rect 180024 636216 180030 636228
rect 485130 636216 485136 636228
rect 485188 636216 485194 636268
rect 387794 636148 387800 636200
rect 387852 636188 387858 636200
rect 391382 636188 391388 636200
rect 387852 636160 391388 636188
rect 387852 636148 387858 636160
rect 391382 636148 391388 636160
rect 391440 636148 391446 636200
rect 38562 635468 38568 635520
rect 38620 635508 38626 635520
rect 72970 635508 72976 635520
rect 38620 635480 72976 635508
rect 38620 635468 38626 635480
rect 72970 635468 72976 635480
rect 73028 635468 73034 635520
rect 156690 635468 156696 635520
rect 156748 635508 156754 635520
rect 375374 635508 375380 635520
rect 156748 635480 375380 635508
rect 156748 635468 156754 635480
rect 375374 635468 375380 635480
rect 375432 635468 375438 635520
rect 247586 635400 247592 635452
rect 247644 635440 247650 635452
rect 471422 635440 471428 635452
rect 247644 635412 471428 635440
rect 247644 635400 247650 635412
rect 471422 635400 471428 635412
rect 471480 635400 471486 635452
rect 92474 635332 92480 635384
rect 92532 635372 92538 635384
rect 342622 635372 342628 635384
rect 92532 635344 342628 635372
rect 92532 635332 92538 635344
rect 342622 635332 342628 635344
rect 342680 635332 342686 635384
rect 99374 635264 99380 635316
rect 99432 635304 99438 635316
rect 391290 635304 391296 635316
rect 99432 635276 391296 635304
rect 99432 635264 99438 635276
rect 391290 635264 391296 635276
rect 391348 635264 391354 635316
rect 95142 635196 95148 635248
rect 95200 635236 95206 635248
rect 386138 635236 386144 635248
rect 95200 635208 386144 635236
rect 95200 635196 95206 635208
rect 386138 635196 386144 635208
rect 386196 635196 386202 635248
rect 109126 635128 109132 635180
rect 109184 635168 109190 635180
rect 412450 635168 412456 635180
rect 109184 635140 412456 635168
rect 109184 635128 109190 635140
rect 412450 635128 412456 635140
rect 412508 635128 412514 635180
rect 104802 635060 104808 635112
rect 104860 635100 104866 635112
rect 410518 635100 410524 635112
rect 104860 635072 410524 635100
rect 104860 635060 104866 635072
rect 410518 635060 410524 635072
rect 410576 635060 410582 635112
rect 98086 634992 98092 635044
rect 98144 635032 98150 635044
rect 409414 635032 409420 635044
rect 98144 635004 409420 635032
rect 98144 634992 98150 635004
rect 409414 634992 409420 635004
rect 409472 634992 409478 635044
rect 96522 634924 96528 634976
rect 96580 634964 96586 634976
rect 407758 634964 407764 634976
rect 96580 634936 407764 634964
rect 96580 634924 96586 634936
rect 407758 634924 407764 634936
rect 407816 634924 407822 634976
rect 101674 634856 101680 634908
rect 101732 634896 101738 634908
rect 414474 634896 414480 634908
rect 101732 634868 414480 634896
rect 101732 634856 101738 634868
rect 414474 634856 414480 634868
rect 414532 634856 414538 634908
rect 97810 634788 97816 634840
rect 97868 634828 97874 634840
rect 411438 634828 411444 634840
rect 97868 634800 411444 634828
rect 97868 634788 97874 634800
rect 411438 634788 411444 634800
rect 411496 634788 411502 634840
rect 151078 634448 151084 634500
rect 151136 634488 151142 634500
rect 376754 634488 376760 634500
rect 151136 634460 376760 634488
rect 151136 634448 151142 634460
rect 376754 634448 376760 634460
rect 376812 634448 376818 634500
rect 171962 634380 171968 634432
rect 172020 634420 172026 634432
rect 186958 634420 186964 634432
rect 172020 634392 186964 634420
rect 172020 634380 172026 634392
rect 186958 634380 186964 634392
rect 187016 634380 187022 634432
rect 371878 634380 371884 634432
rect 371936 634420 371942 634432
rect 387702 634420 387708 634432
rect 371936 634392 387708 634420
rect 371936 634380 371942 634392
rect 387702 634380 387708 634392
rect 387760 634380 387766 634432
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 31570 632108 31576 632120
rect 3476 632080 31576 632108
rect 3476 632068 3482 632080
rect 31570 632068 31576 632080
rect 31628 632108 31634 632120
rect 31628 632080 55214 632108
rect 31628 632068 31634 632080
rect 55186 632040 55214 632080
rect 58618 632040 58624 632052
rect 55186 632012 58624 632040
rect 58618 632000 58624 632012
rect 58676 632000 58682 632052
rect 146938 630640 146944 630692
rect 146996 630680 147002 630692
rect 148318 630680 148324 630692
rect 146996 630652 148324 630680
rect 146996 630640 147002 630652
rect 148318 630640 148324 630652
rect 148376 630640 148382 630692
rect 387702 627172 387708 627224
rect 387760 627212 387766 627224
rect 400766 627212 400772 627224
rect 387760 627184 400772 627212
rect 387760 627172 387766 627184
rect 400766 627172 400772 627184
rect 400824 627172 400830 627224
rect 377214 622412 377220 622464
rect 377272 622452 377278 622464
rect 380158 622452 380164 622464
rect 377272 622424 380164 622452
rect 377272 622412 377278 622424
rect 380158 622412 380164 622424
rect 380216 622412 380222 622464
rect 391382 621664 391388 621716
rect 391440 621704 391446 621716
rect 398098 621704 398104 621716
rect 391440 621676 398104 621704
rect 391440 621664 391446 621676
rect 398098 621664 398104 621676
rect 398156 621664 398162 621716
rect 400766 621664 400772 621716
rect 400824 621704 400830 621716
rect 406470 621704 406476 621716
rect 400824 621676 406476 621704
rect 400824 621664 400830 621676
rect 406470 621664 406476 621676
rect 406528 621664 406534 621716
rect 144914 620984 144920 621036
rect 144972 621024 144978 621036
rect 146938 621024 146944 621036
rect 144972 620996 146944 621024
rect 144972 620984 144978 620996
rect 146938 620984 146944 620996
rect 146996 620984 147002 621036
rect 282178 619624 282184 619676
rect 282236 619664 282242 619676
rect 298002 619664 298008 619676
rect 282236 619636 298008 619664
rect 282236 619624 282242 619636
rect 298002 619624 298008 619636
rect 298060 619624 298066 619676
rect 142798 619556 142804 619608
rect 142856 619596 142862 619608
rect 144914 619596 144920 619608
rect 142856 619568 144920 619596
rect 142856 619556 142862 619568
rect 144914 619556 144920 619568
rect 144972 619556 144978 619608
rect 289078 618264 289084 618316
rect 289136 618304 289142 618316
rect 298002 618304 298008 618316
rect 289136 618276 298008 618304
rect 289136 618264 289142 618276
rect 298002 618264 298008 618276
rect 298060 618264 298066 618316
rect 260098 617516 260104 617568
rect 260156 617556 260162 617568
rect 282178 617556 282184 617568
rect 260156 617528 282184 617556
rect 260156 617516 260162 617528
rect 282178 617516 282184 617528
rect 282236 617516 282242 617568
rect 540422 617516 540428 617568
rect 540480 617556 540486 617568
rect 580166 617556 580172 617568
rect 540480 617528 580172 617556
rect 540480 617516 540486 617528
rect 580166 617516 580172 617528
rect 580224 617516 580230 617568
rect 293218 616836 293224 616888
rect 293276 616876 293282 616888
rect 298002 616876 298008 616888
rect 293276 616848 298008 616876
rect 293276 616836 293282 616848
rect 298002 616836 298008 616848
rect 298060 616836 298066 616888
rect 542906 616836 542912 616888
rect 542964 616876 542970 616888
rect 545574 616876 545580 616888
rect 542964 616848 545580 616876
rect 542964 616836 542970 616848
rect 545574 616836 545580 616848
rect 545632 616836 545638 616888
rect 159358 613368 159364 613420
rect 159416 613408 159422 613420
rect 171962 613408 171968 613420
rect 159416 613380 171968 613408
rect 159416 613368 159422 613380
rect 171962 613368 171968 613380
rect 172020 613368 172026 613420
rect 292022 612688 292028 612740
rect 292080 612728 292086 612740
rect 298002 612728 298008 612740
rect 292080 612700 298008 612728
rect 292080 612688 292086 612700
rect 298002 612688 298008 612700
rect 298060 612688 298066 612740
rect 398098 612008 398104 612060
rect 398156 612048 398162 612060
rect 410610 612048 410616 612060
rect 398156 612020 410616 612048
rect 398156 612008 398162 612020
rect 410610 612008 410616 612020
rect 410668 612008 410674 612060
rect 142890 611328 142896 611380
rect 142948 611368 142954 611380
rect 144270 611368 144276 611380
rect 142948 611340 144276 611368
rect 142948 611328 142954 611340
rect 144270 611328 144276 611340
rect 144328 611328 144334 611380
rect 175182 610648 175188 610700
rect 175240 610688 175246 610700
rect 179046 610688 179052 610700
rect 175240 610660 179052 610688
rect 175240 610648 175246 610660
rect 179046 610648 179052 610660
rect 179104 610648 179110 610700
rect 406470 610580 406476 610632
rect 406528 610620 406534 610632
rect 420178 610620 420184 610632
rect 406528 610592 420184 610620
rect 406528 610580 406534 610592
rect 420178 610580 420184 610592
rect 420236 610580 420242 610632
rect 377030 604528 377036 604580
rect 377088 604568 377094 604580
rect 379790 604568 379796 604580
rect 377088 604540 379796 604568
rect 377088 604528 377094 604540
rect 379790 604528 379796 604540
rect 379848 604528 379854 604580
rect 378042 604460 378048 604512
rect 378100 604500 378106 604512
rect 386414 604500 386420 604512
rect 378100 604472 386420 604500
rect 378100 604460 378106 604472
rect 386414 604460 386420 604472
rect 386472 604460 386478 604512
rect 410610 604460 410616 604512
rect 410668 604500 410674 604512
rect 413278 604500 413284 604512
rect 410668 604472 413284 604500
rect 410668 604460 410674 604472
rect 413278 604460 413284 604472
rect 413336 604460 413342 604512
rect 540330 604460 540336 604512
rect 540388 604500 540394 604512
rect 541434 604500 541440 604512
rect 540388 604472 541440 604500
rect 540388 604460 540394 604472
rect 541434 604460 541440 604472
rect 541492 604460 541498 604512
rect 286318 603100 286324 603152
rect 286376 603140 286382 603152
rect 297910 603140 297916 603152
rect 286376 603112 297916 603140
rect 286376 603100 286382 603112
rect 297910 603100 297916 603112
rect 297968 603100 297974 603152
rect 136082 602352 136088 602404
rect 136140 602392 136146 602404
rect 159358 602392 159364 602404
rect 136140 602364 159364 602392
rect 136140 602352 136146 602364
rect 159358 602352 159364 602364
rect 159416 602352 159422 602404
rect 539226 600992 539232 601044
rect 539284 601032 539290 601044
rect 540974 601032 540980 601044
rect 539284 601004 540980 601032
rect 539284 600992 539290 601004
rect 540974 600992 540980 601004
rect 541032 600992 541038 601044
rect 488350 600244 488356 600296
rect 488408 600284 488414 600296
rect 498838 600284 498844 600296
rect 488408 600256 498844 600284
rect 488408 600244 488414 600256
rect 498838 600244 498844 600256
rect 498896 600244 498902 600296
rect 537570 600244 537576 600296
rect 537628 600284 537634 600296
rect 540422 600284 540428 600296
rect 537628 600256 540428 600284
rect 537628 600244 537634 600256
rect 540422 600244 540428 600256
rect 540480 600244 540486 600296
rect 488258 600176 488264 600228
rect 488316 600216 488322 600228
rect 510338 600216 510344 600228
rect 488316 600188 510344 600216
rect 488316 600176 488322 600188
rect 510338 600176 510344 600188
rect 510396 600176 510402 600228
rect 488442 600108 488448 600160
rect 488500 600148 488506 600160
rect 524046 600148 524052 600160
rect 488500 600120 524052 600148
rect 488500 600108 488506 600120
rect 524046 600108 524052 600120
rect 524104 600108 524110 600160
rect 489638 600040 489644 600092
rect 489696 600080 489702 600092
rect 525886 600080 525892 600092
rect 489696 600052 525892 600080
rect 489696 600040 489702 600052
rect 525886 600040 525892 600052
rect 525944 600040 525950 600092
rect 462314 599972 462320 600024
rect 462372 600012 462378 600024
rect 499390 600012 499396 600024
rect 462372 599984 499396 600012
rect 462372 599972 462378 599984
rect 499390 599972 499396 599984
rect 499448 599972 499454 600024
rect 485682 599904 485688 599956
rect 485740 599944 485746 599956
rect 529198 599944 529204 599956
rect 485740 599916 529204 599944
rect 485740 599904 485746 599916
rect 529198 599904 529204 599916
rect 529256 599904 529262 599956
rect 486970 599836 486976 599888
rect 487028 599876 487034 599888
rect 530578 599876 530584 599888
rect 487028 599848 530584 599876
rect 487028 599836 487034 599848
rect 530578 599836 530584 599848
rect 530636 599836 530642 599888
rect 485590 599768 485596 599820
rect 485648 599808 485654 599820
rect 531406 599808 531412 599820
rect 485648 599780 531412 599808
rect 485648 599768 485654 599780
rect 531406 599768 531412 599780
rect 531464 599768 531470 599820
rect 486878 599700 486884 599752
rect 486936 599740 486942 599752
rect 532786 599740 532792 599752
rect 486936 599712 532792 599740
rect 486936 599700 486942 599712
rect 532786 599700 532792 599712
rect 532844 599700 532850 599752
rect 489730 599632 489736 599684
rect 489788 599672 489794 599684
rect 535730 599672 535736 599684
rect 489788 599644 535736 599672
rect 489788 599632 489794 599644
rect 535730 599632 535736 599644
rect 535788 599632 535794 599684
rect 413646 599564 413652 599616
rect 413704 599604 413710 599616
rect 499298 599604 499304 599616
rect 413704 599576 499304 599604
rect 413704 599564 413710 599576
rect 499298 599564 499304 599576
rect 499356 599564 499362 599616
rect 519722 598884 519728 598936
rect 519780 598924 519786 598936
rect 532970 598924 532976 598936
rect 519780 598896 532976 598924
rect 519780 598884 519786 598896
rect 532970 598884 532976 598896
rect 533028 598884 533034 598936
rect 515582 598816 515588 598868
rect 515640 598856 515646 598868
rect 529842 598856 529848 598868
rect 515640 598828 529848 598856
rect 515640 598816 515646 598828
rect 529842 598816 529848 598828
rect 529900 598816 529906 598868
rect 518342 598748 518348 598800
rect 518400 598788 518406 598800
rect 531314 598788 531320 598800
rect 518400 598760 531320 598788
rect 518400 598748 518406 598760
rect 531314 598748 531320 598760
rect 531372 598748 531378 598800
rect 512822 598272 512828 598324
rect 512880 598312 512886 598324
rect 527266 598312 527272 598324
rect 512880 598284 527272 598312
rect 512880 598272 512886 598284
rect 527266 598272 527272 598284
rect 527324 598272 527330 598324
rect 493502 598204 493508 598256
rect 493560 598244 493566 598256
rect 498930 598244 498936 598256
rect 493560 598216 498936 598244
rect 493560 598204 493566 598216
rect 498930 598204 498936 598216
rect 498988 598204 498994 598256
rect 514202 598204 514208 598256
rect 514260 598244 514266 598256
rect 535546 598244 535552 598256
rect 514260 598216 535552 598244
rect 514260 598204 514266 598216
rect 535546 598204 535552 598216
rect 535604 598204 535610 598256
rect 492122 598136 492128 598188
rect 492180 598176 492186 598188
rect 498746 598176 498752 598188
rect 492180 598148 498752 598176
rect 492180 598136 492186 598148
rect 498746 598136 498752 598148
rect 498804 598136 498810 598188
rect 531222 598136 531228 598188
rect 531280 598176 531286 598188
rect 536282 598176 536288 598188
rect 531280 598148 536288 598176
rect 531280 598136 531286 598148
rect 536282 598136 536288 598148
rect 536340 598136 536346 598188
rect 496262 598068 496268 598120
rect 496320 598108 496326 598120
rect 499114 598108 499120 598120
rect 496320 598080 499120 598108
rect 496320 598068 496326 598080
rect 499114 598068 499120 598080
rect 499172 598068 499178 598120
rect 518158 597524 518164 597576
rect 518216 597564 518222 597576
rect 521102 597564 521108 597576
rect 518216 597536 521108 597564
rect 518216 597524 518222 597536
rect 521102 597524 521108 597536
rect 521160 597524 521166 597576
rect 536098 597524 536104 597576
rect 536156 597564 536162 597576
rect 539042 597564 539048 597576
rect 536156 597536 539048 597564
rect 536156 597524 536162 597536
rect 539042 597524 539048 597536
rect 539100 597524 539106 597576
rect 378042 593444 378048 593496
rect 378100 593484 378106 593496
rect 385034 593484 385040 593496
rect 378100 593456 385040 593484
rect 378100 593444 378106 593456
rect 385034 593444 385040 593456
rect 385092 593444 385098 593496
rect 377950 593376 377956 593428
rect 378008 593416 378014 593428
rect 386598 593416 386604 593428
rect 378008 593388 386604 593416
rect 378008 593376 378014 593388
rect 386598 593376 386604 593388
rect 386656 593376 386662 593428
rect 141418 593308 141424 593360
rect 141476 593348 141482 593360
rect 142890 593348 142896 593360
rect 141476 593320 142896 593348
rect 141476 593308 141482 593320
rect 142890 593308 142896 593320
rect 142948 593308 142954 593360
rect 378042 592288 378048 592340
rect 378100 592328 378106 592340
rect 382826 592328 382832 592340
rect 378100 592300 382832 592328
rect 378100 592288 378106 592300
rect 382826 592288 382832 592300
rect 382884 592288 382890 592340
rect 378042 592084 378048 592136
rect 378100 592124 378106 592136
rect 385310 592124 385316 592136
rect 378100 592096 385316 592124
rect 378100 592084 378106 592096
rect 385310 592084 385316 592096
rect 385368 592084 385374 592136
rect 45278 592016 45284 592068
rect 45336 592056 45342 592068
rect 57514 592056 57520 592068
rect 45336 592028 57520 592056
rect 45336 592016 45342 592028
rect 57514 592016 57520 592028
rect 57572 592016 57578 592068
rect 134518 591336 134524 591388
rect 134576 591376 134582 591388
rect 136082 591376 136088 591388
rect 134576 591348 136088 591376
rect 134576 591336 134582 591348
rect 136082 591336 136088 591348
rect 136140 591336 136146 591388
rect 378042 590656 378048 590708
rect 378100 590696 378106 590708
rect 385218 590696 385224 590708
rect 378100 590668 385224 590696
rect 378100 590656 378106 590668
rect 385218 590656 385224 590668
rect 385276 590656 385282 590708
rect 378042 589908 378048 589960
rect 378100 589948 378106 589960
rect 385402 589948 385408 589960
rect 378100 589920 385408 589948
rect 378100 589908 378106 589920
rect 385402 589908 385408 589920
rect 385460 589908 385466 589960
rect 420178 589908 420184 589960
rect 420236 589948 420242 589960
rect 428458 589948 428464 589960
rect 420236 589920 428464 589948
rect 420236 589908 420242 589920
rect 428458 589908 428464 589920
rect 428516 589908 428522 589960
rect 378042 589296 378048 589348
rect 378100 589336 378106 589348
rect 382458 589336 382464 589348
rect 378100 589308 382464 589336
rect 378100 589296 378106 589308
rect 382458 589296 382464 589308
rect 382516 589296 382522 589348
rect 378042 587936 378048 587988
rect 378100 587976 378106 587988
rect 382274 587976 382280 587988
rect 378100 587948 382280 587976
rect 378100 587936 378106 587948
rect 382274 587936 382280 587948
rect 382332 587936 382338 587988
rect 376938 587868 376944 587920
rect 376996 587908 377002 587920
rect 379606 587908 379612 587920
rect 376996 587880 379612 587908
rect 376996 587868 377002 587880
rect 379606 587868 379612 587880
rect 379664 587868 379670 587920
rect 413278 587800 413284 587852
rect 413336 587840 413342 587852
rect 416130 587840 416136 587852
rect 413336 587812 416136 587840
rect 413336 587800 413342 587812
rect 416130 587800 416136 587812
rect 416188 587800 416194 587852
rect 377766 586916 377772 586968
rect 377824 586956 377830 586968
rect 381262 586956 381268 586968
rect 377824 586928 381268 586956
rect 377824 586916 377830 586928
rect 381262 586916 381268 586928
rect 381320 586916 381326 586968
rect 162302 586576 162308 586628
rect 162360 586616 162366 586628
rect 170858 586616 170864 586628
rect 162360 586588 170864 586616
rect 162360 586576 162366 586588
rect 170858 586576 170864 586588
rect 170916 586576 170922 586628
rect 378042 586576 378048 586628
rect 378100 586616 378106 586628
rect 383746 586616 383752 586628
rect 378100 586588 383752 586616
rect 378100 586576 378106 586588
rect 383746 586576 383752 586588
rect 383804 586576 383810 586628
rect 141510 586508 141516 586560
rect 141568 586548 141574 586560
rect 142798 586548 142804 586560
rect 141568 586520 142804 586548
rect 141568 586508 141574 586520
rect 142798 586508 142804 586520
rect 142856 586508 142862 586560
rect 162578 586508 162584 586560
rect 162636 586548 162642 586560
rect 169478 586548 169484 586560
rect 162636 586520 169484 586548
rect 162636 586508 162642 586520
rect 169478 586508 169484 586520
rect 169536 586508 169542 586560
rect 378042 585148 378048 585200
rect 378100 585188 378106 585200
rect 382366 585188 382372 585200
rect 378100 585160 382372 585188
rect 378100 585148 378106 585160
rect 382366 585148 382372 585160
rect 382424 585148 382430 585200
rect 258718 584400 258724 584452
rect 258776 584440 258782 584452
rect 258902 584440 258908 584452
rect 258776 584412 258908 584440
rect 258776 584400 258782 584412
rect 258902 584400 258908 584412
rect 258960 584400 258966 584452
rect 378042 584128 378048 584180
rect 378100 584168 378106 584180
rect 383654 584168 383660 584180
rect 378100 584140 383660 584168
rect 378100 584128 378106 584140
rect 383654 584128 383660 584140
rect 383712 584128 383718 584180
rect 140038 583720 140044 583772
rect 140096 583760 140102 583772
rect 141510 583760 141516 583772
rect 140096 583732 141516 583760
rect 140096 583720 140102 583732
rect 141510 583720 141516 583732
rect 141568 583720 141574 583772
rect 378042 583720 378048 583772
rect 378100 583760 378106 583772
rect 382734 583760 382740 583772
rect 378100 583732 382740 583760
rect 378100 583720 378106 583732
rect 382734 583720 382740 583732
rect 382792 583720 382798 583772
rect 378042 582496 378048 582548
rect 378100 582536 378106 582548
rect 382642 582536 382648 582548
rect 378100 582508 382648 582536
rect 378100 582496 378106 582508
rect 382642 582496 382648 582508
rect 382700 582496 382706 582548
rect 378042 582360 378048 582412
rect 378100 582400 378106 582412
rect 382550 582400 382556 582412
rect 378100 582372 382556 582400
rect 378100 582360 378106 582372
rect 382550 582360 382556 582372
rect 382608 582360 382614 582412
rect 490374 581612 490380 581664
rect 490432 581652 490438 581664
rect 493318 581652 493324 581664
rect 490432 581624 493324 581652
rect 490432 581612 490438 581624
rect 493318 581612 493324 581624
rect 493376 581612 493382 581664
rect 377858 581000 377864 581052
rect 377916 581040 377922 581052
rect 381446 581040 381452 581052
rect 377916 581012 381452 581040
rect 377916 581000 377922 581012
rect 381446 581000 381452 581012
rect 381504 581000 381510 581052
rect 165062 579776 165068 579828
rect 165120 579816 165126 579828
rect 173710 579816 173716 579828
rect 165120 579788 173716 579816
rect 165120 579776 165126 579788
rect 173710 579776 173716 579788
rect 173768 579776 173774 579828
rect 377582 579708 377588 579760
rect 377640 579748 377646 579760
rect 380894 579748 380900 579760
rect 377640 579720 380900 579748
rect 377640 579708 377646 579720
rect 380894 579708 380900 579720
rect 380952 579708 380958 579760
rect 3418 579640 3424 579692
rect 3476 579680 3482 579692
rect 41506 579680 41512 579692
rect 3476 579652 41512 579680
rect 3476 579640 3482 579652
rect 41506 579640 41512 579652
rect 41564 579640 41570 579692
rect 377122 579640 377128 579692
rect 377180 579680 377186 579692
rect 379882 579680 379888 579692
rect 377180 579652 379888 579680
rect 377180 579640 377186 579652
rect 379882 579640 379888 579652
rect 379940 579640 379946 579692
rect 377858 578280 377864 578332
rect 377916 578320 377922 578332
rect 381354 578320 381360 578332
rect 377916 578292 381360 578320
rect 377916 578280 377922 578292
rect 381354 578280 381360 578292
rect 381412 578280 381418 578332
rect 377030 578212 377036 578264
rect 377088 578252 377094 578264
rect 379698 578252 379704 578264
rect 377088 578224 379704 578252
rect 377088 578212 377094 578224
rect 379698 578212 379704 578224
rect 379756 578212 379762 578264
rect 377122 575492 377128 575544
rect 377180 575532 377186 575544
rect 379974 575532 379980 575544
rect 377180 575504 379980 575532
rect 377180 575492 377186 575504
rect 379974 575492 379980 575504
rect 380032 575492 380038 575544
rect 416130 575492 416136 575544
rect 416188 575532 416194 575544
rect 419626 575532 419632 575544
rect 416188 575504 419632 575532
rect 416188 575492 416194 575504
rect 419626 575492 419632 575504
rect 419684 575492 419690 575544
rect 378042 572704 378048 572756
rect 378100 572744 378106 572756
rect 386690 572744 386696 572756
rect 378100 572716 386696 572744
rect 378100 572704 378106 572716
rect 386690 572704 386696 572716
rect 386748 572704 386754 572756
rect 378042 571888 378048 571940
rect 378100 571928 378106 571940
rect 383838 571928 383844 571940
rect 378100 571900 383844 571928
rect 378100 571888 378106 571900
rect 383838 571888 383844 571900
rect 383896 571888 383902 571940
rect 378042 571344 378048 571396
rect 378100 571384 378106 571396
rect 383930 571384 383936 571396
rect 378100 571356 383936 571384
rect 378100 571344 378106 571356
rect 383930 571344 383936 571356
rect 383988 571344 383994 571396
rect 428458 571276 428464 571328
rect 428516 571316 428522 571328
rect 433978 571316 433984 571328
rect 428516 571288 433984 571316
rect 428516 571276 428522 571288
rect 433978 571276 433984 571288
rect 434036 571276 434042 571328
rect 419626 570596 419632 570648
rect 419684 570636 419690 570648
rect 429194 570636 429200 570648
rect 419684 570608 429200 570636
rect 419684 570596 419690 570608
rect 429194 570596 429200 570608
rect 429252 570596 429258 570648
rect 169294 569780 169300 569832
rect 169352 569820 169358 569832
rect 171134 569820 171140 569832
rect 169352 569792 171140 569820
rect 169352 569780 169358 569792
rect 171134 569780 171140 569792
rect 171192 569780 171198 569832
rect 164970 569644 164976 569696
rect 165028 569684 165034 569696
rect 172422 569684 172428 569696
rect 165028 569656 172428 569684
rect 165028 569644 165034 569656
rect 172422 569644 172428 569656
rect 172480 569644 172486 569696
rect 377030 568556 377036 568608
rect 377088 568596 377094 568608
rect 379514 568596 379520 568608
rect 377088 568568 379520 568596
rect 377088 568556 377094 568568
rect 379514 568556 379520 568568
rect 379572 568556 379578 568608
rect 493318 568488 493324 568540
rect 493376 568528 493382 568540
rect 496078 568528 496084 568540
rect 493376 568500 496084 568528
rect 493376 568488 493382 568500
rect 496078 568488 496084 568500
rect 496136 568488 496142 568540
rect 377766 567808 377772 567860
rect 377824 567848 377830 567860
rect 381170 567848 381176 567860
rect 377824 567820 381176 567848
rect 377824 567808 377830 567820
rect 381170 567808 381176 567820
rect 381228 567808 381234 567860
rect 429194 567196 429200 567248
rect 429252 567236 429258 567248
rect 432046 567236 432052 567248
rect 429252 567208 432052 567236
rect 429252 567196 429258 567208
rect 432046 567196 432052 567208
rect 432104 567196 432110 567248
rect 543734 564340 543740 564392
rect 543792 564380 543798 564392
rect 580166 564380 580172 564392
rect 543792 564352 580172 564380
rect 543792 564340 543798 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 537754 563660 537760 563712
rect 537812 563700 537818 563712
rect 543734 563700 543740 563712
rect 537812 563672 543740 563700
rect 537812 563660 537818 563672
rect 543734 563660 543740 563672
rect 543792 563660 543798 563712
rect 169110 562300 169116 562352
rect 169168 562340 169174 562352
rect 170122 562340 170128 562352
rect 169168 562312 170128 562340
rect 169168 562300 169174 562312
rect 170122 562300 170128 562312
rect 170180 562300 170186 562352
rect 178402 562300 178408 562352
rect 178460 562340 178466 562352
rect 178678 562340 178684 562352
rect 178460 562312 178684 562340
rect 178460 562300 178466 562312
rect 178678 562300 178684 562312
rect 178736 562300 178742 562352
rect 432046 562300 432052 562352
rect 432104 562340 432110 562352
rect 444282 562340 444288 562352
rect 432104 562312 444288 562340
rect 432104 562300 432110 562312
rect 444282 562300 444288 562312
rect 444340 562300 444346 562352
rect 140038 561824 140044 561876
rect 140096 561824 140102 561876
rect 140056 561728 140084 561824
rect 138032 561700 140084 561728
rect 135162 561620 135168 561672
rect 135220 561660 135226 561672
rect 138032 561660 138060 561700
rect 259178 561688 259184 561740
rect 259236 561728 259242 561740
rect 299658 561728 299664 561740
rect 259236 561700 299664 561728
rect 259236 561688 259242 561700
rect 299658 561688 299664 561700
rect 299716 561688 299722 561740
rect 135220 561632 138060 561660
rect 135220 561620 135226 561632
rect 310486 561224 313274 561252
rect 299566 561144 299572 561196
rect 299624 561184 299630 561196
rect 310486 561184 310514 561224
rect 299624 561156 310514 561184
rect 313246 561184 313274 561224
rect 313246 561156 314654 561184
rect 299624 561144 299630 561156
rect 314626 561116 314654 561156
rect 314626 561088 316034 561116
rect 254486 561008 254492 561060
rect 254544 561048 254550 561060
rect 316006 561048 316034 561088
rect 254544 561020 309134 561048
rect 316006 561020 317414 561048
rect 254544 561008 254550 561020
rect 299566 560980 299572 560992
rect 253584 560952 299572 560980
rect 253584 560652 253612 560952
rect 299566 560940 299572 560952
rect 299624 560940 299630 560992
rect 294046 560872 294052 560924
rect 294104 560912 294110 560924
rect 297910 560912 297916 560924
rect 294104 560884 297916 560912
rect 294104 560872 294110 560884
rect 297910 560872 297916 560884
rect 297968 560872 297974 560924
rect 309106 560776 309134 561020
rect 317386 560980 317414 561020
rect 525978 560980 525984 560992
rect 317386 560952 525984 560980
rect 525978 560940 525984 560952
rect 526036 560940 526042 560992
rect 316006 560884 318794 560912
rect 316006 560844 316034 560884
rect 311866 560816 316034 560844
rect 311866 560776 311894 560816
rect 309106 560748 311894 560776
rect 254670 560668 254676 560720
rect 254728 560708 254734 560720
rect 293954 560708 293960 560720
rect 254728 560680 293960 560708
rect 254728 560668 254734 560680
rect 293954 560668 293960 560680
rect 294012 560668 294018 560720
rect 253566 560600 253572 560652
rect 253624 560600 253630 560652
rect 254854 560600 254860 560652
rect 254912 560640 254918 560652
rect 318766 560640 318794 560884
rect 319346 560640 319352 560652
rect 254912 560612 300808 560640
rect 318766 560612 319352 560640
rect 254912 560600 254918 560612
rect 254394 560532 254400 560584
rect 254452 560572 254458 560584
rect 300578 560572 300584 560584
rect 254452 560544 300584 560572
rect 254452 560532 254458 560544
rect 300578 560532 300584 560544
rect 300636 560532 300642 560584
rect 253474 560464 253480 560516
rect 253532 560504 253538 560516
rect 300670 560504 300676 560516
rect 253532 560476 300676 560504
rect 253532 560464 253538 560476
rect 300670 560464 300676 560476
rect 300728 560464 300734 560516
rect 246574 560396 246580 560448
rect 246632 560436 246638 560448
rect 299566 560436 299572 560448
rect 246632 560408 299572 560436
rect 246632 560396 246638 560408
rect 299566 560396 299572 560408
rect 299624 560396 299630 560448
rect 169202 560328 169208 560380
rect 169260 560368 169266 560380
rect 172238 560368 172244 560380
rect 169260 560340 172244 560368
rect 169260 560328 169266 560340
rect 172238 560328 172244 560340
rect 172296 560328 172302 560380
rect 300780 560368 300808 560612
rect 319346 560600 319352 560612
rect 319404 560600 319410 560652
rect 300780 560340 300900 560368
rect 59538 560260 59544 560312
rect 59596 560300 59602 560312
rect 60734 560300 60740 560312
rect 59596 560272 60740 560300
rect 59596 560260 59602 560272
rect 60734 560260 60740 560272
rect 60792 560260 60798 560312
rect 179046 560260 179052 560312
rect 179104 560300 179110 560312
rect 245470 560300 245476 560312
rect 179104 560272 245476 560300
rect 179104 560260 179110 560272
rect 245470 560260 245476 560272
rect 245528 560260 245534 560312
rect 287790 560260 287796 560312
rect 287848 560300 287854 560312
rect 287848 560272 300808 560300
rect 287848 560260 287854 560272
rect 45278 560192 45284 560244
rect 45336 560232 45342 560244
rect 162486 560232 162492 560244
rect 45336 560204 162492 560232
rect 45336 560192 45342 560204
rect 162486 560192 162492 560204
rect 162544 560192 162550 560244
rect 168006 560192 168012 560244
rect 168064 560232 168070 560244
rect 172330 560232 172336 560244
rect 168064 560204 172336 560232
rect 168064 560192 168070 560204
rect 172330 560192 172336 560204
rect 172388 560192 172394 560244
rect 175734 560192 175740 560244
rect 175792 560232 175798 560244
rect 297634 560232 297640 560244
rect 175792 560204 297640 560232
rect 175792 560192 175798 560204
rect 297634 560192 297640 560204
rect 297692 560192 297698 560244
rect 300780 560164 300808 560272
rect 300872 560232 300900 560340
rect 315390 560232 315396 560244
rect 300872 560204 315396 560232
rect 315390 560192 315396 560204
rect 315448 560192 315454 560244
rect 318334 560164 318340 560176
rect 300780 560136 318340 560164
rect 318334 560124 318340 560136
rect 318392 560124 318398 560176
rect 165522 560056 165528 560108
rect 165580 560096 165586 560108
rect 173710 560096 173716 560108
rect 165580 560068 173716 560096
rect 165580 560056 165586 560068
rect 173710 560056 173716 560068
rect 173768 560056 173774 560108
rect 299658 560056 299664 560108
rect 299716 560096 299722 560108
rect 306374 560096 306380 560108
rect 299716 560068 306380 560096
rect 299716 560056 299722 560068
rect 306374 560056 306380 560068
rect 306432 560056 306438 560108
rect 216674 559580 216680 559632
rect 216732 559620 216738 559632
rect 357802 559620 357808 559632
rect 216732 559592 357808 559620
rect 216732 559580 216738 559592
rect 357802 559580 357808 559592
rect 357860 559580 357866 559632
rect 444282 559580 444288 559632
rect 444340 559620 444346 559632
rect 459094 559620 459100 559632
rect 444340 559592 459100 559620
rect 444340 559580 444346 559592
rect 459094 559580 459100 559592
rect 459152 559580 459158 559632
rect 91186 559512 91192 559564
rect 91244 559552 91250 559564
rect 141418 559552 141424 559564
rect 91244 559524 141424 559552
rect 91244 559512 91250 559524
rect 141418 559512 141424 559524
rect 141476 559512 141482 559564
rect 177206 559512 177212 559564
rect 177264 559552 177270 559564
rect 514846 559552 514852 559564
rect 177264 559524 514852 559552
rect 177264 559512 177270 559524
rect 514846 559512 514852 559524
rect 514904 559512 514910 559564
rect 169846 559444 169852 559496
rect 169904 559484 169910 559496
rect 367922 559484 367928 559496
rect 169904 559456 367928 559484
rect 169904 559444 169910 559456
rect 367922 559444 367928 559456
rect 367980 559444 367986 559496
rect 169754 559376 169760 559428
rect 169812 559416 169818 559428
rect 368934 559416 368940 559428
rect 169812 559388 368940 559416
rect 169812 559376 169818 559388
rect 368934 559376 368940 559388
rect 368992 559376 368998 559428
rect 233694 559308 233700 559360
rect 233752 559348 233758 559360
rect 500218 559348 500224 559360
rect 233752 559320 500224 559348
rect 233752 559308 233758 559320
rect 500218 559308 500224 559320
rect 500276 559308 500282 559360
rect 60642 559240 60648 559292
rect 60700 559280 60706 559292
rect 369946 559280 369952 559292
rect 60700 559252 369952 559280
rect 60700 559240 60706 559252
rect 369946 559240 369952 559252
rect 370004 559240 370010 559292
rect 57238 559172 57244 559224
rect 57296 559212 57302 559224
rect 370958 559212 370964 559224
rect 57296 559184 370964 559212
rect 57296 559172 57302 559184
rect 370958 559172 370964 559184
rect 371016 559172 371022 559224
rect 56962 559104 56968 559156
rect 57020 559144 57026 559156
rect 371970 559144 371976 559156
rect 57020 559116 371976 559144
rect 57020 559104 57026 559116
rect 371970 559104 371976 559116
rect 372028 559104 372034 559156
rect 57514 559036 57520 559088
rect 57572 559076 57578 559088
rect 373258 559076 373264 559088
rect 57572 559048 373264 559076
rect 57572 559036 57578 559048
rect 373258 559036 373264 559048
rect 373316 559036 373322 559088
rect 166534 558968 166540 559020
rect 166592 559008 166598 559020
rect 511994 559008 512000 559020
rect 166592 558980 512000 559008
rect 166592 558968 166598 558980
rect 511994 558968 512000 558980
rect 512052 558968 512058 559020
rect 166810 558900 166816 558952
rect 166868 558940 166874 558952
rect 520734 558940 520740 558952
rect 166868 558912 520740 558940
rect 166868 558900 166874 558912
rect 520734 558900 520740 558912
rect 520792 558900 520798 558952
rect 53834 558832 53840 558884
rect 53892 558872 53898 558884
rect 372338 558872 372344 558884
rect 53892 558844 372344 558872
rect 53892 558832 53898 558844
rect 372338 558832 372344 558844
rect 372396 558832 372402 558884
rect 53926 558764 53932 558816
rect 53984 558804 53990 558816
rect 367278 558804 367284 558816
rect 53984 558776 367284 558804
rect 53984 558764 53990 558776
rect 367278 558764 367284 558776
rect 367336 558764 367342 558816
rect 56042 558696 56048 558748
rect 56100 558736 56106 558748
rect 361206 558736 361212 558748
rect 56100 558708 361212 558736
rect 56100 558696 56106 558708
rect 361206 558696 361212 558708
rect 361264 558696 361270 558748
rect 59262 558628 59268 558680
rect 59320 558668 59326 558680
rect 357158 558668 357164 558680
rect 59320 558640 357164 558668
rect 59320 558628 59326 558640
rect 357158 558628 357164 558640
rect 357216 558628 357222 558680
rect 63586 558560 63592 558612
rect 63644 558600 63650 558612
rect 355134 558600 355140 558612
rect 63644 558572 355140 558600
rect 63644 558560 63650 558572
rect 355134 558560 355140 558572
rect 355192 558560 355198 558612
rect 89622 558492 89628 558544
rect 89680 558532 89686 558544
rect 91186 558532 91192 558544
rect 89680 558504 91192 558532
rect 89680 558492 89686 558504
rect 91186 558492 91192 558504
rect 91244 558492 91250 558544
rect 231762 558492 231768 558544
rect 231820 558532 231826 558544
rect 297542 558532 297548 558544
rect 231820 558504 297548 558532
rect 231820 558492 231826 558504
rect 297542 558492 297548 558504
rect 297600 558492 297606 558544
rect 300670 558492 300676 558544
rect 300728 558532 300734 558544
rect 314654 558532 314660 558544
rect 300728 558504 314660 558532
rect 300728 558492 300734 558504
rect 314654 558492 314660 558504
rect 314712 558492 314718 558544
rect 245654 558424 245660 558476
rect 245712 558464 245718 558476
rect 245712 558436 277394 558464
rect 245712 558424 245718 558436
rect 199930 558288 199936 558340
rect 199988 558328 199994 558340
rect 251818 558328 251824 558340
rect 199988 558300 251824 558328
rect 199988 558288 199994 558300
rect 251818 558288 251824 558300
rect 251876 558288 251882 558340
rect 277366 558328 277394 558436
rect 293954 558424 293960 558476
rect 294012 558464 294018 558476
rect 353110 558464 353116 558476
rect 294012 558436 353116 558464
rect 294012 558424 294018 558436
rect 353110 558424 353116 558436
rect 353168 558424 353174 558476
rect 293310 558356 293316 558408
rect 293368 558396 293374 558408
rect 303522 558396 303528 558408
rect 293368 558368 303528 558396
rect 293368 558356 293374 558368
rect 303522 558356 303528 558368
rect 303580 558356 303586 558408
rect 294046 558328 294052 558340
rect 277366 558300 294052 558328
rect 294046 558288 294052 558300
rect 294104 558288 294110 558340
rect 300578 558288 300584 558340
rect 300636 558328 300642 558340
rect 521930 558328 521936 558340
rect 300636 558300 521936 558328
rect 300636 558288 300642 558300
rect 521930 558288 521936 558300
rect 521988 558288 521994 558340
rect 177298 558220 177304 558272
rect 177356 558260 177362 558272
rect 503990 558260 503996 558272
rect 177356 558232 503996 558260
rect 177356 558220 177362 558232
rect 503990 558220 503996 558232
rect 504048 558220 504054 558272
rect 104894 558152 104900 558204
rect 104952 558192 104958 558204
rect 135162 558192 135168 558204
rect 104952 558164 135168 558192
rect 104952 558152 104958 558164
rect 135162 558152 135168 558164
rect 135220 558152 135226 558204
rect 177574 558152 177580 558204
rect 177632 558192 177638 558204
rect 512178 558192 512184 558204
rect 177632 558164 512184 558192
rect 177632 558152 177638 558164
rect 512178 558152 512184 558164
rect 512236 558152 512242 558204
rect 252462 557676 252468 557728
rect 252520 557716 252526 557728
rect 346670 557716 346676 557728
rect 252520 557688 346676 557716
rect 252520 557676 252526 557688
rect 346670 557676 346676 557688
rect 346728 557676 346734 557728
rect 41506 557648 41512 557660
rect 41432 557620 41512 557648
rect 37090 557540 37096 557592
rect 37148 557580 37154 557592
rect 41432 557580 41460 557620
rect 41506 557608 41512 557620
rect 41564 557608 41570 557660
rect 180702 557608 180708 557660
rect 180760 557648 180766 557660
rect 524690 557648 524696 557660
rect 180760 557620 524696 557648
rect 180760 557608 180766 557620
rect 524690 557608 524696 557620
rect 524748 557608 524754 557660
rect 37148 557552 41460 557580
rect 37148 557540 37154 557552
rect 41432 557444 41460 557552
rect 180610 557540 180616 557592
rect 180668 557580 180674 557592
rect 537018 557580 537024 557592
rect 180668 557552 537024 557580
rect 180668 557540 180674 557552
rect 537018 557540 537024 557552
rect 537076 557540 537082 557592
rect 53834 557472 53840 557524
rect 53892 557512 53898 557524
rect 297726 557512 297732 557524
rect 53892 557484 297732 557512
rect 53892 557472 53898 557484
rect 297726 557472 297732 557484
rect 297784 557472 297790 557524
rect 156598 557444 156604 557456
rect 41432 557416 156604 557444
rect 156598 557404 156604 557416
rect 156656 557404 156662 557456
rect 202046 557404 202052 557456
rect 202104 557444 202110 557456
rect 254394 557444 254400 557456
rect 202104 557416 254400 557444
rect 202104 557404 202110 557416
rect 254394 557404 254400 557416
rect 254452 557404 254458 557456
rect 128262 557064 128268 557116
rect 128320 557104 128326 557116
rect 174906 557104 174912 557116
rect 128320 557076 174912 557104
rect 128320 557064 128326 557076
rect 174906 557064 174912 557076
rect 174964 557064 174970 557116
rect 57606 556996 57612 557048
rect 57664 557036 57670 557048
rect 170858 557036 170864 557048
rect 57664 557008 170864 557036
rect 57664 556996 57670 557008
rect 170858 556996 170864 557008
rect 170916 556996 170922 557048
rect 250438 556996 250444 557048
rect 250496 557036 250502 557048
rect 293218 557036 293224 557048
rect 250496 557008 293224 557036
rect 250496 556996 250502 557008
rect 293218 556996 293224 557008
rect 293276 556996 293282 557048
rect 137738 556928 137744 556980
rect 137796 556968 137802 556980
rect 258994 556968 259000 556980
rect 137796 556940 259000 556968
rect 137796 556928 137802 556940
rect 258994 556928 259000 556940
rect 259052 556928 259058 556980
rect 280798 556928 280804 556980
rect 280856 556968 280862 556980
rect 378778 556968 378784 556980
rect 280856 556940 378784 556968
rect 280856 556928 280862 556940
rect 378778 556928 378784 556940
rect 378836 556928 378842 556980
rect 91094 556860 91100 556912
rect 91152 556900 91158 556912
rect 104894 556900 104900 556912
rect 91152 556872 104900 556900
rect 91152 556860 91158 556872
rect 104894 556860 104900 556872
rect 104952 556860 104958 556912
rect 137922 556860 137928 556912
rect 137980 556900 137986 556912
rect 331950 556900 331956 556912
rect 137980 556872 331956 556900
rect 137980 556860 137986 556872
rect 331950 556860 331956 556872
rect 332008 556860 332014 556912
rect 61378 556792 61384 556844
rect 61436 556832 61442 556844
rect 375926 556832 375932 556844
rect 61436 556804 375932 556832
rect 61436 556792 61442 556804
rect 375926 556792 375932 556804
rect 375984 556792 375990 556844
rect 255038 556656 255044 556708
rect 255096 556696 255102 556708
rect 260098 556696 260104 556708
rect 255096 556668 260104 556696
rect 255096 556656 255102 556668
rect 260098 556656 260104 556668
rect 260156 556656 260162 556708
rect 230382 556588 230388 556640
rect 230440 556628 230446 556640
rect 448882 556628 448888 556640
rect 230440 556600 448888 556628
rect 230440 556588 230446 556600
rect 448882 556588 448888 556600
rect 448940 556588 448946 556640
rect 227714 556520 227720 556572
rect 227772 556560 227778 556572
rect 449894 556560 449900 556572
rect 227772 556532 449900 556560
rect 227772 556520 227778 556532
rect 449894 556520 449900 556532
rect 449952 556520 449958 556572
rect 179414 556452 179420 556504
rect 179472 556492 179478 556504
rect 450906 556492 450912 556504
rect 179472 556464 450912 556492
rect 179472 556452 179478 556464
rect 450906 556452 450912 556464
rect 450964 556452 450970 556504
rect 178126 556384 178132 556436
rect 178184 556424 178190 556436
rect 452930 556424 452936 556436
rect 178184 556396 452936 556424
rect 178184 556384 178190 556396
rect 452930 556384 452936 556396
rect 452988 556384 452994 556436
rect 178034 556316 178040 556368
rect 178092 556356 178098 556368
rect 453942 556356 453948 556368
rect 178092 556328 453948 556356
rect 178092 556316 178098 556328
rect 453942 556316 453948 556328
rect 454000 556316 454006 556368
rect 137462 556248 137468 556300
rect 137520 556288 137526 556300
rect 137738 556288 137744 556300
rect 137520 556260 137744 556288
rect 137520 556248 137526 556260
rect 137738 556248 137744 556260
rect 137796 556248 137802 556300
rect 175826 556248 175832 556300
rect 175884 556288 175890 556300
rect 454954 556288 454960 556300
rect 175884 556260 454960 556288
rect 175884 556248 175890 556260
rect 454954 556248 454960 556260
rect 455012 556248 455018 556300
rect 56042 556180 56048 556232
rect 56100 556220 56106 556232
rect 56502 556220 56508 556232
rect 56100 556192 56508 556220
rect 56100 556180 56106 556192
rect 56502 556180 56508 556192
rect 56560 556180 56566 556232
rect 86862 556180 86868 556232
rect 86920 556220 86926 556232
rect 89622 556220 89628 556232
rect 86920 556192 89628 556220
rect 86920 556180 86926 556192
rect 89622 556180 89628 556192
rect 89680 556180 89686 556232
rect 175182 556180 175188 556232
rect 175240 556220 175246 556232
rect 509970 556220 509976 556232
rect 175240 556192 509976 556220
rect 175240 556180 175246 556192
rect 509970 556180 509976 556192
rect 510028 556180 510034 556232
rect 137186 556112 137192 556164
rect 137244 556152 137250 556164
rect 137462 556152 137468 556164
rect 137244 556124 137468 556152
rect 137244 556112 137250 556124
rect 137462 556112 137468 556124
rect 137520 556112 137526 556164
rect 56502 556044 56508 556096
rect 56560 556084 56566 556096
rect 379974 556084 379980 556096
rect 56560 556056 379980 556084
rect 56560 556044 56566 556056
rect 379974 556044 379980 556056
rect 380032 556044 380038 556096
rect 137186 555976 137192 556028
rect 137244 556016 137250 556028
rect 376938 556016 376944 556028
rect 137244 555988 376944 556016
rect 137244 555976 137250 555988
rect 376938 555976 376944 555988
rect 376996 555976 377002 556028
rect 53834 555908 53840 555960
rect 53892 555948 53898 555960
rect 381446 555948 381452 555960
rect 53892 555920 381452 555948
rect 53892 555908 53898 555920
rect 381446 555908 381452 555920
rect 381504 555908 381510 555960
rect 137462 555568 137468 555620
rect 137520 555608 137526 555620
rect 271138 555608 271144 555620
rect 137520 555580 271144 555608
rect 137520 555568 137526 555580
rect 271138 555568 271144 555580
rect 271196 555568 271202 555620
rect 137646 555500 137652 555552
rect 137704 555540 137710 555552
rect 347130 555540 347136 555552
rect 137704 555512 347136 555540
rect 137704 555500 137710 555512
rect 347130 555500 347136 555512
rect 347188 555500 347194 555552
rect 175826 555432 175832 555484
rect 175884 555472 175890 555484
rect 507854 555472 507860 555484
rect 175884 555444 507860 555472
rect 175884 555432 175890 555444
rect 507854 555432 507860 555444
rect 507912 555432 507918 555484
rect 247034 555160 247040 555212
rect 247092 555200 247098 555212
rect 434714 555200 434720 555212
rect 247092 555172 434720 555200
rect 247092 555160 247098 555172
rect 434714 555160 434720 555172
rect 434772 555160 434778 555212
rect 226334 555092 226340 555144
rect 226392 555132 226398 555144
rect 460014 555132 460020 555144
rect 226392 555104 460020 555132
rect 226392 555092 226398 555104
rect 460014 555092 460020 555104
rect 460072 555092 460078 555144
rect 179414 555024 179420 555076
rect 179472 555064 179478 555076
rect 473170 555064 473176 555076
rect 179472 555036 473176 555064
rect 179472 555024 179478 555036
rect 473170 555024 473176 555036
rect 473228 555024 473234 555076
rect 178034 554956 178040 555008
rect 178092 554996 178098 555008
rect 475194 554996 475200 555008
rect 178092 554968 475200 554996
rect 178092 554956 178098 554968
rect 475194 554956 475200 554968
rect 475252 554956 475258 555008
rect 220170 554888 220176 554940
rect 220228 554928 220234 554940
rect 523034 554928 523040 554940
rect 220228 554900 523040 554928
rect 220228 554888 220234 554900
rect 523034 554888 523040 554900
rect 523092 554888 523098 554940
rect 185762 554820 185768 554872
rect 185820 554860 185826 554872
rect 543734 554860 543740 554872
rect 185820 554832 543740 554860
rect 185820 554820 185826 554832
rect 543734 554820 543740 554832
rect 543792 554820 543798 554872
rect 78582 554752 78588 554804
rect 78640 554792 78646 554804
rect 86862 554792 86868 554804
rect 78640 554764 86868 554792
rect 78640 554752 78646 554764
rect 86862 554752 86868 554764
rect 86920 554752 86926 554804
rect 151354 554752 151360 554804
rect 151412 554792 151418 554804
rect 510154 554792 510160 554804
rect 151412 554764 510160 554792
rect 151412 554752 151418 554764
rect 510154 554752 510160 554764
rect 510212 554752 510218 554804
rect 57330 554684 57336 554736
rect 57388 554724 57394 554736
rect 375834 554724 375840 554736
rect 57388 554696 375840 554724
rect 57388 554684 57394 554696
rect 375834 554684 375840 554696
rect 375892 554684 375898 554736
rect 59998 554616 60004 554668
rect 60056 554656 60062 554668
rect 323762 554656 323768 554668
rect 60056 554628 323768 554656
rect 60056 554616 60062 554628
rect 323762 554616 323768 554628
rect 323820 554616 323826 554668
rect 173802 554548 173808 554600
rect 173860 554588 173866 554600
rect 378686 554588 378692 554600
rect 173860 554560 378692 554588
rect 173860 554548 173866 554560
rect 378686 554548 378692 554560
rect 378744 554548 378750 554600
rect 178034 554480 178040 554532
rect 178092 554520 178098 554532
rect 376846 554520 376852 554532
rect 178092 554492 376852 554520
rect 178092 554480 178098 554492
rect 376846 554480 376852 554492
rect 376904 554480 376910 554532
rect 230382 554412 230388 554464
rect 230440 554452 230446 554464
rect 376754 554452 376760 554464
rect 230440 554424 376760 554452
rect 230440 554412 230446 554424
rect 376754 554412 376760 554424
rect 376812 554412 376818 554464
rect 240042 554344 240048 554396
rect 240100 554384 240106 554396
rect 376018 554384 376024 554396
rect 240100 554356 376024 554384
rect 240100 554344 240106 554356
rect 376018 554344 376024 554356
rect 376076 554344 376082 554396
rect 192938 554276 192944 554328
rect 192996 554316 193002 554328
rect 253566 554316 253572 554328
rect 192996 554288 253572 554316
rect 192996 554276 193002 554288
rect 253566 554276 253572 554288
rect 253624 554276 253630 554328
rect 256694 554276 256700 554328
rect 256752 554316 256758 554328
rect 376110 554316 376116 554328
rect 256752 554288 376116 554316
rect 256752 554276 256758 554288
rect 376110 554276 376116 554288
rect 376168 554276 376174 554328
rect 179046 554140 179052 554192
rect 179104 554180 179110 554192
rect 477218 554180 477224 554192
rect 179104 554152 477224 554180
rect 179104 554140 179110 554152
rect 477218 554140 477224 554152
rect 477276 554140 477282 554192
rect 174630 554072 174636 554124
rect 174688 554112 174694 554124
rect 482278 554112 482284 554124
rect 174688 554084 482284 554112
rect 174688 554072 174694 554084
rect 482278 554072 482284 554084
rect 482336 554072 482342 554124
rect 57606 554004 57612 554056
rect 57664 554044 57670 554056
rect 375742 554044 375748 554056
rect 57664 554016 375748 554044
rect 57664 554004 57670 554016
rect 375742 554004 375748 554016
rect 375800 554004 375806 554056
rect 496078 553528 496084 553580
rect 496136 553568 496142 553580
rect 497458 553568 497464 553580
rect 496136 553540 497464 553568
rect 496136 553528 496142 553540
rect 497458 553528 497464 553540
rect 497516 553528 497522 553580
rect 219158 553460 219164 553512
rect 219216 553500 219222 553512
rect 523126 553500 523132 553512
rect 219216 553472 523132 553500
rect 219216 553460 219222 553472
rect 523126 553460 523132 553472
rect 523184 553460 523190 553512
rect 177942 553392 177948 553444
rect 178000 553432 178006 553444
rect 513558 553432 513564 553444
rect 178000 553404 513564 553432
rect 178000 553392 178006 553404
rect 513558 553392 513564 553404
rect 513616 553392 513622 553444
rect 59170 553324 59176 553376
rect 59228 553364 59234 553376
rect 379790 553364 379796 553376
rect 59228 553336 379796 553364
rect 59228 553324 59234 553336
rect 379790 553324 379796 553336
rect 379848 553324 379854 553376
rect 56502 553256 56508 553308
rect 56560 553296 56566 553308
rect 369302 553296 369308 553308
rect 56560 553268 369308 553296
rect 56560 553256 56566 553268
rect 369302 553256 369308 553268
rect 369360 553256 369366 553308
rect 98638 553188 98644 553240
rect 98696 553228 98702 553240
rect 378134 553228 378140 553240
rect 98696 553200 378140 553228
rect 98696 553188 98702 553200
rect 378134 553188 378140 553200
rect 378192 553188 378198 553240
rect 97902 553120 97908 553172
rect 97960 553160 97966 553172
rect 326798 553160 326804 553172
rect 97960 553132 326804 553160
rect 97960 553120 97966 553132
rect 326798 553120 326804 553132
rect 326856 553120 326862 553172
rect 60826 553052 60832 553104
rect 60884 553092 60890 553104
rect 156690 553092 156696 553104
rect 60884 553064 156696 553092
rect 60884 553052 60890 553064
rect 156690 553052 156696 553064
rect 156748 553052 156754 553104
rect 191742 553052 191748 553104
rect 191800 553092 191806 553104
rect 253014 553092 253020 553104
rect 191800 553064 253020 553092
rect 191800 553052 191806 553064
rect 253014 553052 253020 553064
rect 253072 553052 253078 553104
rect 170766 552780 170772 552832
rect 170824 552820 170830 552832
rect 463050 552820 463056 552832
rect 170824 552792 463056 552820
rect 170824 552780 170830 552792
rect 463050 552780 463056 552792
rect 463108 552780 463114 552832
rect 208118 552712 208124 552764
rect 208176 552752 208182 552764
rect 530026 552752 530032 552764
rect 208176 552724 530032 552752
rect 208176 552712 208182 552724
rect 530026 552712 530032 552724
rect 530084 552712 530090 552764
rect 184842 552644 184848 552696
rect 184900 552684 184906 552696
rect 519354 552684 519360 552696
rect 184900 552656 519360 552684
rect 184900 552644 184906 552656
rect 519354 552644 519360 552656
rect 519412 552644 519418 552696
rect 253198 552236 253204 552288
rect 253256 552276 253262 552288
rect 343634 552276 343640 552288
rect 253256 552248 343640 552276
rect 253256 552236 253262 552248
rect 343634 552236 343640 552248
rect 343692 552236 343698 552288
rect 88978 552168 88984 552220
rect 89036 552208 89042 552220
rect 91094 552208 91100 552220
rect 89036 552180 91100 552208
rect 89036 552168 89042 552180
rect 91094 552168 91100 552180
rect 91152 552168 91158 552220
rect 249702 552168 249708 552220
rect 249760 552208 249766 552220
rect 344646 552208 344652 552220
rect 249760 552180 344652 552208
rect 249760 552168 249766 552180
rect 344646 552168 344652 552180
rect 344704 552168 344710 552220
rect 114462 552100 114468 552152
rect 114520 552140 114526 552152
rect 351730 552140 351736 552152
rect 114520 552112 351736 552140
rect 114520 552100 114526 552112
rect 351730 552100 351736 552112
rect 351788 552100 351794 552152
rect 234614 552032 234620 552084
rect 234672 552072 234678 552084
rect 512914 552072 512920 552084
rect 234672 552044 512920 552072
rect 234672 552032 234678 552044
rect 512914 552032 512920 552044
rect 512972 552032 512978 552084
rect 81434 551964 81440 552016
rect 81492 552004 81498 552016
rect 346026 552004 346032 552016
rect 81492 551976 346032 552004
rect 81492 551964 81498 551976
rect 346026 551964 346032 551976
rect 346084 551964 346090 552016
rect 433978 551964 433984 552016
rect 434036 552004 434042 552016
rect 436094 552004 436100 552016
rect 434036 551976 436100 552004
rect 434036 551964 434042 551976
rect 436094 551964 436100 551976
rect 436152 551964 436158 552016
rect 490466 551964 490472 552016
rect 490524 552004 490530 552016
rect 493318 552004 493324 552016
rect 490524 551976 493324 552004
rect 490524 551964 490530 551976
rect 493318 551964 493324 551976
rect 493376 551964 493382 552016
rect 111794 551896 111800 551948
rect 111852 551936 111858 551948
rect 374638 551936 374644 551948
rect 111852 551908 374644 551936
rect 111852 551896 111858 551908
rect 374638 551896 374644 551908
rect 374696 551896 374702 551948
rect 172422 551828 172428 551880
rect 172480 551868 172486 551880
rect 381262 551868 381268 551880
rect 172480 551840 381268 551868
rect 172480 551828 172486 551840
rect 381262 551828 381268 551840
rect 381320 551828 381326 551880
rect 118694 551760 118700 551812
rect 118752 551800 118758 551812
rect 317690 551800 317696 551812
rect 118752 551772 317696 551800
rect 118752 551760 118758 551772
rect 317690 551760 317696 551772
rect 317748 551760 317754 551812
rect 175826 551692 175832 551744
rect 175884 551732 175890 551744
rect 297450 551732 297456 551744
rect 175884 551704 297456 551732
rect 175884 551692 175890 551704
rect 297450 551692 297456 551704
rect 297508 551692 297514 551744
rect 204070 551420 204076 551472
rect 204128 551460 204134 551472
rect 507394 551460 507400 551472
rect 204128 551432 507400 551460
rect 204128 551420 204134 551432
rect 507394 551420 507400 551432
rect 507452 551420 507458 551472
rect 174262 551352 174268 551404
rect 174320 551392 174326 551404
rect 486326 551392 486332 551404
rect 174320 551364 486332 551392
rect 174320 551352 174326 551364
rect 486326 551352 486332 551364
rect 486384 551352 486390 551404
rect 189902 551284 189908 551336
rect 189960 551324 189966 551336
rect 508038 551324 508044 551336
rect 189960 551296 508044 551324
rect 189960 551284 189966 551296
rect 508038 551284 508044 551296
rect 508096 551284 508102 551336
rect 235994 550808 236000 550860
rect 236052 550848 236058 550860
rect 360838 550848 360844 550860
rect 236052 550820 360844 550848
rect 236052 550808 236058 550820
rect 360838 550808 360844 550820
rect 360896 550808 360902 550860
rect 224218 550740 224224 550792
rect 224276 550780 224282 550792
rect 518894 550780 518900 550792
rect 224276 550752 518900 550780
rect 224276 550740 224282 550752
rect 518894 550740 518900 550752
rect 518952 550740 518958 550792
rect 180058 550672 180064 550724
rect 180116 550712 180122 550724
rect 526254 550712 526260 550724
rect 180116 550684 526260 550712
rect 180116 550672 180122 550684
rect 526254 550672 526260 550684
rect 526312 550672 526318 550724
rect 163498 550604 163504 550656
rect 163556 550644 163562 550656
rect 509234 550644 509240 550656
rect 163556 550616 509240 550644
rect 163556 550604 163562 550616
rect 509234 550604 509240 550616
rect 509292 550604 509298 550656
rect 75914 550536 75920 550588
rect 75972 550576 75978 550588
rect 78582 550576 78588 550588
rect 75972 550548 78588 550576
rect 75972 550536 75978 550548
rect 78582 550536 78588 550548
rect 78640 550536 78646 550588
rect 80054 550536 80060 550588
rect 80112 550576 80118 550588
rect 344002 550576 344008 550588
rect 80112 550548 344008 550576
rect 80112 550536 80118 550548
rect 344002 550536 344008 550548
rect 344060 550536 344066 550588
rect 99374 550468 99380 550520
rect 99432 550508 99438 550520
rect 327810 550508 327816 550520
rect 99432 550480 327816 550508
rect 99432 550468 99438 550480
rect 327810 550468 327816 550480
rect 327868 550468 327874 550520
rect 92474 550400 92480 550452
rect 92532 550440 92538 550452
rect 153930 550440 153936 550452
rect 92532 550412 153936 550440
rect 92532 550400 92538 550412
rect 153930 550400 153936 550412
rect 153988 550400 153994 550452
rect 173802 550400 173808 550452
rect 173860 550440 173866 550452
rect 379514 550440 379520 550452
rect 173860 550412 379520 550440
rect 173860 550400 173866 550412
rect 379514 550400 379520 550412
rect 379572 550400 379578 550452
rect 168374 550332 168380 550384
rect 168432 550372 168438 550384
rect 304534 550372 304540 550384
rect 168432 550344 304540 550372
rect 168432 550332 168438 550344
rect 304534 550332 304540 550344
rect 304592 550332 304598 550384
rect 137738 550128 137744 550180
rect 137796 550168 137802 550180
rect 418798 550168 418804 550180
rect 137796 550140 418804 550168
rect 137796 550128 137802 550140
rect 418798 550128 418804 550140
rect 418856 550128 418862 550180
rect 226058 550060 226064 550112
rect 226116 550100 226122 550112
rect 510798 550100 510804 550112
rect 226116 550072 510804 550100
rect 226116 550060 226122 550072
rect 510798 550060 510804 550072
rect 510856 550060 510862 550112
rect 210878 549992 210884 550044
rect 210936 550032 210942 550044
rect 506566 550032 506572 550044
rect 210936 550004 506572 550032
rect 210936 549992 210942 550004
rect 506566 549992 506572 550004
rect 506624 549992 506630 550044
rect 60090 549924 60096 549976
rect 60148 549964 60154 549976
rect 378594 549964 378600 549976
rect 60148 549936 378600 549964
rect 60148 549924 60154 549936
rect 378594 549924 378600 549936
rect 378652 549924 378658 549976
rect 79594 549856 79600 549908
rect 79652 549896 79658 549908
rect 88978 549896 88984 549908
rect 79652 549868 88984 549896
rect 79652 549856 79658 549868
rect 88978 549856 88984 549868
rect 89036 549856 89042 549908
rect 177390 549856 177396 549908
rect 177448 549896 177454 549908
rect 514938 549896 514944 549908
rect 177448 549868 514944 549896
rect 177448 549856 177454 549868
rect 514938 549856 514944 549868
rect 514996 549856 515002 549908
rect 131114 549380 131120 549432
rect 131172 549420 131178 549432
rect 372982 549420 372988 549432
rect 131172 549392 372988 549420
rect 131172 549380 131178 549392
rect 372982 549380 372988 549392
rect 373040 549380 373046 549432
rect 221182 549312 221188 549364
rect 221240 549352 221246 549364
rect 524414 549352 524420 549364
rect 221240 549324 524420 549352
rect 221240 549312 221246 549324
rect 524414 549312 524420 549324
rect 524472 549312 524478 549364
rect 176562 549244 176568 549296
rect 176620 549284 176626 549296
rect 537110 549284 537116 549296
rect 176620 549256 537116 549284
rect 176620 549244 176626 549256
rect 537110 549244 537116 549256
rect 537168 549244 537174 549296
rect 79318 549176 79324 549228
rect 79376 549216 79382 549228
rect 380158 549216 380164 549228
rect 79376 549188 380164 549216
rect 79376 549176 79382 549188
rect 380158 549176 380164 549188
rect 380216 549176 380222 549228
rect 110414 549108 110420 549160
rect 110472 549148 110478 549160
rect 354122 549148 354128 549160
rect 110472 549120 354128 549148
rect 110472 549108 110478 549120
rect 354122 549108 354128 549120
rect 354180 549108 354186 549160
rect 178034 549040 178040 549092
rect 178092 549080 178098 549092
rect 381354 549080 381360 549092
rect 178092 549052 381360 549080
rect 178092 549040 178098 549052
rect 381354 549040 381360 549052
rect 381412 549040 381418 549092
rect 169754 548972 169760 549024
rect 169812 549012 169818 549024
rect 348050 549012 348056 549024
rect 169812 548984 348056 549012
rect 169812 548972 169818 548984
rect 348050 548972 348056 548984
rect 348108 548972 348114 549024
rect 175182 548904 175188 548956
rect 175240 548944 175246 548956
rect 254486 548944 254492 548956
rect 175240 548916 254492 548944
rect 175240 548904 175246 548916
rect 254486 548904 254492 548916
rect 254544 548904 254550 548956
rect 459094 548768 459100 548820
rect 459152 548808 459158 548820
rect 466914 548808 466920 548820
rect 459152 548780 466920 548808
rect 459152 548768 459158 548780
rect 466914 548768 466920 548780
rect 466972 548768 466978 548820
rect 198734 548700 198740 548752
rect 198792 548740 198798 548752
rect 505370 548740 505376 548752
rect 198792 548712 505376 548740
rect 198792 548700 198798 548712
rect 505370 548700 505376 548712
rect 505428 548700 505434 548752
rect 211890 548632 211896 548684
rect 211948 548672 211954 548684
rect 526070 548672 526076 548684
rect 211948 548644 526076 548672
rect 211948 548632 211954 548644
rect 526070 548632 526076 548644
rect 526128 548632 526134 548684
rect 200758 548564 200764 548616
rect 200816 548604 200822 548616
rect 523494 548604 523500 548616
rect 200816 548576 523500 548604
rect 200816 548564 200822 548576
rect 523494 548564 523500 548576
rect 523552 548564 523558 548616
rect 166350 548496 166356 548548
rect 166408 548536 166414 548548
rect 492398 548536 492404 548548
rect 166408 548508 492404 548536
rect 166408 548496 166414 548508
rect 492398 548496 492404 548508
rect 492456 548496 492462 548548
rect 436094 548360 436100 548412
rect 436152 548400 436158 548412
rect 441614 548400 441620 548412
rect 436152 548372 441620 548400
rect 436152 548360 436158 548372
rect 441614 548360 441620 548372
rect 441672 548360 441678 548412
rect 227714 548088 227720 548140
rect 227772 548128 227778 548140
rect 462038 548128 462044 548140
rect 227772 548100 462044 548128
rect 227772 548088 227778 548100
rect 462038 548088 462044 548100
rect 462096 548088 462102 548140
rect 253198 548020 253204 548072
rect 253256 548060 253262 548072
rect 500310 548060 500316 548072
rect 253256 548032 500316 548060
rect 253256 548020 253262 548032
rect 500310 548020 500316 548032
rect 500368 548020 500374 548072
rect 161474 547952 161480 548004
rect 161532 547992 161538 548004
rect 506474 547992 506480 548004
rect 161532 547964 506480 547992
rect 161532 547952 161538 547964
rect 506474 547952 506480 547964
rect 506532 547952 506538 548004
rect 93670 547884 93676 547936
rect 93728 547924 93734 547936
rect 520642 547924 520648 547936
rect 93728 547896 520648 547924
rect 93728 547884 93734 547896
rect 520642 547884 520648 547896
rect 520700 547884 520706 547936
rect 67542 547816 67548 547868
rect 67600 547856 67606 547868
rect 347038 547856 347044 547868
rect 67600 547828 347044 547856
rect 67600 547816 67606 547828
rect 347038 547816 347044 547828
rect 347096 547816 347102 547868
rect 88978 547748 88984 547800
rect 89036 547788 89042 547800
rect 151078 547788 151084 547800
rect 89036 547760 151084 547788
rect 89036 547748 89042 547760
rect 151078 547748 151084 547760
rect 151136 547748 151142 547800
rect 166166 547748 166172 547800
rect 166224 547788 166230 547800
rect 383930 547788 383936 547800
rect 166224 547760 383936 547788
rect 166224 547748 166230 547760
rect 383930 547748 383936 547760
rect 383988 547748 383994 547800
rect 136542 547680 136548 547732
rect 136600 547720 136606 547732
rect 320726 547720 320732 547732
rect 136600 547692 320732 547720
rect 136600 547680 136606 547692
rect 320726 547680 320732 547692
rect 320784 547680 320790 547732
rect 172054 547272 172060 547324
rect 172112 547312 172118 547324
rect 467006 547312 467012 547324
rect 172112 547284 467012 547312
rect 172112 547272 172118 547284
rect 467006 547272 467012 547284
rect 467064 547272 467070 547324
rect 185578 547204 185584 547256
rect 185636 547244 185642 547256
rect 508130 547244 508136 547256
rect 185636 547216 508136 547244
rect 185636 547204 185642 547216
rect 508130 547204 508136 547216
rect 508188 547204 508194 547256
rect 182542 547136 182548 547188
rect 182600 547176 182606 547188
rect 527358 547176 527364 547188
rect 182600 547148 527364 547176
rect 182600 547136 182606 547148
rect 527358 547136 527364 547148
rect 527416 547136 527422 547188
rect 231762 546796 231768 546848
rect 231820 546836 231826 546848
rect 365898 546836 365904 546848
rect 231820 546808 365904 546836
rect 231820 546796 231826 546808
rect 365898 546796 365904 546808
rect 365956 546796 365962 546848
rect 246298 546728 246304 546780
rect 246356 546768 246362 546780
rect 496078 546768 496084 546780
rect 246356 546740 496084 546768
rect 246356 546728 246362 546740
rect 496078 546728 496084 546740
rect 496136 546728 496142 546780
rect 187786 546660 187792 546712
rect 187844 546700 187850 546712
rect 503714 546700 503720 546712
rect 187844 546672 503720 546700
rect 187844 546660 187850 546672
rect 503714 546660 503720 546672
rect 503772 546660 503778 546712
rect 175642 546592 175648 546644
rect 175700 546632 175706 546644
rect 531314 546632 531320 546644
rect 175700 546604 531320 546632
rect 175700 546592 175706 546604
rect 531314 546592 531320 546604
rect 531372 546592 531378 546644
rect 175182 546524 175188 546576
rect 175240 546564 175246 546576
rect 540330 546564 540336 546576
rect 175240 546536 540336 546564
rect 175240 546524 175246 546536
rect 540330 546524 540336 546536
rect 540388 546524 540394 546576
rect 77294 546456 77300 546508
rect 77352 546496 77358 546508
rect 79594 546496 79600 546508
rect 77352 546468 79600 546496
rect 77352 546456 77358 546468
rect 79594 546456 79600 546468
rect 79652 546456 79658 546508
rect 90634 546456 90640 546508
rect 90692 546496 90698 546508
rect 520550 546496 520556 546508
rect 90692 546468 520556 546496
rect 90692 546456 90698 546468
rect 520550 546456 520556 546468
rect 520608 546456 520614 546508
rect 56502 546388 56508 546440
rect 56560 546428 56566 546440
rect 359182 546428 359188 546440
rect 56560 546400 359188 546428
rect 56560 546388 56566 546400
rect 359182 546388 359188 546400
rect 359240 546388 359246 546440
rect 75822 546320 75828 546372
rect 75880 546360 75886 546372
rect 350074 546360 350080 546372
rect 75880 546332 350080 546360
rect 75880 546320 75886 546332
rect 350074 546320 350080 546332
rect 350132 546320 350138 546372
rect 86862 546252 86868 546304
rect 86920 546292 86926 546304
rect 335906 546292 335912 546304
rect 86920 546264 335912 546292
rect 86920 546252 86926 546264
rect 335906 546252 335912 546264
rect 335964 546252 335970 546304
rect 126882 546184 126888 546236
rect 126940 546224 126946 546236
rect 313642 546224 313648 546236
rect 126940 546196 313648 546224
rect 126940 546184 126946 546196
rect 313642 546184 313648 546196
rect 313700 546184 313706 546236
rect 224126 546116 224132 546168
rect 224184 546156 224190 546168
rect 307570 546156 307576 546168
rect 224184 546128 307576 546156
rect 224184 546116 224190 546128
rect 307570 546116 307576 546128
rect 307628 546116 307634 546168
rect 299658 546048 299664 546100
rect 299716 546088 299722 546100
rect 538398 546088 538404 546100
rect 299716 546060 538404 546088
rect 299716 546048 299722 546060
rect 538398 546048 538404 546060
rect 538456 546048 538462 546100
rect 289630 545980 289636 546032
rect 289688 546020 289694 546032
rect 541526 546020 541532 546032
rect 289688 545992 541532 546020
rect 289688 545980 289694 545992
rect 541526 545980 541532 545992
rect 541584 545980 541590 546032
rect 173434 545912 173440 545964
rect 173492 545952 173498 545964
rect 483290 545952 483296 545964
rect 173492 545924 483296 545952
rect 173492 545912 173498 545924
rect 483290 545912 483296 545924
rect 483348 545912 483354 545964
rect 196710 545844 196716 545896
rect 196768 545884 196774 545896
rect 528922 545884 528928 545896
rect 196768 545856 528928 545884
rect 196768 545844 196774 545856
rect 528922 545844 528928 545856
rect 528980 545844 528986 545896
rect 183554 545776 183560 545828
rect 183612 545816 183618 545828
rect 528830 545816 528836 545828
rect 183612 545788 528836 545816
rect 183612 545776 183618 545788
rect 528830 545776 528836 545788
rect 528888 545776 528894 545828
rect 179598 545708 179604 545760
rect 179656 545748 179662 545760
rect 538490 545748 538496 545760
rect 179656 545720 538496 545748
rect 179656 545708 179662 545720
rect 538490 545708 538496 545720
rect 538548 545708 538554 545760
rect 192846 545164 192852 545216
rect 192904 545204 192910 545216
rect 253934 545204 253940 545216
rect 192904 545176 253940 545204
rect 192904 545164 192910 545176
rect 253934 545164 253940 545176
rect 253992 545164 253998 545216
rect 441614 545164 441620 545216
rect 441672 545204 441678 545216
rect 444374 545204 444380 545216
rect 441672 545176 444380 545204
rect 441672 545164 441678 545176
rect 444374 545164 444380 545176
rect 444432 545164 444438 545216
rect 493318 545164 493324 545216
rect 493376 545204 493382 545216
rect 496170 545204 496176 545216
rect 493376 545176 496176 545204
rect 493376 545164 493382 545176
rect 496170 545164 496176 545176
rect 496228 545164 496234 545216
rect 218146 545096 218152 545148
rect 218204 545136 218210 545148
rect 522574 545136 522580 545148
rect 218204 545108 522580 545136
rect 218204 545096 218210 545108
rect 522574 545096 522580 545108
rect 522632 545096 522638 545148
rect 75822 545028 75828 545080
rect 75880 545068 75886 545080
rect 364242 545068 364248 545080
rect 75880 545040 364248 545068
rect 75880 545028 75886 545040
rect 364242 545028 364248 545040
rect 364300 545028 364306 545080
rect 88242 544960 88248 545012
rect 88300 545000 88306 545012
rect 329834 545000 329840 545012
rect 88300 544972 329840 545000
rect 88300 544960 88306 544972
rect 329834 544960 329840 544972
rect 329892 544960 329898 545012
rect 131114 544892 131120 544944
rect 131172 544932 131178 544944
rect 324774 544932 324780 544944
rect 131172 544904 324780 544932
rect 131172 544892 131178 544904
rect 324774 544892 324780 544904
rect 324832 544892 324838 544944
rect 169754 544824 169760 544876
rect 169812 544864 169818 544876
rect 253474 544864 253480 544876
rect 169812 544836 253480 544864
rect 169812 544824 169818 544836
rect 253474 544824 253480 544836
rect 253532 544824 253538 544876
rect 216674 544756 216680 544808
rect 216732 544796 216738 544808
rect 250438 544796 250444 544808
rect 216732 544768 250444 544796
rect 216732 544756 216738 544768
rect 250438 544756 250444 544768
rect 250496 544756 250502 544808
rect 251818 544620 251824 544672
rect 251876 544660 251882 544672
rect 545666 544660 545672 544672
rect 251876 544632 545672 544660
rect 251876 544620 251882 544632
rect 545666 544620 545672 544632
rect 545724 544620 545730 544672
rect 170582 544552 170588 544604
rect 170640 544592 170646 544604
rect 465074 544592 465080 544604
rect 170640 544564 465080 544592
rect 170640 544552 170646 544564
rect 465074 544552 465080 544564
rect 465132 544552 465138 544604
rect 202782 544484 202788 544536
rect 202840 544524 202846 544536
rect 506658 544524 506664 544536
rect 202840 544496 506664 544524
rect 202840 544484 202846 544496
rect 506658 544484 506664 544496
rect 506716 544484 506722 544536
rect 209866 544416 209872 544468
rect 209924 544456 209930 544468
rect 530210 544456 530216 544468
rect 209924 544428 530216 544456
rect 209924 544416 209930 544428
rect 530210 544416 530216 544428
rect 530268 544416 530274 544468
rect 177482 544348 177488 544400
rect 177540 544388 177546 544400
rect 515122 544388 515128 544400
rect 177540 544360 515128 544388
rect 177540 544348 177546 544360
rect 515122 544348 515128 544360
rect 515180 544348 515186 544400
rect 252462 543872 252468 543924
rect 252520 543912 252526 543924
rect 526162 543912 526168 543924
rect 252520 543884 526168 543912
rect 252520 543872 252526 543884
rect 526162 543872 526168 543884
rect 526220 543872 526226 543924
rect 181714 543804 181720 543856
rect 181772 543844 181778 543856
rect 539870 543844 539876 543856
rect 181772 543816 539876 543844
rect 181772 543804 181778 543816
rect 539870 543804 539876 543816
rect 539928 543804 539934 543856
rect 75730 543776 75736 543788
rect 74506 543748 75736 543776
rect 72418 543668 72424 543720
rect 72476 543708 72482 543720
rect 74506 543708 74534 543748
rect 75730 543736 75736 543748
rect 75788 543736 75794 543788
rect 94682 543736 94688 543788
rect 94740 543776 94746 543788
rect 523402 543776 523408 543788
rect 94740 543748 523408 543776
rect 94740 543736 94746 543748
rect 523402 543736 523408 543748
rect 523460 543736 523466 543788
rect 72476 543680 74534 543708
rect 72476 543668 72482 543680
rect 128722 543668 128728 543720
rect 128780 543708 128786 543720
rect 134518 543708 134524 543720
rect 128780 543680 134524 543708
rect 128780 543668 128786 543680
rect 134518 543668 134524 543680
rect 134576 543668 134582 543720
rect 362218 543708 362224 543720
rect 142126 543680 362224 543708
rect 127618 543600 127624 543652
rect 127676 543640 127682 543652
rect 142126 543640 142154 543680
rect 362218 543668 362224 543680
rect 362276 543668 362282 543720
rect 127676 543612 142154 543640
rect 127676 543600 127682 543612
rect 208394 543600 208400 543652
rect 208452 543640 208458 543652
rect 360194 543640 360200 543652
rect 208452 543612 360200 543640
rect 208452 543600 208458 543612
rect 360194 543600 360200 543612
rect 360252 543600 360258 543652
rect 240042 543532 240048 543584
rect 240100 543572 240106 543584
rect 325786 543572 325792 543584
rect 240100 543544 325792 543572
rect 240100 543532 240106 543544
rect 325786 543532 325792 543544
rect 325844 543532 325850 543584
rect 244274 543464 244280 543516
rect 244332 543504 244338 543516
rect 259178 543504 259184 543516
rect 244332 543476 259184 543504
rect 244332 543464 244338 543476
rect 259178 543464 259184 543476
rect 259236 543464 259242 543516
rect 160738 543260 160744 543312
rect 160796 543300 160802 543312
rect 255038 543300 255044 543312
rect 160796 543272 255044 543300
rect 160796 543260 160802 543272
rect 255038 543260 255044 543272
rect 255096 543260 255102 543312
rect 191098 543192 191104 543244
rect 191156 543232 191162 543244
rect 382826 543232 382832 543244
rect 191156 543204 382832 543232
rect 191156 543192 191162 543204
rect 382826 543192 382832 543204
rect 382884 543192 382890 543244
rect 194686 543124 194692 543176
rect 194744 543164 194750 543176
rect 503806 543164 503812 543176
rect 194744 543136 503812 543164
rect 194744 543124 194750 543136
rect 503806 543124 503812 543136
rect 503864 543124 503870 543176
rect 173250 543056 173256 543108
rect 173308 543096 173314 543108
rect 485314 543096 485320 543108
rect 173308 543068 485320 543096
rect 173308 543056 173314 543068
rect 485314 543056 485320 543068
rect 485372 543056 485378 543108
rect 193674 542988 193680 543040
rect 193732 543028 193738 543040
rect 532970 543028 532976 543040
rect 193732 543000 532976 543028
rect 193732 542988 193738 543000
rect 532970 542988 532976 543000
rect 533028 542988 533034 543040
rect 466914 542920 466920 542972
rect 466972 542960 466978 542972
rect 470134 542960 470140 542972
rect 466972 542932 470140 542960
rect 466972 542920 466978 542932
rect 470134 542920 470140 542932
rect 470192 542920 470198 542972
rect 299198 542580 299204 542632
rect 299256 542620 299262 542632
rect 511166 542620 511172 542632
rect 299256 542592 511172 542620
rect 299256 542580 299262 542592
rect 511166 542580 511172 542592
rect 511224 542580 511230 542632
rect 242802 542512 242808 542564
rect 242860 542552 242866 542564
rect 503898 542552 503904 542564
rect 242860 542524 503904 542552
rect 242860 542512 242866 542524
rect 503898 542512 503904 542524
rect 503956 542512 503962 542564
rect 172606 542444 172612 542496
rect 172664 542484 172670 542496
rect 517698 542484 517704 542496
rect 172664 542456 517704 542484
rect 172664 542444 172670 542456
rect 517698 542444 517704 542456
rect 517756 542444 517762 542496
rect 91646 542376 91652 542428
rect 91704 542416 91710 542428
rect 517790 542416 517796 542428
rect 91704 542388 517796 542416
rect 91704 542376 91710 542388
rect 517790 542376 517796 542388
rect 517848 542376 517854 542428
rect 82814 542308 82820 542360
rect 82872 542348 82878 542360
rect 363230 542348 363236 542360
rect 82872 542320 363236 542348
rect 82872 542308 82878 542320
rect 363230 542308 363236 542320
rect 363288 542308 363294 542360
rect 178034 542240 178040 542292
rect 178092 542280 178098 542292
rect 383838 542280 383844 542292
rect 178092 542252 383844 542280
rect 178092 542240 178098 542252
rect 383838 542240 383844 542252
rect 383896 542240 383902 542292
rect 128354 542172 128360 542224
rect 128412 542212 128418 542224
rect 328822 542212 328828 542224
rect 128412 542184 328828 542212
rect 128412 542172 128418 542184
rect 328822 542172 328828 542184
rect 328880 542172 328886 542224
rect 129734 542104 129740 542156
rect 129792 542144 129798 542156
rect 316678 542144 316684 542156
rect 129792 542116 316684 542144
rect 129792 542104 129798 542116
rect 316678 542104 316684 542116
rect 316736 542104 316742 542156
rect 291838 541832 291844 541884
rect 291896 541872 291902 541884
rect 536282 541872 536288 541884
rect 291896 541844 536288 541872
rect 291896 541832 291902 541844
rect 536282 541832 536288 541844
rect 536340 541832 536346 541884
rect 171962 541764 171968 541816
rect 172020 541804 172026 541816
rect 468110 541804 468116 541816
rect 172020 541776 468116 541804
rect 172020 541764 172026 541776
rect 468110 541764 468116 541776
rect 468168 541764 468174 541816
rect 179690 541696 179696 541748
rect 179748 541736 179754 541748
rect 517974 541736 517980 541748
rect 179748 541708 517980 541736
rect 179748 541696 179754 541708
rect 517974 541696 517980 541708
rect 518032 541696 518038 541748
rect 181530 541628 181536 541680
rect 181588 541668 181594 541680
rect 527450 541668 527456 541680
rect 181588 541640 527456 541668
rect 181588 541628 181594 541640
rect 527450 541628 527456 541640
rect 527508 541628 527514 541680
rect 235994 541220 236000 541272
rect 236052 541260 236058 541272
rect 506750 541260 506756 541272
rect 236052 541232 506756 541260
rect 236052 541220 236058 541232
rect 506750 541220 506756 541232
rect 506808 541220 506814 541272
rect 172422 541152 172428 541204
rect 172480 541192 172486 541204
rect 516594 541192 516600 541204
rect 172480 541164 516600 541192
rect 172480 541152 172486 541164
rect 516594 541152 516600 541164
rect 516652 541152 516658 541204
rect 178678 541084 178684 541136
rect 178736 541124 178742 541136
rect 524506 541124 524512 541136
rect 178736 541096 524512 541124
rect 178736 541084 178742 541096
rect 524506 541084 524512 541096
rect 524564 541084 524570 541136
rect 148318 541016 148324 541068
rect 148376 541056 148382 541068
rect 506474 541056 506480 541068
rect 148376 541028 506480 541056
rect 148376 541016 148382 541028
rect 506474 541016 506480 541028
rect 506532 541016 506538 541068
rect 92658 540948 92664 541000
rect 92716 540988 92722 541000
rect 516502 540988 516508 541000
rect 92716 540960 516508 540988
rect 92716 540948 92722 540960
rect 516502 540948 516508 540960
rect 516560 540948 516566 541000
rect 91094 540880 91100 540932
rect 91152 540920 91158 540932
rect 368290 540920 368296 540932
rect 91152 540892 368296 540920
rect 91152 540880 91158 540892
rect 368290 540880 368296 540892
rect 368348 540880 368354 540932
rect 444374 540880 444380 540932
rect 444432 540920 444438 540932
rect 447226 540920 447232 540932
rect 444432 540892 447232 540920
rect 444432 540880 444438 540892
rect 447226 540880 447232 540892
rect 447284 540880 447290 540932
rect 107562 540812 107568 540864
rect 107620 540852 107626 540864
rect 345014 540852 345020 540864
rect 107620 540824 345020 540852
rect 107620 540812 107626 540824
rect 345014 540812 345020 540824
rect 345072 540812 345078 540864
rect 218054 540744 218060 540796
rect 218112 540784 218118 540796
rect 374730 540784 374736 540796
rect 218112 540756 374736 540784
rect 218112 540744 218118 540756
rect 374730 540744 374736 540756
rect 374788 540744 374794 540796
rect 169754 540676 169760 540728
rect 169812 540716 169818 540728
rect 254854 540716 254860 540728
rect 169812 540688 254860 540716
rect 169812 540676 169818 540688
rect 254854 540676 254860 540688
rect 254912 540676 254918 540728
rect 187602 540336 187608 540388
rect 187660 540376 187666 540388
rect 508222 540376 508228 540388
rect 187660 540348 508228 540376
rect 187660 540336 187666 540348
rect 508222 540336 508228 540348
rect 508280 540336 508286 540388
rect 177666 540268 177672 540320
rect 177724 540308 177730 540320
rect 515306 540308 515312 540320
rect 177724 540280 515312 540308
rect 177724 540268 177730 540280
rect 515306 540268 515312 540280
rect 515364 540268 515370 540320
rect 73154 540200 73160 540252
rect 73212 540240 73218 540252
rect 77294 540240 77300 540252
rect 73212 540212 77300 540240
rect 73212 540200 73218 540212
rect 77294 540200 77300 540212
rect 77352 540200 77358 540252
rect 92014 540200 92020 540252
rect 92072 540240 92078 540252
rect 144178 540240 144184 540252
rect 92072 540212 144184 540240
rect 92072 540200 92078 540212
rect 144178 540200 144184 540212
rect 144236 540200 144242 540252
rect 190638 540200 190644 540252
rect 190696 540240 190702 540252
rect 530118 540240 530124 540252
rect 190696 540212 530124 540240
rect 190696 540200 190702 540212
rect 530118 540200 530124 540212
rect 530176 540200 530182 540252
rect 244274 539928 244280 539980
rect 244332 539968 244338 539980
rect 254762 539968 254768 539980
rect 244332 539940 254768 539968
rect 244332 539928 244338 539940
rect 254762 539928 254768 539940
rect 254820 539928 254826 539980
rect 247034 539860 247040 539912
rect 247092 539900 247098 539912
rect 354766 539900 354772 539912
rect 247092 539872 354772 539900
rect 247092 539860 247098 539872
rect 354766 539860 354772 539872
rect 354824 539860 354830 539912
rect 175182 539792 175188 539844
rect 175240 539832 175246 539844
rect 466086 539832 466092 539844
rect 175240 539804 466092 539832
rect 175240 539792 175246 539804
rect 466086 539792 466092 539804
rect 466144 539792 466150 539844
rect 217134 539724 217140 539776
rect 217192 539764 217198 539776
rect 521654 539764 521660 539776
rect 217192 539736 521660 539764
rect 217192 539724 217198 539736
rect 521654 539724 521660 539736
rect 521712 539724 521718 539776
rect 158438 539656 158444 539708
rect 158496 539696 158502 539708
rect 500402 539696 500408 539708
rect 158496 539668 500408 539696
rect 158496 539656 158502 539668
rect 500402 539656 500408 539668
rect 500460 539656 500466 539708
rect 88610 539588 88616 539640
rect 88668 539628 88674 539640
rect 521654 539628 521660 539640
rect 88668 539600 521660 539628
rect 88668 539588 88674 539600
rect 521654 539588 521660 539600
rect 521712 539588 521718 539640
rect 60826 539520 60832 539572
rect 60884 539560 60890 539572
rect 371326 539560 371332 539572
rect 60884 539532 371332 539560
rect 60884 539520 60890 539532
rect 371326 539520 371332 539532
rect 371384 539520 371390 539572
rect 86862 539452 86868 539504
rect 86920 539492 86926 539504
rect 352098 539492 352104 539504
rect 86920 539464 352104 539492
rect 86920 539452 86926 539464
rect 352098 539452 352104 539464
rect 352156 539452 352162 539504
rect 100754 539384 100760 539436
rect 100812 539424 100818 539436
rect 340966 539424 340972 539436
rect 100812 539396 340972 539424
rect 100812 539384 100818 539396
rect 340966 539384 340972 539396
rect 341024 539384 341030 539436
rect 124858 539316 124864 539368
rect 124916 539356 124922 539368
rect 128722 539356 128728 539368
rect 124916 539328 128728 539356
rect 124916 539316 124922 539328
rect 128722 539316 128728 539328
rect 128780 539316 128786 539368
rect 136542 539316 136548 539368
rect 136600 539356 136606 539368
rect 331858 539356 331864 539368
rect 136600 539328 331864 539356
rect 136600 539316 136606 539328
rect 331858 539316 331864 539328
rect 331916 539316 331922 539368
rect 222102 539248 222108 539300
rect 222160 539288 222166 539300
rect 386598 539288 386604 539300
rect 222160 539260 386604 539288
rect 222160 539248 222166 539260
rect 386598 539248 386604 539260
rect 386656 539248 386662 539300
rect 206830 538908 206836 538960
rect 206888 538948 206894 538960
rect 506842 538948 506848 538960
rect 206888 538920 506848 538948
rect 206888 538908 206894 538920
rect 506842 538908 506848 538920
rect 506900 538908 506906 538960
rect 174538 538840 174544 538892
rect 174596 538880 174602 538892
rect 479242 538880 479248 538892
rect 174596 538852 479248 538880
rect 174596 538840 174602 538852
rect 479242 538840 479248 538852
rect 479300 538840 479306 538892
rect 104802 538500 104808 538552
rect 104860 538540 104866 538552
rect 375006 538540 375012 538552
rect 104860 538512 375012 538540
rect 104860 538500 104866 538512
rect 375006 538500 375012 538512
rect 375064 538500 375070 538552
rect 225506 538432 225512 538484
rect 225564 538472 225570 538484
rect 501046 538472 501052 538484
rect 225564 538444 501052 538472
rect 225564 538432 225570 538444
rect 501046 538432 501052 538444
rect 501104 538432 501110 538484
rect 156414 538364 156420 538416
rect 156472 538404 156478 538416
rect 496262 538404 496268 538416
rect 156472 538376 496268 538404
rect 156472 538364 156478 538376
rect 496262 538364 496268 538376
rect 496320 538364 496326 538416
rect 170582 538296 170588 538348
rect 170640 538336 170646 538348
rect 516134 538336 516140 538348
rect 170640 538308 516140 538336
rect 170640 538296 170646 538308
rect 516134 538296 516140 538308
rect 516192 538296 516198 538348
rect 179690 538228 179696 538280
rect 179748 538268 179754 538280
rect 536834 538268 536840 538280
rect 179748 538240 536840 538268
rect 179748 538228 179754 538240
rect 536834 538228 536840 538240
rect 536892 538228 536898 538280
rect 85482 538160 85488 538212
rect 85540 538200 85546 538212
rect 373350 538200 373356 538212
rect 85540 538172 373356 538200
rect 85540 538160 85546 538172
rect 373350 538160 373356 538172
rect 373408 538160 373414 538212
rect 117222 538092 117228 538144
rect 117280 538132 117286 538144
rect 330846 538132 330852 538144
rect 117280 538104 330852 538132
rect 117280 538092 117286 538104
rect 330846 538092 330852 538104
rect 330904 538092 330910 538144
rect 252462 538024 252468 538076
rect 252520 538064 252526 538076
rect 311618 538064 311624 538076
rect 252520 538036 311624 538064
rect 252520 538024 252526 538036
rect 311618 538024 311624 538036
rect 311676 538024 311682 538076
rect 205818 537616 205824 537668
rect 205876 537656 205882 537668
rect 505554 537656 505560 537668
rect 205876 537628 505560 537656
rect 205876 537616 205882 537628
rect 505554 537616 505560 537628
rect 505612 537616 505618 537668
rect 175918 537548 175924 537600
rect 175976 537588 175982 537600
rect 478322 537588 478328 537600
rect 175976 537560 478328 537588
rect 175976 537548 175982 537560
rect 478322 537548 478328 537560
rect 478380 537548 478386 537600
rect 172882 537480 172888 537532
rect 172940 537520 172946 537532
rect 488350 537520 488356 537532
rect 172940 537492 488356 537520
rect 172940 537480 172946 537492
rect 488350 537480 488356 537492
rect 488408 537480 488414 537532
rect 109034 537140 109040 537192
rect 109092 537180 109098 537192
rect 376018 537180 376024 537192
rect 109092 537152 376024 537180
rect 109092 537140 109098 537152
rect 376018 537140 376024 537152
rect 376076 537140 376082 537192
rect 213086 537072 213092 537124
rect 213144 537112 213150 537124
rect 518434 537112 518440 537124
rect 213144 537084 518440 537112
rect 213144 537072 213150 537084
rect 518434 537072 518440 537084
rect 518492 537072 518498 537124
rect 180702 537004 180708 537056
rect 180760 537044 180766 537056
rect 511534 537044 511540 537056
rect 180760 537016 511540 537044
rect 180760 537004 180766 537016
rect 511534 537004 511540 537016
rect 511592 537004 511598 537056
rect 190822 536936 190828 536988
rect 190880 536976 190886 536988
rect 543826 536976 543832 536988
rect 190880 536948 543832 536976
rect 190880 536936 190886 536948
rect 543826 536936 543832 536948
rect 543884 536936 543890 536988
rect 72418 536908 72424 536920
rect 69124 536880 72424 536908
rect 69124 536840 69152 536880
rect 72418 536868 72424 536880
rect 72476 536868 72482 536920
rect 166902 536868 166908 536920
rect 166960 536908 166966 536920
rect 527634 536908 527640 536920
rect 166960 536880 527640 536908
rect 166960 536868 166966 536880
rect 527634 536868 527640 536880
rect 527692 536868 527698 536920
rect 73154 536840 73160 536852
rect 68940 536812 69152 536840
rect 70412 536812 73160 536840
rect 66254 536732 66260 536784
rect 66312 536772 66318 536784
rect 68940 536772 68968 536812
rect 66312 536744 68968 536772
rect 66312 536732 66318 536744
rect 69014 536732 69020 536784
rect 69072 536772 69078 536784
rect 70412 536772 70440 536812
rect 73154 536800 73160 536812
rect 73212 536800 73218 536852
rect 84562 536800 84568 536852
rect 84620 536840 84626 536852
rect 520458 536840 520464 536852
rect 84620 536812 520464 536840
rect 84620 536800 84626 536812
rect 520458 536800 520464 536812
rect 520516 536800 520522 536852
rect 69072 536744 70440 536772
rect 69072 536732 69078 536744
rect 89714 536732 89720 536784
rect 89772 536772 89778 536784
rect 370314 536772 370320 536784
rect 89772 536744 370320 536772
rect 89772 536732 89778 536744
rect 370314 536732 370320 536744
rect 370372 536732 370378 536784
rect 109034 536664 109040 536716
rect 109092 536704 109098 536716
rect 342990 536704 342996 536716
rect 109092 536676 342996 536704
rect 109092 536664 109098 536676
rect 342990 536664 342996 536676
rect 343048 536664 343054 536716
rect 117222 536596 117228 536648
rect 117280 536636 117286 536648
rect 297358 536636 297364 536648
rect 117280 536608 297364 536636
rect 117280 536596 117286 536608
rect 297358 536596 297364 536608
rect 297416 536596 297422 536648
rect 168374 536528 168380 536580
rect 168432 536568 168438 536580
rect 301498 536568 301504 536580
rect 168432 536540 301504 536568
rect 168432 536528 168438 536540
rect 301498 536528 301504 536540
rect 301556 536528 301562 536580
rect 479702 536392 479708 536444
rect 479760 536432 479766 536444
rect 530394 536432 530400 536444
rect 479760 536404 530400 536432
rect 479760 536392 479766 536404
rect 530394 536392 530400 536404
rect 530452 536392 530458 536444
rect 447226 536324 447232 536376
rect 447284 536364 447290 536376
rect 456794 536364 456800 536376
rect 447284 536336 456800 536364
rect 447284 536324 447290 536336
rect 456794 536324 456800 536336
rect 456852 536324 456858 536376
rect 472986 536324 472992 536376
rect 473044 536364 473050 536376
rect 537294 536364 537300 536376
rect 473044 536336 537300 536364
rect 473044 536324 473050 536336
rect 537294 536324 537300 536336
rect 537352 536324 537358 536376
rect 456150 536256 456156 536308
rect 456208 536296 456214 536308
rect 535822 536296 535828 536308
rect 456208 536268 535828 536296
rect 456208 536256 456214 536268
rect 535822 536256 535828 536268
rect 535880 536256 535886 536308
rect 174722 536188 174728 536240
rect 174780 536228 174786 536240
rect 457990 536228 457996 536240
rect 174780 536200 457996 536228
rect 174780 536188 174786 536200
rect 457990 536188 457996 536200
rect 458048 536188 458054 536240
rect 459002 536188 459008 536240
rect 459060 536228 459066 536240
rect 524598 536228 524604 536240
rect 459060 536200 524604 536228
rect 459060 536188 459066 536200
rect 524598 536188 524604 536200
rect 524656 536188 524662 536240
rect 171778 536120 171784 536172
rect 171836 536160 171842 536172
rect 490374 536160 490380 536172
rect 171836 536132 490380 536160
rect 171836 536120 171842 536132
rect 490374 536120 490380 536132
rect 490432 536120 490438 536172
rect 186590 536052 186596 536104
rect 186648 536092 186654 536104
rect 508314 536092 508320 536104
rect 186648 536064 508320 536092
rect 186648 536052 186654 536064
rect 508314 536052 508320 536064
rect 508372 536052 508378 536104
rect 299382 535780 299388 535832
rect 299440 535820 299446 535832
rect 353754 535820 353760 535832
rect 299440 535792 353760 535820
rect 299440 535780 299446 535792
rect 353754 535780 353760 535792
rect 353812 535780 353818 535832
rect 175918 535712 175924 535764
rect 175976 535752 175982 535764
rect 355778 535752 355784 535764
rect 175976 535724 355784 535752
rect 175976 535712 175982 535724
rect 355778 535712 355784 535724
rect 355836 535712 355842 535764
rect 216122 535644 216128 535696
rect 216180 535684 216186 535696
rect 520274 535684 520280 535696
rect 216180 535656 520280 535684
rect 216180 535644 216186 535656
rect 520274 535644 520280 535656
rect 520332 535644 520338 535696
rect 241330 535576 241336 535628
rect 241388 535616 241394 535628
rect 545758 535616 545764 535628
rect 241388 535588 545764 535616
rect 241388 535576 241394 535588
rect 545758 535576 545764 535588
rect 545816 535576 545822 535628
rect 191834 535508 191840 535560
rect 191892 535548 191898 535560
rect 535362 535548 535368 535560
rect 191892 535520 535368 535548
rect 191892 535508 191898 535520
rect 535362 535508 535368 535520
rect 535420 535508 535426 535560
rect 85574 535440 85580 535492
rect 85632 535480 85638 535492
rect 519170 535480 519176 535492
rect 85632 535452 519176 535480
rect 85632 535440 85638 535452
rect 519170 535440 519176 535452
rect 519228 535440 519234 535492
rect 100754 535372 100760 535424
rect 100812 535412 100818 535424
rect 358170 535412 358176 535424
rect 100812 535384 358176 535412
rect 100812 535372 100818 535384
rect 358170 535372 358176 535384
rect 358228 535372 358234 535424
rect 169754 535304 169760 535356
rect 169812 535344 169818 535356
rect 334894 535344 334900 535356
rect 169812 535316 334900 535344
rect 169812 535304 169818 535316
rect 334894 535304 334900 535316
rect 334952 535304 334958 535356
rect 251082 535236 251088 535288
rect 251140 535276 251146 535288
rect 309594 535276 309600 535288
rect 251140 535248 309600 535276
rect 251140 535236 251146 535248
rect 309594 535236 309600 535248
rect 309652 535236 309658 535288
rect 60734 534896 60740 534948
rect 60792 534936 60798 534948
rect 348694 534936 348700 534948
rect 60792 534908 348700 534936
rect 60792 534896 60798 534908
rect 348694 534896 348700 534908
rect 348752 534896 348758 534948
rect 470134 534896 470140 534948
rect 470192 534936 470198 534948
rect 475838 534936 475844 534948
rect 470192 534908 475844 534936
rect 470192 534896 470198 534908
rect 475838 534896 475844 534908
rect 475896 534896 475902 534948
rect 212902 534828 212908 534880
rect 212960 534868 212966 534880
rect 506934 534868 506940 534880
rect 212960 534840 506940 534868
rect 212960 534828 212966 534840
rect 506934 534828 506940 534840
rect 506992 534828 506998 534880
rect 197722 534760 197728 534812
rect 197780 534800 197786 534812
rect 505738 534800 505744 534812
rect 197780 534772 505744 534800
rect 197780 534760 197786 534772
rect 505738 534760 505744 534772
rect 505796 534760 505802 534812
rect 63586 534692 63592 534744
rect 63644 534732 63650 534744
rect 69014 534732 69020 534744
rect 63644 534704 69020 534732
rect 63644 534692 63650 534704
rect 69014 534692 69020 534704
rect 69072 534692 69078 534744
rect 177758 534692 177764 534744
rect 177816 534732 177822 534744
rect 513834 534732 513840 534744
rect 177816 534704 513840 534732
rect 177816 534692 177822 534704
rect 513834 534692 513840 534704
rect 513892 534692 513898 534744
rect 108298 534352 108304 534404
rect 108356 534392 108362 534404
rect 377030 534392 377036 534404
rect 108356 534364 377036 534392
rect 108356 534352 108362 534364
rect 377030 534352 377036 534364
rect 377088 534352 377094 534404
rect 211062 534284 211068 534336
rect 211120 534324 211126 534336
rect 497550 534324 497556 534336
rect 211120 534296 497556 534324
rect 211120 534284 211126 534296
rect 497550 534284 497556 534296
rect 497608 534284 497614 534336
rect 209038 534216 209044 534268
rect 209096 534256 209102 534268
rect 527174 534256 527180 534268
rect 209096 534228 527180 534256
rect 209096 534216 209102 534228
rect 527174 534216 527180 534228
rect 527232 534216 527238 534268
rect 154390 534148 154396 534200
rect 154448 534188 154454 534200
rect 499574 534188 499580 534200
rect 154448 534160 499580 534188
rect 154448 534148 154454 534160
rect 499574 534148 499580 534160
rect 499632 534148 499638 534200
rect 157978 534080 157984 534132
rect 158036 534120 158042 534132
rect 160738 534120 160744 534132
rect 158036 534092 160744 534120
rect 158036 534080 158042 534092
rect 160738 534080 160744 534092
rect 160796 534080 160802 534132
rect 167546 534080 167552 534132
rect 167604 534120 167610 534132
rect 517054 534120 517060 534132
rect 167604 534092 517060 534120
rect 167604 534080 167610 534092
rect 517054 534080 517060 534092
rect 517112 534080 517118 534132
rect 106182 534012 106188 534064
rect 106240 534052 106246 534064
rect 366266 534052 366272 534064
rect 106240 534024 366272 534052
rect 106240 534012 106246 534024
rect 366266 534012 366272 534024
rect 366324 534012 366330 534064
rect 115842 533944 115848 533996
rect 115900 533984 115906 533996
rect 332870 533984 332876 533996
rect 115900 533956 332876 533984
rect 115900 533944 115906 533956
rect 332870 533944 332876 533956
rect 332928 533944 332934 533996
rect 175918 533876 175924 533928
rect 175976 533916 175982 533928
rect 339954 533916 339960 533928
rect 175976 533888 339960 533916
rect 175976 533876 175982 533888
rect 339954 533876 339960 533888
rect 340012 533876 340018 533928
rect 223482 533808 223488 533860
rect 223540 533848 223546 533860
rect 337930 533848 337936 533860
rect 223540 533820 337936 533848
rect 223540 533808 223546 533820
rect 337930 533808 337936 533820
rect 337988 533808 337994 533860
rect 195698 533536 195704 533588
rect 195756 533576 195762 533588
rect 505646 533576 505652 533588
rect 195756 533548 505652 533576
rect 195756 533536 195762 533548
rect 505646 533536 505652 533548
rect 505704 533536 505710 533588
rect 171870 533468 171876 533520
rect 171928 533508 171934 533520
rect 484302 533508 484308 533520
rect 171928 533480 484308 533508
rect 171928 533468 171934 533480
rect 484302 533468 484308 533480
rect 484360 533468 484366 533520
rect 489362 533468 489368 533520
rect 489420 533508 489426 533520
rect 544470 533508 544476 533520
rect 489420 533480 544476 533508
rect 489420 533468 489426 533480
rect 544470 533468 544476 533480
rect 544528 533468 544534 533520
rect 188614 533400 188620 533452
rect 188672 533440 188678 533452
rect 505462 533440 505468 533452
rect 188672 533412 505468 533440
rect 188672 533400 188678 533412
rect 505462 533400 505468 533412
rect 505520 533400 505526 533452
rect 177114 533332 177120 533384
rect 177172 533372 177178 533384
rect 513742 533372 513748 533384
rect 177172 533344 513748 533372
rect 177172 533332 177178 533344
rect 513742 533332 513748 533344
rect 513800 533332 513806 533384
rect 485038 533060 485044 533112
rect 485096 533100 485102 533112
rect 513926 533100 513932 533112
rect 485096 533072 513932 533100
rect 485096 533060 485102 533072
rect 513926 533060 513932 533072
rect 513984 533060 513990 533112
rect 251818 532992 251824 533044
rect 251876 533032 251882 533044
rect 509786 533032 509792 533044
rect 251876 533004 509792 533032
rect 251876 532992 251882 533004
rect 509786 532992 509792 533004
rect 509844 532992 509850 533044
rect 215110 532924 215116 532976
rect 215168 532964 215174 532976
rect 519078 532964 519084 532976
rect 215168 532936 519084 532964
rect 215168 532924 215174 532936
rect 519078 532924 519084 532936
rect 519136 532924 519142 532976
rect 194870 532856 194876 532908
rect 194928 532896 194934 532908
rect 538214 532896 538220 532908
rect 194928 532868 538220 532896
rect 194928 532856 194934 532868
rect 538214 532856 538220 532868
rect 538272 532856 538278 532908
rect 169570 532788 169576 532840
rect 169628 532828 169634 532840
rect 514754 532828 514760 532840
rect 169628 532800 514760 532828
rect 169628 532788 169634 532800
rect 514754 532788 514760 532800
rect 514812 532788 514818 532840
rect 83550 532720 83556 532772
rect 83608 532760 83614 532772
rect 518986 532760 518992 532772
rect 83608 532732 518992 532760
rect 83608 532720 83614 532732
rect 518986 532720 518992 532732
rect 519044 532720 519050 532772
rect 59630 532652 59636 532704
rect 59688 532692 59694 532704
rect 376294 532692 376300 532704
rect 59688 532664 376300 532692
rect 59688 532652 59694 532664
rect 376294 532652 376300 532664
rect 376352 532652 376358 532704
rect 215294 532584 215300 532636
rect 215352 532624 215358 532636
rect 374546 532624 374552 532636
rect 215352 532596 374552 532624
rect 215352 532584 215358 532596
rect 374546 532584 374552 532596
rect 374604 532584 374610 532636
rect 175458 532108 175464 532160
rect 175516 532148 175522 532160
rect 487338 532148 487344 532160
rect 175516 532120 487344 532148
rect 175516 532108 175522 532120
rect 487338 532108 487344 532120
rect 487396 532108 487402 532160
rect 57330 532040 57336 532092
rect 57388 532080 57394 532092
rect 376202 532080 376208 532092
rect 57388 532052 376208 532080
rect 57388 532040 57394 532052
rect 376202 532040 376208 532052
rect 376260 532040 376266 532092
rect 57422 531972 57428 532024
rect 57480 532012 57486 532024
rect 378318 532012 378324 532024
rect 57480 531984 378324 532012
rect 57480 531972 57486 531984
rect 378318 531972 378324 531984
rect 378376 531972 378382 532024
rect 254854 531700 254860 531752
rect 254912 531740 254918 531752
rect 521654 531740 521660 531752
rect 254912 531712 521660 531740
rect 254912 531700 254918 531712
rect 521654 531700 521660 531712
rect 521712 531700 521718 531752
rect 214098 531632 214104 531684
rect 214156 531672 214162 531684
rect 517606 531672 517612 531684
rect 214156 531644 517612 531672
rect 214156 531632 214162 531644
rect 517606 531632 517612 531644
rect 517664 531632 517670 531684
rect 198918 531564 198924 531616
rect 198976 531604 198982 531616
rect 507854 531604 507860 531616
rect 198976 531576 507860 531604
rect 198976 531564 198982 531576
rect 507854 531564 507860 531576
rect 507912 531564 507918 531616
rect 208026 531496 208032 531548
rect 208084 531536 208090 531548
rect 525794 531536 525800 531548
rect 208084 531508 525800 531536
rect 208084 531496 208090 531508
rect 525794 531496 525800 531508
rect 525852 531496 525858 531548
rect 168558 531428 168564 531480
rect 168616 531468 168622 531480
rect 499574 531468 499580 531480
rect 168616 531440 499580 531468
rect 168616 531428 168622 531440
rect 499574 531428 499580 531440
rect 499632 531428 499638 531480
rect 177942 531360 177948 531412
rect 178000 531400 178006 531412
rect 512822 531400 512828 531412
rect 178000 531372 512828 531400
rect 178000 531360 178006 531372
rect 512822 531360 512828 531372
rect 512880 531360 512886 531412
rect 529842 531400 529848 531412
rect 518866 531372 529848 531400
rect 66162 531332 66168 531344
rect 63512 531304 66168 531332
rect 62850 531224 62856 531276
rect 62908 531264 62914 531276
rect 63512 531264 63540 531304
rect 66162 531292 66168 531304
rect 66220 531292 66226 531344
rect 184750 531292 184756 531344
rect 184808 531332 184814 531344
rect 518866 531332 518894 531372
rect 529842 531360 529848 531372
rect 529900 531360 529906 531412
rect 184808 531304 518894 531332
rect 184808 531292 184814 531304
rect 62908 531236 63540 531264
rect 62908 531224 62914 531236
rect 166166 531224 166172 531276
rect 166224 531264 166230 531276
rect 374822 531264 374828 531276
rect 166224 531236 374828 531264
rect 166224 531224 166230 531236
rect 374822 531224 374828 531236
rect 374880 531224 374886 531276
rect 178218 531156 178224 531208
rect 178276 531196 178282 531208
rect 287790 531196 287796 531208
rect 178276 531168 287796 531196
rect 178276 531156 178282 531168
rect 287790 531156 287796 531168
rect 287848 531156 287854 531208
rect 178126 531088 178132 531140
rect 178184 531128 178190 531140
rect 280798 531128 280804 531140
rect 178184 531100 280804 531128
rect 178184 531088 178190 531100
rect 280798 531088 280804 531100
rect 280856 531088 280862 531140
rect 489454 531088 489460 531140
rect 489512 531128 489518 531140
rect 538582 531128 538588 531140
rect 489512 531100 538588 531128
rect 489512 531088 489518 531100
rect 538582 531088 538588 531100
rect 538640 531088 538646 531140
rect 476758 531020 476764 531072
rect 476816 531060 476822 531072
rect 534902 531060 534908 531072
rect 476816 531032 534908 531060
rect 476816 531020 476822 531032
rect 534902 531020 534908 531032
rect 534960 531020 534966 531072
rect 178862 530952 178868 531004
rect 178920 530952 178926 531004
rect 472894 530952 472900 531004
rect 472952 530992 472958 531004
rect 533246 530992 533252 531004
rect 472952 530964 533252 530992
rect 472952 530952 472958 530964
rect 533246 530952 533252 530964
rect 533304 530952 533310 531004
rect 178880 530800 178908 530952
rect 471514 530884 471520 530936
rect 471572 530924 471578 530936
rect 533338 530924 533344 530936
rect 471572 530896 533344 530924
rect 471572 530884 471578 530896
rect 533338 530884 533344 530896
rect 533396 530884 533402 530936
rect 464522 530816 464528 530868
rect 464580 530856 464586 530868
rect 530670 530856 530676 530868
rect 464580 530828 530676 530856
rect 464580 530816 464586 530828
rect 530670 530816 530676 530828
rect 530728 530816 530734 530868
rect 178862 530748 178868 530800
rect 178920 530748 178926 530800
rect 464338 530748 464344 530800
rect 464396 530788 464402 530800
rect 531682 530788 531688 530800
rect 464396 530760 531688 530788
rect 464396 530748 464402 530760
rect 531682 530748 531688 530760
rect 531740 530748 531746 530800
rect 465810 530680 465816 530732
rect 465868 530720 465874 530732
rect 534718 530720 534724 530732
rect 465868 530692 534724 530720
rect 465868 530680 465874 530692
rect 534718 530680 534724 530692
rect 534776 530680 534782 530732
rect 464614 530612 464620 530664
rect 464672 530652 464678 530664
rect 534534 530652 534540 530664
rect 464672 530624 534540 530652
rect 464672 530612 464678 530624
rect 534534 530612 534540 530624
rect 534592 530612 534598 530664
rect 137278 530544 137284 530596
rect 137336 530584 137342 530596
rect 342898 530584 342904 530596
rect 137336 530556 342904 530584
rect 137336 530544 137342 530556
rect 342898 530544 342904 530556
rect 342956 530544 342962 530596
rect 464430 530544 464436 530596
rect 464488 530584 464494 530596
rect 534626 530584 534632 530596
rect 464488 530556 534632 530584
rect 464488 530544 464494 530556
rect 534626 530544 534632 530556
rect 534684 530544 534690 530596
rect 164142 530476 164148 530528
rect 164200 530516 164206 530528
rect 313182 530516 313188 530528
rect 164200 530488 313188 530516
rect 164200 530476 164206 530488
rect 313182 530476 313188 530488
rect 313240 530476 313246 530528
rect 175918 530408 175924 530460
rect 175976 530448 175982 530460
rect 374086 530448 374092 530460
rect 175976 530420 374092 530448
rect 175976 530408 175982 530420
rect 374086 530408 374092 530420
rect 374144 530408 374150 530460
rect 256694 530340 256700 530392
rect 256752 530380 256758 530392
rect 469122 530380 469128 530392
rect 256752 530352 469128 530380
rect 256752 530340 256758 530352
rect 469122 530340 469128 530352
rect 469180 530340 469186 530392
rect 60182 530272 60188 530324
rect 60240 530312 60246 530324
rect 60240 530284 60734 530312
rect 60240 530272 60246 530284
rect 60706 530108 60734 530284
rect 285766 530272 285772 530324
rect 285824 530312 285830 530324
rect 521746 530312 521752 530324
rect 285824 530284 521752 530312
rect 285824 530272 285830 530284
rect 521746 530272 521752 530284
rect 521804 530272 521810 530324
rect 178034 530204 178040 530256
rect 178092 530244 178098 530256
rect 470134 530244 470140 530256
rect 178092 530216 470140 530244
rect 178092 530204 178098 530216
rect 470134 530204 470140 530216
rect 470192 530204 470198 530256
rect 62758 530136 62764 530188
rect 62816 530176 62822 530188
rect 138198 530176 138204 530188
rect 62816 530148 138204 530176
rect 62816 530136 62822 530148
rect 138198 530136 138204 530148
rect 138256 530136 138262 530188
rect 173802 530136 173808 530188
rect 173860 530176 173866 530188
rect 472158 530176 472164 530188
rect 173860 530148 472164 530176
rect 173860 530136 173866 530148
rect 472158 530136 472164 530148
rect 472216 530136 472222 530188
rect 140222 530108 140228 530120
rect 60706 530080 140228 530108
rect 140222 530068 140228 530080
rect 140280 530068 140286 530120
rect 212074 530068 212080 530120
rect 212132 530108 212138 530120
rect 516226 530108 516232 530120
rect 212132 530080 516232 530108
rect 212132 530068 212138 530080
rect 516226 530068 516232 530080
rect 516284 530068 516290 530120
rect 60274 530000 60280 530052
rect 60332 530040 60338 530052
rect 147306 530040 147312 530052
rect 60332 530012 147312 530040
rect 60332 530000 60338 530012
rect 147306 530000 147312 530012
rect 147364 530000 147370 530052
rect 195882 530000 195888 530052
rect 195940 530040 195946 530052
rect 541066 530040 541072 530052
rect 195940 530012 541072 530040
rect 195940 530000 195946 530012
rect 541066 530000 541072 530012
rect 541124 530000 541130 530052
rect 53742 529932 53748 529984
rect 53800 529972 53806 529984
rect 144270 529972 144276 529984
rect 53800 529944 144276 529972
rect 53800 529932 53806 529944
rect 144270 529932 144276 529944
rect 144328 529932 144334 529984
rect 183738 529932 183744 529984
rect 183796 529972 183802 529984
rect 540974 529972 540980 529984
rect 183796 529944 540980 529972
rect 183796 529932 183802 529944
rect 540974 529932 540980 529944
rect 541032 529932 541038 529984
rect 177850 529864 177856 529916
rect 177908 529904 177914 529916
rect 500954 529904 500960 529916
rect 177908 529876 500960 529904
rect 177908 529864 177914 529876
rect 500954 529864 500960 529876
rect 501012 529864 501018 529916
rect 96522 529796 96528 529848
rect 96580 529836 96586 529848
rect 382734 529836 382740 529848
rect 96580 529808 382740 529836
rect 96580 529796 96586 529808
rect 382734 529796 382740 529808
rect 382792 529796 382798 529848
rect 95142 529728 95148 529780
rect 95200 529768 95206 529780
rect 333882 529768 333888 529780
rect 95200 529740 333888 529768
rect 95200 529728 95206 529740
rect 333882 529728 333888 529740
rect 333940 529728 333946 529780
rect 95050 529660 95056 529712
rect 95108 529700 95114 529712
rect 321738 529700 321744 529712
rect 95108 529672 321744 529700
rect 95108 529660 95114 529672
rect 321738 529660 321744 529672
rect 321796 529660 321802 529712
rect 285674 529592 285680 529644
rect 285732 529632 285738 529644
rect 379882 529632 379888 529644
rect 285732 529604 379888 529632
rect 285732 529592 285738 529604
rect 379882 529592 379888 529604
rect 379940 529592 379946 529644
rect 456794 529524 456800 529576
rect 456852 529564 456858 529576
rect 501874 529564 501880 529576
rect 456852 529536 501880 529564
rect 456852 529524 456858 529536
rect 501874 529524 501880 529536
rect 501932 529524 501938 529576
rect 458818 529456 458824 529508
rect 458876 529496 458882 529508
rect 531590 529496 531596 529508
rect 458876 529468 531596 529496
rect 458876 529456 458882 529468
rect 531590 529456 531596 529468
rect 531648 529456 531654 529508
rect 213914 529388 213920 529440
rect 213972 529428 213978 529440
rect 511074 529428 511080 529440
rect 213972 529400 511080 529428
rect 213972 529388 213978 529400
rect 511074 529388 511080 529400
rect 511132 529388 511138 529440
rect 173158 529320 173164 529372
rect 173216 529360 173222 529372
rect 481266 529360 481272 529372
rect 173216 529332 481272 529360
rect 173216 529320 173222 529332
rect 481266 529320 481272 529332
rect 481324 529320 481330 529372
rect 486510 529320 486516 529372
rect 486568 529360 486574 529372
rect 527542 529360 527548 529372
rect 486568 529332 527548 529360
rect 486568 529320 486574 529332
rect 527542 529320 527548 529332
rect 527600 529320 527606 529372
rect 177022 529252 177028 529304
rect 177080 529292 177086 529304
rect 509786 529292 509792 529304
rect 177080 529264 509792 529292
rect 177080 529252 177086 529264
rect 509786 529252 509792 529264
rect 509844 529252 509850 529304
rect 61102 529184 61108 529236
rect 61160 529224 61166 529236
rect 61562 529224 61568 529236
rect 61160 529196 61568 529224
rect 61160 529184 61166 529196
rect 61562 529184 61568 529196
rect 61620 529184 61626 529236
rect 96890 529184 96896 529236
rect 96948 529224 96954 529236
rect 436002 529224 436008 529236
rect 96948 529196 436008 529224
rect 96948 529184 96954 529196
rect 436002 529184 436008 529196
rect 436060 529184 436066 529236
rect 458910 529184 458916 529236
rect 458968 529224 458974 529236
rect 536006 529224 536012 529236
rect 458968 529196 536012 529224
rect 458968 529184 458974 529196
rect 536006 529184 536012 529196
rect 536064 529184 536070 529236
rect 299382 528776 299388 528828
rect 299440 528816 299446 528828
rect 364886 528816 364892 528828
rect 299440 528788 364892 528816
rect 299440 528776 299446 528788
rect 364886 528776 364892 528788
rect 364944 528776 364950 528828
rect 210050 528708 210056 528760
rect 210108 528748 210114 528760
rect 510246 528748 510252 528760
rect 210108 528720 510252 528748
rect 210108 528708 210114 528720
rect 510246 528708 510252 528720
rect 510304 528708 510310 528760
rect 174630 528640 174636 528692
rect 174688 528680 174694 528692
rect 505922 528680 505928 528692
rect 174688 528652 505928 528680
rect 174688 528640 174694 528652
rect 505922 528640 505928 528652
rect 505980 528640 505986 528692
rect 25958 528572 25964 528624
rect 26016 528612 26022 528624
rect 105814 528612 105820 528624
rect 26016 528584 105820 528612
rect 26016 528572 26022 528584
rect 105814 528572 105820 528584
rect 105872 528572 105878 528624
rect 155402 528572 155408 528624
rect 155460 528612 155466 528624
rect 500954 528612 500960 528624
rect 155460 528584 500960 528612
rect 155460 528572 155466 528584
rect 500954 528572 500960 528584
rect 501012 528572 501018 528624
rect 121454 528504 121460 528556
rect 121512 528544 121518 528556
rect 385402 528544 385408 528556
rect 121512 528516 385408 528544
rect 121512 528504 121518 528516
rect 385402 528504 385408 528516
rect 385460 528504 385466 528556
rect 125502 528436 125508 528488
rect 125560 528476 125566 528488
rect 289078 528476 289084 528488
rect 125560 528448 289084 528476
rect 125560 528436 125566 528448
rect 289078 528436 289084 528448
rect 289136 528436 289142 528488
rect 55122 528368 55128 528420
rect 55180 528408 55186 528420
rect 137830 528408 137836 528420
rect 55180 528380 137836 528408
rect 55180 528368 55186 528380
rect 137830 528368 137836 528380
rect 137888 528368 137894 528420
rect 475838 528368 475844 528420
rect 475896 528408 475902 528420
rect 488534 528408 488540 528420
rect 475896 528380 488540 528408
rect 475896 528368 475902 528380
rect 488534 528368 488540 528380
rect 488592 528368 488598 528420
rect 125410 528300 125416 528352
rect 125468 528340 125474 528352
rect 157978 528340 157984 528352
rect 125468 528312 157984 528340
rect 125468 528300 125474 528312
rect 157978 528300 157984 528312
rect 158036 528300 158042 528352
rect 483750 528300 483756 528352
rect 483808 528340 483814 528352
rect 520918 528340 520924 528352
rect 483808 528312 520924 528340
rect 483808 528300 483814 528312
rect 520918 528300 520924 528312
rect 520976 528300 520982 528352
rect 299290 528232 299296 528284
rect 299348 528272 299354 528284
rect 502886 528272 502892 528284
rect 299348 528244 502892 528272
rect 299348 528232 299354 528244
rect 502886 528232 502892 528244
rect 502944 528232 502950 528284
rect 133322 528164 133328 528216
rect 133380 528204 133386 528216
rect 342622 528204 342628 528216
rect 133380 528176 342628 528204
rect 133380 528164 133386 528176
rect 342622 528164 342628 528176
rect 342680 528164 342686 528216
rect 486418 528164 486424 528216
rect 486476 528204 486482 528216
rect 524966 528204 524972 528216
rect 486476 528176 524972 528204
rect 486476 528164 486482 528176
rect 524966 528164 524972 528176
rect 525024 528164 525030 528216
rect 162210 528096 162216 528148
rect 162268 528136 162274 528148
rect 430574 528136 430580 528148
rect 162268 528108 430580 528136
rect 162268 528096 162274 528108
rect 430574 528096 430580 528108
rect 430632 528096 430638 528148
rect 483658 528096 483664 528148
rect 483716 528136 483722 528148
rect 529014 528136 529020 528148
rect 483716 528108 529020 528136
rect 483716 528096 483722 528108
rect 529014 528096 529020 528108
rect 529072 528096 529078 528148
rect 232130 528028 232136 528080
rect 232188 528068 232194 528080
rect 502150 528068 502156 528080
rect 232188 528040 502156 528068
rect 232188 528028 232194 528040
rect 502150 528028 502156 528040
rect 502208 528028 502214 528080
rect 229094 527960 229100 528012
rect 229152 528000 229158 528012
rect 508498 528000 508504 528012
rect 229152 527972 508504 528000
rect 229152 527960 229158 527972
rect 508498 527960 508504 527972
rect 508556 527960 508562 528012
rect 60826 527892 60832 527944
rect 60884 527932 60890 527944
rect 124858 527932 124864 527944
rect 60884 527904 124864 527932
rect 60884 527892 60890 527904
rect 124858 527892 124864 527904
rect 124916 527892 124922 527944
rect 159358 527892 159364 527944
rect 159416 527932 159422 527944
rect 442718 527932 442724 527944
rect 159416 527904 442724 527932
rect 159416 527892 159422 527904
rect 442718 527892 442724 527904
rect 442776 527892 442782 527944
rect 463234 527892 463240 527944
rect 463292 527932 463298 527944
rect 523310 527932 523316 527944
rect 463292 527904 523316 527932
rect 463292 527892 463298 527904
rect 523310 527892 523316 527904
rect 523368 527892 523374 527944
rect 31754 527824 31760 527876
rect 31812 527864 31818 527876
rect 32766 527864 32772 527876
rect 31812 527836 32772 527864
rect 31812 527824 31818 527836
rect 32766 527824 32772 527836
rect 32824 527864 32830 527876
rect 91738 527864 91744 527876
rect 32824 527836 91744 527864
rect 32824 527824 32830 527836
rect 91738 527824 91744 527836
rect 91796 527824 91802 527876
rect 120074 527824 120080 527876
rect 120132 527864 120138 527876
rect 517514 527864 517520 527876
rect 120132 527836 517520 527864
rect 120132 527824 120138 527836
rect 517514 527824 517520 527836
rect 517572 527824 517578 527876
rect 61562 527620 61568 527672
rect 61620 527660 61626 527672
rect 97902 527660 97908 527672
rect 61620 527632 97908 527660
rect 61620 527620 61626 527632
rect 97902 527620 97908 527632
rect 97960 527620 97966 527672
rect 124122 527620 124128 527672
rect 124180 527660 124186 527672
rect 231762 527660 231768 527672
rect 124180 527632 231768 527660
rect 124180 527620 124186 527632
rect 231762 527620 231768 527632
rect 231820 527620 231826 527672
rect 59814 527552 59820 527604
rect 59872 527592 59878 527604
rect 123938 527592 123944 527604
rect 59872 527564 123944 527592
rect 59872 527552 59878 527564
rect 123938 527552 123944 527564
rect 123996 527552 124002 527604
rect 59262 527484 59268 527536
rect 59320 527524 59326 527536
rect 126974 527524 126980 527536
rect 59320 527496 126980 527524
rect 59320 527484 59326 527496
rect 126974 527484 126980 527496
rect 127032 527484 127038 527536
rect 60550 527416 60556 527468
rect 60608 527456 60614 527468
rect 125042 527456 125048 527468
rect 60608 527428 125048 527456
rect 60608 527416 60614 527428
rect 125042 527416 125048 527428
rect 125100 527416 125106 527468
rect 61654 527348 61660 527400
rect 61712 527388 61718 527400
rect 132034 527388 132040 527400
rect 61712 527360 132040 527388
rect 61712 527348 61718 527360
rect 132034 527348 132040 527360
rect 132092 527348 132098 527400
rect 202046 527348 202052 527400
rect 202104 527388 202110 527400
rect 511994 527388 512000 527400
rect 202104 527360 512000 527388
rect 202104 527348 202110 527360
rect 511994 527348 512000 527360
rect 512052 527348 512058 527400
rect 50982 527280 50988 527332
rect 51040 527320 51046 527332
rect 122926 527320 122932 527332
rect 51040 527292 122932 527320
rect 51040 527280 51046 527292
rect 122926 527280 122932 527292
rect 122984 527280 122990 527332
rect 204162 527280 204168 527332
rect 204220 527320 204226 527332
rect 514754 527320 514760 527332
rect 204220 527292 514760 527320
rect 204220 527280 204226 527292
rect 514754 527280 514760 527292
rect 514812 527280 514818 527332
rect 53466 527212 53472 527264
rect 53524 527252 53530 527264
rect 136174 527252 136180 527264
rect 53524 527224 136180 527252
rect 53524 527212 53530 527224
rect 136174 527212 136180 527224
rect 136232 527212 136238 527264
rect 177758 527212 177764 527264
rect 177816 527252 177822 527264
rect 523034 527252 523040 527264
rect 177816 527224 523040 527252
rect 177816 527212 177822 527224
rect 523034 527212 523040 527224
rect 523092 527212 523098 527264
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 31754 527184 31760 527196
rect 3476 527156 31760 527184
rect 3476 527144 3482 527156
rect 31754 527144 31760 527156
rect 31812 527144 31818 527196
rect 46750 527144 46756 527196
rect 46808 527184 46814 527196
rect 130102 527184 130108 527196
rect 46808 527156 130108 527184
rect 46808 527144 46814 527156
rect 130102 527144 130108 527156
rect 130160 527144 130166 527196
rect 189902 527144 189908 527196
rect 189960 527184 189966 527196
rect 545114 527184 545120 527196
rect 189960 527156 545120 527184
rect 189960 527144 189966 527156
rect 545114 527144 545120 527156
rect 545172 527144 545178 527196
rect 62022 527076 62028 527128
rect 62080 527116 62086 527128
rect 365254 527116 365260 527128
rect 62080 527088 365260 527116
rect 62080 527076 62086 527088
rect 365254 527076 365260 527088
rect 365312 527076 365318 527128
rect 111794 527008 111800 527060
rect 111852 527048 111858 527060
rect 341978 527048 341984 527060
rect 111852 527020 341984 527048
rect 111852 527008 111858 527020
rect 341978 527008 341984 527020
rect 342036 527008 342042 527060
rect 178034 526940 178040 526992
rect 178092 526980 178098 526992
rect 374454 526980 374460 526992
rect 178092 526952 374460 526980
rect 178092 526940 178098 526952
rect 374454 526940 374460 526952
rect 374512 526940 374518 526992
rect 214558 526872 214564 526924
rect 214616 526912 214622 526924
rect 385310 526912 385316 526924
rect 214616 526884 385316 526912
rect 214616 526872 214622 526884
rect 385310 526872 385316 526884
rect 385368 526872 385374 526924
rect 233878 526804 233884 526856
rect 233936 526844 233942 526856
rect 383746 526844 383752 526856
rect 233936 526816 383752 526844
rect 233936 526804 233942 526816
rect 383746 526804 383752 526816
rect 383804 526804 383810 526856
rect 106182 526736 106188 526788
rect 106240 526776 106246 526788
rect 254670 526776 254676 526788
rect 106240 526748 254676 526776
rect 106240 526736 106246 526748
rect 254670 526736 254676 526748
rect 254728 526736 254734 526788
rect 249702 526668 249708 526720
rect 249760 526708 249766 526720
rect 286318 526708 286324 526720
rect 249760 526680 286324 526708
rect 249760 526668 249766 526680
rect 286318 526668 286324 526680
rect 286376 526668 286382 526720
rect 501782 526668 501788 526720
rect 501840 526708 501846 526720
rect 517514 526708 517520 526720
rect 501840 526680 517520 526708
rect 501840 526668 501846 526680
rect 517514 526668 517520 526680
rect 517572 526668 517578 526720
rect 483842 526600 483848 526652
rect 483900 526640 483906 526652
rect 527910 526640 527916 526652
rect 483900 526612 527916 526640
rect 483900 526600 483906 526612
rect 527910 526600 527916 526612
rect 527968 526600 527974 526652
rect 485130 526532 485136 526584
rect 485188 526572 485194 526584
rect 534442 526572 534448 526584
rect 485188 526544 534448 526572
rect 485188 526532 485194 526544
rect 534442 526532 534448 526544
rect 534500 526532 534506 526584
rect 462958 526464 462964 526516
rect 463016 526504 463022 526516
rect 513650 526504 513656 526516
rect 463016 526476 513656 526504
rect 463016 526464 463022 526476
rect 513650 526464 513656 526476
rect 513708 526464 513714 526516
rect 59446 526396 59452 526448
rect 59504 526436 59510 526448
rect 135898 526436 135904 526448
rect 59504 526408 135904 526436
rect 59504 526396 59510 526408
rect 135898 526396 135904 526408
rect 135956 526396 135962 526448
rect 176838 526396 176844 526448
rect 176896 526436 176902 526448
rect 285766 526436 285772 526448
rect 176896 526408 285772 526436
rect 176896 526396 176902 526408
rect 285766 526396 285772 526408
rect 285824 526396 285830 526448
rect 287698 526396 287704 526448
rect 287756 526436 287762 526448
rect 522390 526436 522396 526448
rect 287756 526408 522396 526436
rect 287756 526396 287762 526408
rect 522390 526396 522396 526408
rect 522448 526396 522454 526448
rect 59722 526328 59728 526380
rect 59780 526368 59786 526380
rect 112898 526368 112904 526380
rect 59780 526340 112904 526368
rect 59780 526328 59786 526340
rect 112898 526328 112904 526340
rect 112956 526328 112962 526380
rect 61838 526260 61844 526312
rect 61896 526300 61902 526312
rect 114922 526300 114928 526312
rect 61896 526272 114928 526300
rect 61896 526260 61902 526272
rect 114922 526260 114928 526272
rect 114980 526260 114986 526312
rect 47946 526192 47952 526244
rect 48004 526232 48010 526244
rect 109770 526232 109776 526244
rect 48004 526204 109776 526232
rect 48004 526192 48010 526204
rect 109770 526192 109776 526204
rect 109828 526192 109834 526244
rect 288342 526192 288348 526244
rect 288400 526232 288406 526244
rect 501690 526232 501696 526244
rect 288400 526204 501696 526232
rect 288400 526192 288406 526204
rect 501690 526192 501696 526204
rect 501748 526192 501754 526244
rect 46658 526124 46664 526176
rect 46716 526164 46722 526176
rect 108758 526164 108764 526176
rect 46716 526136 108764 526164
rect 46716 526124 46722 526136
rect 108758 526124 108764 526136
rect 108816 526124 108822 526176
rect 152550 526124 152556 526176
rect 152608 526164 152614 526176
rect 247034 526164 247040 526176
rect 152608 526136 247040 526164
rect 152608 526124 152614 526136
rect 247034 526124 247040 526136
rect 247092 526124 247098 526176
rect 256694 526124 256700 526176
rect 256752 526164 256758 526176
rect 499942 526164 499948 526176
rect 256752 526136 499948 526164
rect 256752 526124 256758 526136
rect 499942 526124 499948 526136
rect 500000 526124 500006 526176
rect 25774 526056 25780 526108
rect 25832 526096 25838 526108
rect 95602 526096 95608 526108
rect 25832 526068 95608 526096
rect 25832 526056 25838 526068
rect 95602 526056 95608 526068
rect 95660 526056 95666 526108
rect 237466 526056 237472 526108
rect 237524 526096 237530 526108
rect 515214 526096 515220 526108
rect 237524 526068 515220 526096
rect 237524 526056 237530 526068
rect 515214 526056 515220 526068
rect 515272 526056 515278 526108
rect 39942 525988 39948 526040
rect 40000 526028 40006 526040
rect 110782 526028 110788 526040
rect 40000 526000 110788 526028
rect 40000 525988 40006 526000
rect 110782 525988 110788 526000
rect 110840 525988 110846 526040
rect 200022 525988 200028 526040
rect 200080 526028 200086 526040
rect 498194 526028 498200 526040
rect 200080 526000 498200 526028
rect 200080 525988 200086 526000
rect 498194 525988 498200 526000
rect 498252 525988 498258 526040
rect 40954 525920 40960 525972
rect 41012 525960 41018 525972
rect 116854 525960 116860 525972
rect 41012 525932 116860 525960
rect 41012 525920 41018 525932
rect 116854 525920 116860 525932
rect 116912 525920 116918 525972
rect 198090 525920 198096 525972
rect 198148 525960 198154 525972
rect 510614 525960 510620 525972
rect 198148 525932 510620 525960
rect 198148 525920 198154 525932
rect 510614 525920 510620 525932
rect 510672 525920 510678 525972
rect 58618 525852 58624 525904
rect 58676 525892 58682 525904
rect 143258 525892 143264 525904
rect 58676 525864 143264 525892
rect 58676 525852 58682 525864
rect 143258 525852 143264 525864
rect 143316 525852 143322 525904
rect 173802 525852 173808 525904
rect 173860 525892 173866 525904
rect 519078 525892 519084 525904
rect 173860 525864 519084 525892
rect 173860 525852 173866 525864
rect 519078 525852 519084 525864
rect 519136 525852 519142 525904
rect 60366 525784 60372 525836
rect 60424 525824 60430 525836
rect 63402 525824 63408 525836
rect 60424 525796 63408 525824
rect 60424 525784 60430 525796
rect 63402 525784 63408 525796
rect 63460 525784 63466 525836
rect 82722 525784 82728 525836
rect 82780 525824 82786 525836
rect 516318 525824 516324 525836
rect 82780 525796 516324 525824
rect 82780 525784 82786 525796
rect 516318 525784 516324 525796
rect 516376 525784 516382 525836
rect 69014 525716 69020 525768
rect 69072 525756 69078 525768
rect 386414 525756 386420 525768
rect 69072 525728 386420 525756
rect 69072 525716 69078 525728
rect 386414 525716 386420 525728
rect 386472 525716 386478 525768
rect 70394 525648 70400 525700
rect 70452 525688 70458 525700
rect 382458 525688 382464 525700
rect 70452 525660 382464 525688
rect 70452 525648 70458 525660
rect 382458 525648 382464 525660
rect 382516 525648 382522 525700
rect 247034 525580 247040 525632
rect 247092 525620 247098 525632
rect 511994 525620 512000 525632
rect 247092 525592 512000 525620
rect 247092 525580 247098 525592
rect 511994 525580 512000 525592
rect 512052 525580 512058 525632
rect 117958 525512 117964 525564
rect 118016 525552 118022 525564
rect 379606 525552 379612 525564
rect 118016 525524 379612 525552
rect 118016 525512 118022 525524
rect 379606 525512 379612 525524
rect 379664 525512 379670 525564
rect 247034 525444 247040 525496
rect 247092 525484 247098 525496
rect 379698 525484 379704 525496
rect 247092 525456 379704 525484
rect 247092 525444 247098 525456
rect 379698 525444 379704 525456
rect 379756 525444 379762 525496
rect 498654 525444 498660 525496
rect 498712 525484 498718 525496
rect 499114 525484 499120 525496
rect 498712 525456 499120 525484
rect 498712 525444 498718 525456
rect 499114 525444 499120 525456
rect 499172 525444 499178 525496
rect 224954 525376 224960 525428
rect 225012 525416 225018 525428
rect 308582 525416 308588 525428
rect 225012 525388 308588 525416
rect 225012 525376 225018 525388
rect 308582 525376 308588 525388
rect 308640 525376 308646 525428
rect 478138 525376 478144 525428
rect 478196 525416 478202 525428
rect 519630 525416 519636 525428
rect 478196 525388 519636 525416
rect 478196 525376 478202 525388
rect 519630 525376 519636 525388
rect 519688 525376 519694 525428
rect 482554 525308 482560 525360
rect 482612 525348 482618 525360
rect 527818 525348 527824 525360
rect 482612 525320 527824 525348
rect 482612 525308 482618 525320
rect 527818 525308 527824 525320
rect 527876 525308 527882 525360
rect 472710 525240 472716 525292
rect 472768 525280 472774 525292
rect 525058 525280 525064 525292
rect 472768 525252 525064 525280
rect 472768 525240 472774 525252
rect 525058 525240 525064 525252
rect 525116 525240 525122 525292
rect 186866 525172 186872 525224
rect 186924 525212 186930 525224
rect 253198 525212 253204 525224
rect 186924 525184 253204 525212
rect 186924 525172 186930 525184
rect 253198 525172 253204 525184
rect 253256 525172 253262 525224
rect 469950 525172 469956 525224
rect 470008 525212 470014 525224
rect 529290 525212 529296 525224
rect 470008 525184 529296 525212
rect 470008 525172 470014 525184
rect 529290 525172 529296 525184
rect 529348 525172 529354 525224
rect 159634 525104 159640 525156
rect 159692 525144 159698 525156
rect 246298 525144 246304 525156
rect 159692 525116 246304 525144
rect 159692 525104 159698 525116
rect 246298 525104 246304 525116
rect 246356 525104 246362 525156
rect 467098 525104 467104 525156
rect 467156 525144 467162 525156
rect 529106 525144 529112 525156
rect 467156 525116 529112 525144
rect 467156 525104 467162 525116
rect 529106 525104 529112 525116
rect 529164 525104 529170 525156
rect 53190 525036 53196 525088
rect 53248 525076 53254 525088
rect 349062 525076 349068 525088
rect 53248 525048 349068 525076
rect 53248 525036 53254 525048
rect 349062 525036 349068 525048
rect 349120 525036 349126 525088
rect 453298 525036 453304 525088
rect 453356 525076 453362 525088
rect 526346 525076 526352 525088
rect 453356 525048 526352 525076
rect 453356 525036 453362 525048
rect 526346 525036 526352 525048
rect 526404 525036 526410 525088
rect 29914 524968 29920 525020
rect 29972 525008 29978 525020
rect 97718 525008 97724 525020
rect 29972 524980 97724 525008
rect 29972 524968 29978 524980
rect 97718 524968 97724 524980
rect 97776 524968 97782 525020
rect 60734 524900 60740 524952
rect 60792 524940 60798 524952
rect 71958 524940 71964 524952
rect 60792 524912 71964 524940
rect 60792 524900 60798 524912
rect 71958 524900 71964 524912
rect 72016 524900 72022 524952
rect 62022 524832 62028 524884
rect 62080 524872 62086 524884
rect 122006 524872 122012 524884
rect 62080 524844 122012 524872
rect 62080 524832 62086 524844
rect 122006 524832 122012 524844
rect 122064 524832 122070 524884
rect 41046 524764 41052 524816
rect 41104 524804 41110 524816
rect 101674 524804 101680 524816
rect 41104 524776 101680 524804
rect 41104 524764 41110 524776
rect 101674 524764 101680 524776
rect 101732 524764 101738 524816
rect 285674 524764 285680 524816
rect 285732 524804 285738 524816
rect 505186 524804 505192 524816
rect 285732 524776 505192 524804
rect 285732 524764 285738 524776
rect 505186 524764 505192 524776
rect 505244 524764 505250 524816
rect 29822 524696 29828 524748
rect 29880 524736 29886 524748
rect 99742 524736 99748 524748
rect 29880 524708 99748 524736
rect 29880 524696 29886 524708
rect 99742 524696 99748 524708
rect 99800 524696 99806 524748
rect 222378 524696 222384 524748
rect 222436 524736 222442 524748
rect 525794 524736 525800 524748
rect 222436 524708 525800 524736
rect 222436 524696 222442 524708
rect 525794 524696 525800 524708
rect 525852 524696 525858 524748
rect 31478 524628 31484 524680
rect 31536 524668 31542 524680
rect 102686 524668 102692 524680
rect 31536 524640 102692 524668
rect 31536 524628 31542 524640
rect 102686 524628 102692 524640
rect 102744 524628 102750 524680
rect 197078 524628 197084 524680
rect 197136 524668 197142 524680
rect 500862 524668 500868 524680
rect 197136 524640 500868 524668
rect 197136 524628 197142 524640
rect 500862 524628 500868 524640
rect 500920 524628 500926 524680
rect 27338 524560 27344 524612
rect 27396 524600 27402 524612
rect 100754 524600 100760 524612
rect 27396 524572 100760 524600
rect 27396 524560 27402 524572
rect 100754 524560 100760 524572
rect 100812 524560 100818 524612
rect 201034 524560 201040 524612
rect 201092 524600 201098 524612
rect 509878 524600 509884 524612
rect 201092 524572 509884 524600
rect 201092 524560 201098 524572
rect 509878 524560 509884 524572
rect 509936 524560 509942 524612
rect 44174 524492 44180 524544
rect 44232 524532 44238 524544
rect 144822 524532 144828 524544
rect 44232 524504 144828 524532
rect 44232 524492 44238 524504
rect 144822 524492 144828 524504
rect 144880 524492 144886 524544
rect 177942 524492 177948 524544
rect 178000 524532 178006 524544
rect 507210 524532 507216 524544
rect 178000 524504 507216 524532
rect 178000 524492 178006 524504
rect 507210 524492 507216 524504
rect 507268 524492 507274 524544
rect 54570 524424 54576 524476
rect 54628 524464 54634 524476
rect 71866 524464 71872 524476
rect 54628 524436 71872 524464
rect 54628 524424 54634 524436
rect 71866 524424 71872 524436
rect 71924 524424 71930 524476
rect 87690 524424 87696 524476
rect 87748 524464 87754 524476
rect 519262 524464 519268 524476
rect 87748 524436 519268 524464
rect 87748 524424 87754 524436
rect 519262 524424 519268 524436
rect 519320 524424 519326 524476
rect 57698 524356 57704 524408
rect 57756 524396 57762 524408
rect 378870 524396 378876 524408
rect 57756 524368 378876 524396
rect 57756 524356 57762 524368
rect 378870 524356 378876 524368
rect 378928 524356 378934 524408
rect 68922 524288 68928 524340
rect 68980 524328 68986 524340
rect 385218 524328 385224 524340
rect 68980 524300 385224 524328
rect 68980 524288 68986 524300
rect 385218 524288 385224 524300
rect 385276 524288 385282 524340
rect 78582 524220 78588 524272
rect 78640 524260 78646 524272
rect 383654 524260 383660 524272
rect 78640 524232 383660 524260
rect 78640 524220 78646 524232
rect 383654 524220 383660 524232
rect 383712 524220 383718 524272
rect 53834 524152 53840 524204
rect 53892 524192 53898 524204
rect 351086 524192 351092 524204
rect 53892 524164 351092 524192
rect 53892 524152 53898 524164
rect 351086 524152 351092 524164
rect 351144 524152 351150 524204
rect 241330 524084 241336 524136
rect 241388 524124 241394 524136
rect 382642 524124 382648 524136
rect 241388 524096 382648 524124
rect 241388 524084 241394 524096
rect 382642 524084 382648 524096
rect 382700 524084 382706 524136
rect 470042 523880 470048 523932
rect 470100 523920 470106 523932
rect 515582 523920 515588 523932
rect 470100 523892 515588 523920
rect 470100 523880 470106 523892
rect 515582 523880 515588 523892
rect 515640 523880 515646 523932
rect 480990 523812 480996 523864
rect 481048 523852 481054 523864
rect 530486 523852 530492 523864
rect 481048 523824 530492 523852
rect 481048 523812 481054 523824
rect 530486 523812 530492 523824
rect 530544 523812 530550 523864
rect 489178 523744 489184 523796
rect 489236 523784 489242 523796
rect 541618 523784 541624 523796
rect 489236 523756 541624 523784
rect 489236 523744 489242 523756
rect 541618 523744 541624 523756
rect 541676 523744 541682 523796
rect 27522 523676 27528 523728
rect 27580 523716 27586 523728
rect 44174 523716 44180 523728
rect 27580 523688 44180 523716
rect 27580 523676 27586 523688
rect 44174 523676 44180 523688
rect 44232 523676 44238 523728
rect 58894 523676 58900 523728
rect 58952 523716 58958 523728
rect 356146 523716 356152 523728
rect 58952 523688 356152 523716
rect 58952 523676 58958 523688
rect 356146 523676 356152 523688
rect 356204 523676 356210 523728
rect 456058 523676 456064 523728
rect 456116 523716 456122 523728
rect 533154 523716 533160 523728
rect 456116 523688 533160 523716
rect 456116 523676 456122 523688
rect 533154 523676 533160 523688
rect 533212 523676 533218 523728
rect 500310 523608 500316 523660
rect 500368 523648 500374 523660
rect 505830 523648 505836 523660
rect 500368 523620 505836 523648
rect 500368 523608 500374 523620
rect 505830 523608 505836 523620
rect 505888 523608 505894 523660
rect 510154 523608 510160 523660
rect 510212 523648 510218 523660
rect 511258 523648 511264 523660
rect 510212 523620 511264 523648
rect 510212 523608 510218 523620
rect 511258 523608 511264 523620
rect 511316 523608 511322 523660
rect 50798 523540 50804 523592
rect 50856 523580 50862 523592
rect 69658 523580 69664 523592
rect 50856 523552 69664 523580
rect 50856 523540 50862 523552
rect 69658 523540 69664 523552
rect 69716 523540 69722 523592
rect 489886 523552 491294 523580
rect 26878 523472 26884 523524
rect 26936 523512 26942 523524
rect 129734 523512 129740 523524
rect 26936 523484 129740 523512
rect 26936 523472 26942 523484
rect 129734 523472 129740 523484
rect 129792 523472 129798 523524
rect 177942 523472 177948 523524
rect 178000 523512 178006 523524
rect 489886 523512 489914 523552
rect 178000 523484 489914 523512
rect 491266 523512 491294 523552
rect 500310 523512 500316 523524
rect 491266 523484 500316 523512
rect 178000 523472 178006 523484
rect 500310 523472 500316 523484
rect 500368 523472 500374 523524
rect 55858 523404 55864 523456
rect 55916 523444 55922 523456
rect 71774 523444 71780 523456
rect 55916 523416 71780 523444
rect 55916 523404 55922 523416
rect 71774 523404 71780 523416
rect 71832 523404 71838 523456
rect 481542 523404 481548 523456
rect 481600 523444 481606 523456
rect 522114 523444 522120 523456
rect 481600 523416 522120 523444
rect 481600 523404 481606 523416
rect 522114 523404 522120 523416
rect 522172 523404 522178 523456
rect 42426 523336 42432 523388
rect 42484 523376 42490 523388
rect 103790 523376 103796 523388
rect 42484 523348 103796 523376
rect 42484 523336 42490 523348
rect 103790 523336 103796 523348
rect 103848 523336 103854 523388
rect 203058 523336 203064 523388
rect 203116 523376 203122 523388
rect 500034 523376 500040 523388
rect 203116 523348 500040 523376
rect 203116 523336 203122 523348
rect 500034 523336 500040 523348
rect 500092 523336 500098 523388
rect 500402 523336 500408 523388
rect 500460 523376 500466 523388
rect 503714 523376 503720 523388
rect 500460 523348 503720 523376
rect 500460 523336 500466 523348
rect 503714 523336 503720 523348
rect 503772 523336 503778 523388
rect 29730 523268 29736 523320
rect 29788 523308 29794 523320
rect 98730 523308 98736 523320
rect 29788 523280 98736 523308
rect 29788 523268 29794 523280
rect 98730 523268 98736 523280
rect 98788 523268 98794 523320
rect 223298 523268 223304 523320
rect 223356 523308 223362 523320
rect 525794 523308 525800 523320
rect 223356 523280 525800 523308
rect 223356 523268 223362 523280
rect 525794 523268 525800 523280
rect 525852 523268 525858 523320
rect 28626 523200 28632 523252
rect 28684 523240 28690 523252
rect 104710 523240 104716 523252
rect 28684 523212 104716 523240
rect 28684 523200 28690 523212
rect 104710 523200 104716 523212
rect 104768 523200 104774 523252
rect 206186 523200 206192 523252
rect 206244 523240 206250 523252
rect 516870 523240 516876 523252
rect 206244 523212 516876 523240
rect 206244 523200 206250 523212
rect 516870 523200 516876 523212
rect 516928 523200 516934 523252
rect 60734 523132 60740 523184
rect 60792 523172 60798 523184
rect 139394 523172 139400 523184
rect 60792 523144 139400 523172
rect 60792 523132 60798 523144
rect 139394 523132 139400 523144
rect 139452 523132 139458 523184
rect 496722 523132 496728 523184
rect 496780 523172 496786 523184
rect 545206 523172 545212 523184
rect 496780 523144 545212 523172
rect 496780 523132 496786 523144
rect 545206 523132 545212 523144
rect 545264 523132 545270 523184
rect 25590 523064 25596 523116
rect 25648 523104 25654 523116
rect 117866 523104 117872 523116
rect 25648 523076 117872 523104
rect 25648 523064 25654 523076
rect 117866 523064 117872 523076
rect 117924 523064 117930 523116
rect 182910 523064 182916 523116
rect 182968 523104 182974 523116
rect 528554 523104 528560 523116
rect 182968 523076 528560 523104
rect 182968 523064 182974 523076
rect 528554 523064 528560 523076
rect 528612 523064 528618 523116
rect 52546 522996 52552 523048
rect 52604 523036 52610 523048
rect 68922 523036 68928 523048
rect 52604 523008 68928 523036
rect 52604 522996 52610 523008
rect 68922 522996 68928 523008
rect 68980 522996 68986 523048
rect 171686 522996 171692 523048
rect 171744 523036 171750 523048
rect 518066 523036 518072 523048
rect 171744 523008 518072 523036
rect 171744 522996 171750 523008
rect 518066 522996 518072 523008
rect 518124 522996 518130 523048
rect 59538 522928 59544 522980
rect 59596 522968 59602 522980
rect 60826 522968 60832 522980
rect 59596 522940 60832 522968
rect 59596 522928 59602 522940
rect 60826 522928 60832 522940
rect 60884 522928 60890 522980
rect 178034 522928 178040 522980
rect 178092 522968 178098 522980
rect 378226 522968 378232 522980
rect 178092 522940 378232 522968
rect 178092 522928 178098 522940
rect 378226 522928 378232 522940
rect 378284 522928 378290 522980
rect 395338 522928 395344 522980
rect 395396 522968 395402 522980
rect 396166 522968 396172 522980
rect 395396 522940 396172 522968
rect 395396 522928 395402 522940
rect 396166 522928 396172 522940
rect 396224 522928 396230 522980
rect 400858 522928 400864 522980
rect 400916 522968 400922 522980
rect 402330 522968 402336 522980
rect 400916 522940 402336 522968
rect 400916 522928 400922 522940
rect 402330 522928 402336 522940
rect 402388 522928 402394 522980
rect 403618 522928 403624 522980
rect 403676 522968 403682 522980
rect 404262 522968 404268 522980
rect 403676 522940 404268 522968
rect 403676 522928 403682 522940
rect 404262 522928 404268 522940
rect 404320 522928 404326 522980
rect 407758 522928 407764 522980
rect 407816 522968 407822 522980
rect 410426 522968 410432 522980
rect 407816 522940 410432 522968
rect 407816 522928 407822 522940
rect 410426 522928 410432 522940
rect 410484 522928 410490 522980
rect 410518 522928 410524 522980
rect 410576 522968 410582 522980
rect 413370 522968 413376 522980
rect 410576 522940 413376 522968
rect 410576 522928 410582 522940
rect 413370 522928 413376 522940
rect 413428 522928 413434 522980
rect 414658 522928 414664 522980
rect 414716 522968 414722 522980
rect 415486 522968 415492 522980
rect 414716 522940 415492 522968
rect 414716 522928 414722 522940
rect 415486 522928 415492 522940
rect 415544 522928 415550 522980
rect 500218 522928 500224 522980
rect 500276 522968 500282 522980
rect 500402 522968 500408 522980
rect 500276 522940 500408 522968
rect 500276 522928 500282 522940
rect 500402 522928 500408 522940
rect 500460 522928 500466 522980
rect 184842 522860 184848 522912
rect 184900 522900 184906 522912
rect 369118 522900 369124 522912
rect 184900 522872 369124 522900
rect 184900 522860 184906 522872
rect 369118 522860 369124 522872
rect 369176 522860 369182 522912
rect 373258 522860 373264 522912
rect 373316 522900 373322 522912
rect 373994 522900 374000 522912
rect 373316 522872 374000 522900
rect 373316 522860 373322 522872
rect 373994 522860 374000 522872
rect 374052 522860 374058 522912
rect 488534 522860 488540 522912
rect 488592 522900 488598 522912
rect 497366 522900 497372 522912
rect 488592 522872 497372 522900
rect 488592 522860 488598 522872
rect 497366 522860 497372 522872
rect 497424 522860 497430 522912
rect 224126 522792 224132 522844
rect 224184 522832 224190 522844
rect 385034 522832 385040 522844
rect 224184 522804 385040 522832
rect 224184 522792 224190 522804
rect 385034 522792 385040 522804
rect 385092 522792 385098 522844
rect 475654 522792 475660 522844
rect 475712 522832 475718 522844
rect 518066 522832 518072 522844
rect 475712 522804 518072 522832
rect 475712 522792 475718 522804
rect 518066 522792 518072 522804
rect 518124 522792 518130 522844
rect 227714 522724 227720 522776
rect 227772 522764 227778 522776
rect 386690 522764 386696 522776
rect 227772 522736 386696 522764
rect 227772 522724 227778 522736
rect 386690 522724 386696 522736
rect 386748 522724 386754 522776
rect 436002 522724 436008 522776
rect 436060 522764 436066 522776
rect 491294 522764 491300 522776
rect 436060 522736 491300 522764
rect 436060 522724 436066 522736
rect 491294 522724 491300 522736
rect 491352 522724 491358 522776
rect 226334 522656 226340 522708
rect 226392 522696 226398 522708
rect 382550 522696 382556 522708
rect 226392 522668 382556 522696
rect 226392 522656 226398 522668
rect 382550 522656 382556 522668
rect 382608 522656 382614 522708
rect 391290 522656 391296 522708
rect 391348 522696 391354 522708
rect 408402 522696 408408 522708
rect 391348 522668 408408 522696
rect 391348 522656 391354 522668
rect 408402 522656 408408 522668
rect 408460 522656 408466 522708
rect 418798 522656 418804 522708
rect 418856 522696 418862 522708
rect 489270 522696 489276 522708
rect 418856 522668 489276 522696
rect 418856 522656 418862 522668
rect 489270 522656 489276 522668
rect 489328 522656 489334 522708
rect 496078 522656 496084 522708
rect 496136 522696 496142 522708
rect 505278 522696 505284 522708
rect 496136 522668 505284 522696
rect 496136 522656 496142 522668
rect 505278 522656 505284 522668
rect 505336 522656 505342 522708
rect 42334 522588 42340 522640
rect 42392 522628 42398 522640
rect 70394 522628 70400 522640
rect 42392 522600 70400 522628
rect 42392 522588 42398 522600
rect 70394 522588 70400 522600
rect 70452 522588 70458 522640
rect 347130 522588 347136 522640
rect 347188 522628 347194 522640
rect 476114 522628 476120 522640
rect 347188 522600 476120 522628
rect 347188 522588 347194 522600
rect 476114 522588 476120 522600
rect 476172 522588 476178 522640
rect 496262 522588 496268 522640
rect 496320 522628 496326 522640
rect 513374 522628 513380 522640
rect 496320 522600 513380 522628
rect 496320 522588 496326 522600
rect 513374 522588 513380 522600
rect 513432 522588 513438 522640
rect 43898 522520 43904 522572
rect 43956 522560 43962 522572
rect 69382 522560 69388 522572
rect 43956 522532 69388 522560
rect 43956 522520 43962 522532
rect 69382 522520 69388 522532
rect 69440 522520 69446 522572
rect 69658 522520 69664 522572
rect 69716 522560 69722 522572
rect 111794 522560 111800 522572
rect 69716 522532 111800 522560
rect 69716 522520 69722 522532
rect 111794 522520 111800 522532
rect 111852 522520 111858 522572
rect 313182 522520 313188 522572
rect 313240 522560 313246 522572
rect 474090 522560 474096 522572
rect 313240 522532 474096 522560
rect 313240 522520 313246 522532
rect 474090 522520 474096 522532
rect 474148 522520 474154 522572
rect 475470 522520 475476 522572
rect 475528 522560 475534 522572
rect 522206 522560 522212 522572
rect 475528 522532 522212 522560
rect 475528 522520 475534 522532
rect 522206 522520 522212 522532
rect 522264 522520 522270 522572
rect 97902 522452 97908 522504
rect 97960 522492 97966 522504
rect 153378 522492 153384 522504
rect 97960 522464 153384 522492
rect 97960 522452 97966 522464
rect 153378 522452 153384 522464
rect 153436 522452 153442 522504
rect 174906 522452 174912 522504
rect 174964 522492 174970 522504
rect 337470 522492 337476 522504
rect 174964 522464 337476 522492
rect 174964 522452 174970 522464
rect 337470 522452 337476 522464
rect 337528 522452 337534 522504
rect 342898 522452 342904 522504
rect 342956 522492 342962 522504
rect 480254 522492 480260 522504
rect 342956 522464 480260 522492
rect 342956 522452 342962 522464
rect 480254 522452 480260 522464
rect 480312 522452 480318 522504
rect 482370 522452 482376 522504
rect 482428 522492 482434 522504
rect 516778 522492 516784 522504
rect 482428 522464 516784 522492
rect 482428 522452 482434 522464
rect 516778 522452 516784 522464
rect 516836 522452 516842 522504
rect 52822 522384 52828 522436
rect 52880 522424 52886 522436
rect 59814 522424 59820 522436
rect 52880 522396 59820 522424
rect 52880 522384 52886 522396
rect 59814 522384 59820 522396
rect 59872 522384 59878 522436
rect 68922 522384 68928 522436
rect 68980 522424 68986 522436
rect 118878 522424 118884 522436
rect 68980 522396 118884 522424
rect 68980 522384 68986 522396
rect 118878 522384 118884 522396
rect 118936 522384 118942 522436
rect 129734 522384 129740 522436
rect 129792 522424 129798 522436
rect 142154 522424 142160 522436
rect 129792 522396 142160 522424
rect 129792 522384 129798 522396
rect 142154 522384 142160 522396
rect 142212 522384 142218 522436
rect 150342 522384 150348 522436
rect 150400 522424 150406 522436
rect 251818 522424 251824 522436
rect 150400 522396 251824 522424
rect 150400 522384 150406 522396
rect 251818 522384 251824 522396
rect 251876 522384 251882 522436
rect 271138 522384 271144 522436
rect 271196 522424 271202 522436
rect 435726 522424 435732 522436
rect 271196 522396 435732 522424
rect 271196 522384 271202 522396
rect 435726 522384 435732 522396
rect 435784 522384 435790 522436
rect 472802 522384 472808 522436
rect 472860 522424 472866 522436
rect 521010 522424 521016 522436
rect 472860 522396 521016 522424
rect 472860 522384 472866 522396
rect 521010 522384 521016 522396
rect 521068 522384 521074 522436
rect 52454 522316 52460 522368
rect 52512 522356 52518 522368
rect 60734 522356 60740 522368
rect 52512 522328 60740 522356
rect 52512 522316 52518 522328
rect 60734 522316 60740 522328
rect 60792 522316 60798 522368
rect 89622 522316 89628 522368
rect 89680 522356 89686 522368
rect 254854 522356 254860 522368
rect 89680 522328 254860 522356
rect 89680 522316 89686 522328
rect 254854 522316 254860 522328
rect 254912 522316 254918 522368
rect 258994 522316 259000 522368
rect 259052 522356 259058 522368
rect 456978 522356 456984 522368
rect 259052 522328 456984 522356
rect 259052 522316 259058 522328
rect 456978 522316 456984 522328
rect 457036 522316 457042 522368
rect 472618 522316 472624 522368
rect 472676 522356 472682 522368
rect 526530 522356 526536 522368
rect 472676 522328 526536 522356
rect 472676 522316 472682 522328
rect 526530 522316 526536 522328
rect 526588 522316 526594 522368
rect 27154 522248 27160 522300
rect 27212 522288 27218 522300
rect 41414 522288 41420 522300
rect 27212 522260 41420 522288
rect 27212 522248 27218 522260
rect 41414 522248 41420 522260
rect 41472 522248 41478 522300
rect 43806 522248 43812 522300
rect 43864 522288 43870 522300
rect 67358 522288 67364 522300
rect 43864 522260 67364 522288
rect 43864 522248 43870 522260
rect 67358 522248 67364 522260
rect 67416 522248 67422 522300
rect 71774 522248 71780 522300
rect 71832 522288 71838 522300
rect 139210 522288 139216 522300
rect 71832 522260 139216 522288
rect 71832 522248 71838 522260
rect 139210 522248 139216 522260
rect 139268 522248 139274 522300
rect 139394 522248 139400 522300
rect 139452 522288 139458 522300
rect 157334 522288 157340 522300
rect 139452 522260 157340 522288
rect 139452 522248 139458 522260
rect 157334 522248 157340 522260
rect 157392 522248 157398 522300
rect 170858 522248 170864 522300
rect 170916 522288 170922 522300
rect 378042 522288 378048 522300
rect 170916 522260 378048 522288
rect 170916 522248 170922 522260
rect 378042 522248 378048 522260
rect 378100 522248 378106 522300
rect 380894 522248 380900 522300
rect 380952 522288 380958 522300
rect 380952 522260 509234 522288
rect 380952 522248 380958 522260
rect 44082 522180 44088 522232
rect 44140 522220 44146 522232
rect 68370 522220 68376 522232
rect 44140 522192 68376 522220
rect 44140 522180 44146 522192
rect 68370 522180 68376 522192
rect 68428 522180 68434 522232
rect 253198 522180 253204 522232
rect 253256 522220 253262 522232
rect 381170 522220 381176 522232
rect 253256 522192 381176 522220
rect 253256 522180 253262 522192
rect 381170 522180 381176 522192
rect 381228 522180 381234 522232
rect 45278 522112 45284 522164
rect 45336 522152 45342 522164
rect 77478 522152 77484 522164
rect 45336 522124 77484 522152
rect 45336 522112 45342 522124
rect 77478 522112 77484 522124
rect 77536 522112 77542 522164
rect 331950 522112 331956 522164
rect 332008 522152 332014 522164
rect 451918 522152 451924 522164
rect 332008 522124 451924 522152
rect 332008 522112 332014 522124
rect 451918 522112 451924 522124
rect 451976 522112 451982 522164
rect 45094 522044 45100 522096
rect 45152 522084 45158 522096
rect 78490 522084 78496 522096
rect 45152 522056 78496 522084
rect 45152 522044 45158 522056
rect 78490 522044 78496 522056
rect 78548 522044 78554 522096
rect 369118 522044 369124 522096
rect 369176 522084 369182 522096
rect 375558 522084 375564 522096
rect 369176 522056 375564 522084
rect 369176 522044 369182 522056
rect 375558 522044 375564 522056
rect 375616 522044 375622 522096
rect 471054 522084 471060 522096
rect 383626 522056 471060 522084
rect 107838 522016 107844 522028
rect 60936 521988 107844 522016
rect 60936 521960 60964 521988
rect 107838 521976 107844 521988
rect 107896 521976 107902 522028
rect 374086 521976 374092 522028
rect 374144 522016 374150 522028
rect 383626 522016 383654 522056
rect 471054 522044 471060 522056
rect 471112 522044 471118 522096
rect 374144 521988 383654 522016
rect 509206 522016 509234 522260
rect 517514 522248 517520 522300
rect 517572 522288 517578 522300
rect 538674 522288 538680 522300
rect 517572 522260 538680 522288
rect 517572 522248 517578 522260
rect 538674 522248 538680 522260
rect 538732 522248 538738 522300
rect 517514 522016 517520 522028
rect 509206 521988 517520 522016
rect 374144 521976 374150 521988
rect 517514 521976 517520 521988
rect 517572 521976 517578 522028
rect 60918 521908 60924 521960
rect 60976 521908 60982 521960
rect 125962 521948 125968 521960
rect 61028 521920 125968 521948
rect 60826 521840 60832 521892
rect 60884 521880 60890 521892
rect 61028 521880 61056 521920
rect 125962 521908 125968 521920
rect 126020 521908 126026 521960
rect 144822 521908 144828 521960
rect 144880 521948 144886 521960
rect 149238 521948 149244 521960
rect 144880 521920 149244 521948
rect 144880 521908 144886 521920
rect 149238 521908 149244 521920
rect 149296 521908 149302 521960
rect 60884 521852 61056 521880
rect 60884 521840 60890 521852
rect 61102 521840 61108 521892
rect 61160 521880 61166 521892
rect 131114 521880 131120 521892
rect 61160 521852 131120 521880
rect 61160 521840 61166 521852
rect 131114 521840 131120 521852
rect 131172 521840 131178 521892
rect 205174 521840 205180 521892
rect 205232 521880 205238 521892
rect 303614 521880 303620 521892
rect 205232 521852 303620 521880
rect 205232 521840 205238 521852
rect 303614 521840 303620 521852
rect 303672 521840 303678 521892
rect 497458 521840 497464 521892
rect 497516 521880 497522 521892
rect 500954 521880 500960 521892
rect 497516 521852 500960 521880
rect 497516 521840 497522 521852
rect 500954 521840 500960 521852
rect 501012 521840 501018 521892
rect 42610 521772 42616 521824
rect 42668 521812 42674 521824
rect 115934 521812 115940 521824
rect 42668 521784 115940 521812
rect 42668 521772 42674 521784
rect 115934 521772 115940 521784
rect 115992 521772 115998 521824
rect 160554 521772 160560 521824
rect 160612 521812 160618 521824
rect 269022 521812 269028 521824
rect 160612 521784 269028 521812
rect 160612 521772 160618 521784
rect 269022 521772 269028 521784
rect 269080 521772 269086 521824
rect 376662 521772 376668 521824
rect 376720 521812 376726 521824
rect 500586 521812 500592 521824
rect 376720 521784 500592 521812
rect 376720 521772 376726 521784
rect 500586 521772 500592 521784
rect 500644 521772 500650 521824
rect 43806 521704 43812 521756
rect 43864 521744 43870 521756
rect 129090 521744 129096 521756
rect 43864 521716 129096 521744
rect 43864 521704 43870 521716
rect 129090 521704 129096 521716
rect 129148 521704 129154 521756
rect 145466 521704 145472 521756
rect 145524 521744 145530 521756
rect 256694 521744 256700 521756
rect 145524 521716 256700 521744
rect 145524 521704 145530 521716
rect 256694 521704 256700 521716
rect 256752 521704 256758 521756
rect 377950 521704 377956 521756
rect 378008 521744 378014 521756
rect 508590 521744 508596 521756
rect 378008 521716 508596 521744
rect 378008 521704 378014 521716
rect 508590 521704 508596 521716
rect 508648 521704 508654 521756
rect 45186 521636 45192 521688
rect 45244 521676 45250 521688
rect 79410 521676 79416 521688
rect 45244 521648 79416 521676
rect 45244 521636 45250 521648
rect 79410 521636 79416 521648
rect 79468 521636 79474 521688
rect 81618 521636 81624 521688
rect 81676 521676 81682 521688
rect 313274 521676 313280 521688
rect 81676 521648 313280 521676
rect 81676 521636 81682 521648
rect 313274 521636 313280 521648
rect 313332 521636 313338 521688
rect 378778 521636 378784 521688
rect 378836 521676 378842 521688
rect 523218 521676 523224 521688
rect 378836 521648 523224 521676
rect 378836 521636 378842 521648
rect 523218 521636 523224 521648
rect 523276 521636 523282 521688
rect 50982 521568 50988 521620
rect 51040 521608 51046 521620
rect 51040 521580 58388 521608
rect 51040 521568 51046 521580
rect 58360 521472 58388 521580
rect 59354 521568 59360 521620
rect 59412 521608 59418 521620
rect 62850 521608 62856 521620
rect 59412 521580 62856 521608
rect 59412 521568 59418 521580
rect 62850 521568 62856 521580
rect 62908 521568 62914 521620
rect 167086 521568 167092 521620
rect 167144 521608 167150 521620
rect 382274 521608 382280 521620
rect 167144 521580 382280 521608
rect 167144 521568 167150 521580
rect 382274 521568 382280 521580
rect 382332 521568 382338 521620
rect 479518 521568 479524 521620
rect 479576 521608 479582 521620
rect 500126 521608 500132 521620
rect 479576 521580 500132 521608
rect 479576 521568 479582 521580
rect 500126 521568 500132 521580
rect 500184 521568 500190 521620
rect 510246 521568 510252 521620
rect 510304 521608 510310 521620
rect 513466 521608 513472 521620
rect 510304 521580 513472 521608
rect 510304 521568 510310 521580
rect 513466 521568 513472 521580
rect 513524 521568 513530 521620
rect 58434 521500 58440 521552
rect 58492 521540 58498 521552
rect 59446 521540 59452 521552
rect 58492 521512 59452 521540
rect 58492 521500 58498 521512
rect 59446 521500 59452 521512
rect 59504 521500 59510 521552
rect 59722 521500 59728 521552
rect 59780 521500 59786 521552
rect 168374 521500 168380 521552
rect 168432 521540 168438 521552
rect 382366 521540 382372 521552
rect 168432 521512 382372 521540
rect 168432 521500 168438 521512
rect 382366 521500 382372 521512
rect 382424 521500 382430 521552
rect 497550 521500 497556 521552
rect 497608 521540 497614 521552
rect 514754 521540 514760 521552
rect 497608 521512 514760 521540
rect 497608 521500 497614 521512
rect 514754 521500 514760 521512
rect 514812 521500 514818 521552
rect 59740 521472 59768 521500
rect 58360 521444 59768 521472
rect 60550 521432 60556 521484
rect 60608 521432 60614 521484
rect 166258 521432 166264 521484
rect 166316 521472 166322 521484
rect 338942 521472 338948 521484
rect 166316 521444 338948 521472
rect 166316 521432 166322 521444
rect 338942 521432 338948 521444
rect 339000 521432 339006 521484
rect 51534 521364 51540 521416
rect 51592 521404 51598 521416
rect 60568 521404 60596 521432
rect 51592 521376 60596 521404
rect 51592 521364 51598 521376
rect 166994 521364 167000 521416
rect 167052 521404 167058 521416
rect 191098 521404 191104 521416
rect 167052 521376 191104 521404
rect 167052 521364 167058 521376
rect 191098 521364 191104 521376
rect 191156 521364 191162 521416
rect 220722 521364 220728 521416
rect 220780 521404 220786 521416
rect 380986 521404 380992 521416
rect 220780 521376 380992 521404
rect 220780 521364 220786 521376
rect 380986 521364 380992 521376
rect 381044 521364 381050 521416
rect 231762 521296 231768 521348
rect 231820 521336 231826 521348
rect 312630 521336 312636 521348
rect 231820 521308 312636 521336
rect 231820 521296 231826 521308
rect 312630 521296 312636 521308
rect 312688 521296 312694 521348
rect 498746 521296 498752 521348
rect 498804 521336 498810 521348
rect 501230 521336 501236 521348
rect 498804 521308 501236 521336
rect 498804 521296 498810 521308
rect 501230 521296 501236 521308
rect 501288 521296 501294 521348
rect 43622 521228 43628 521280
rect 43680 521268 43686 521280
rect 73338 521268 73344 521280
rect 43680 521240 73344 521268
rect 43680 521228 43686 521240
rect 73338 521228 73344 521240
rect 73396 521228 73402 521280
rect 222102 521228 222108 521280
rect 222160 521268 222166 521280
rect 293310 521268 293316 521280
rect 222160 521240 293316 521268
rect 222160 521228 222166 521240
rect 293310 521228 293316 521240
rect 293368 521228 293374 521280
rect 499022 521228 499028 521280
rect 499080 521268 499086 521280
rect 501782 521268 501788 521280
rect 499080 521240 501788 521268
rect 499080 521228 499086 521240
rect 501782 521228 501788 521240
rect 501840 521228 501846 521280
rect 41138 521160 41144 521212
rect 41196 521200 41202 521212
rect 74442 521200 74448 521212
rect 41196 521172 74448 521200
rect 41196 521160 41202 521172
rect 74442 521160 74448 521172
rect 74500 521160 74506 521212
rect 498930 521160 498936 521212
rect 498988 521200 498994 521212
rect 501322 521200 501328 521212
rect 498988 521172 501328 521200
rect 498988 521160 498994 521172
rect 501322 521160 501328 521172
rect 501380 521160 501386 521212
rect 48774 521092 48780 521144
rect 48832 521132 48838 521144
rect 96614 521132 96620 521144
rect 48832 521104 96620 521132
rect 48832 521092 48838 521104
rect 96614 521092 96620 521104
rect 96672 521092 96678 521144
rect 471238 521092 471244 521144
rect 471296 521132 471302 521144
rect 518250 521132 518256 521144
rect 471296 521104 518256 521132
rect 471296 521092 471302 521104
rect 518250 521092 518256 521104
rect 518308 521092 518314 521144
rect 59630 521024 59636 521076
rect 59688 521064 59694 521076
rect 61838 521064 61844 521076
rect 59688 521036 61844 521064
rect 59688 521024 59694 521036
rect 61838 521024 61844 521036
rect 61896 521024 61902 521076
rect 146478 521024 146484 521076
rect 146536 521064 146542 521076
rect 285674 521064 285680 521076
rect 146536 521036 285680 521064
rect 146536 521024 146542 521036
rect 285674 521024 285680 521036
rect 285732 521024 285738 521076
rect 471422 521024 471428 521076
rect 471480 521064 471486 521076
rect 530302 521064 530308 521076
rect 471480 521036 530308 521064
rect 471480 521024 471486 521036
rect 530302 521024 530308 521036
rect 530360 521024 530366 521076
rect 53742 520956 53748 521008
rect 53800 520996 53806 521008
rect 59262 520996 59268 521008
rect 53800 520968 59268 520996
rect 53800 520956 53806 520968
rect 59262 520956 59268 520968
rect 59320 520956 59326 521008
rect 71866 520956 71872 521008
rect 71924 520996 71930 521008
rect 133138 520996 133144 521008
rect 71924 520968 133144 520996
rect 71924 520956 71930 520968
rect 133138 520956 133144 520968
rect 133196 520956 133202 521008
rect 254762 520956 254768 521008
rect 254820 520996 254826 521008
rect 524874 520996 524880 521008
rect 254820 520968 524880 520996
rect 254820 520956 254826 520968
rect 524874 520956 524880 520968
rect 524932 520956 524938 521008
rect 34422 520888 34428 520940
rect 34480 520928 34486 520940
rect 52454 520928 52460 520940
rect 34480 520900 52460 520928
rect 34480 520888 34486 520900
rect 52454 520888 52460 520900
rect 52512 520888 52518 520940
rect 59814 520888 59820 520940
rect 59872 520928 59878 520940
rect 62758 520928 62764 520940
rect 59872 520900 62764 520928
rect 59872 520888 59878 520900
rect 62758 520888 62764 520900
rect 62816 520888 62822 520940
rect 71958 520888 71964 520940
rect 72016 520928 72022 520940
rect 141142 520928 141148 520940
rect 72016 520900 141148 520928
rect 72016 520888 72022 520900
rect 141142 520888 141148 520900
rect 141200 520888 141206 520940
rect 193950 520888 193956 520940
rect 194008 520928 194014 520940
rect 496722 520928 496728 520940
rect 194008 520900 496728 520928
rect 194008 520888 194014 520900
rect 496722 520888 496728 520900
rect 496780 520888 496786 520940
rect 499206 520888 499212 520940
rect 499264 520928 499270 520940
rect 500770 520928 500776 520940
rect 499264 520900 500776 520928
rect 499264 520888 499270 520900
rect 500770 520888 500776 520900
rect 500828 520888 500834 520940
rect 505922 520888 505928 520940
rect 505980 520928 505986 520940
rect 520366 520928 520372 520940
rect 505980 520900 520372 520928
rect 505980 520888 505986 520900
rect 520366 520888 520372 520900
rect 520424 520888 520430 520940
rect 42242 520820 42248 520872
rect 42300 520860 42306 520872
rect 71314 520860 71320 520872
rect 42300 520832 71320 520860
rect 42300 520820 42306 520832
rect 71314 520820 71320 520832
rect 71372 520820 71378 520872
rect 498838 520820 498844 520872
rect 498896 520860 498902 520872
rect 500678 520860 500684 520872
rect 498896 520832 500684 520860
rect 498896 520820 498902 520832
rect 500678 520820 500684 520832
rect 500736 520820 500742 520872
rect 45370 520752 45376 520804
rect 45428 520792 45434 520804
rect 76466 520792 76472 520804
rect 45428 520764 76472 520792
rect 45428 520752 45434 520764
rect 76466 520752 76472 520764
rect 76524 520752 76530 520804
rect 504266 520792 504272 520804
rect 495406 520764 504272 520792
rect 40862 520684 40868 520736
rect 40920 520724 40926 520736
rect 75362 520724 75368 520736
rect 40920 520696 75368 520724
rect 40920 520684 40926 520696
rect 75362 520684 75368 520696
rect 75420 520684 75426 520736
rect 59262 520616 59268 520668
rect 59320 520656 59326 520668
rect 59722 520656 59728 520668
rect 59320 520628 59728 520656
rect 59320 520616 59326 520628
rect 59722 520616 59728 520628
rect 59780 520616 59786 520668
rect 59998 520616 60004 520668
rect 60056 520656 60062 520668
rect 106826 520656 106832 520668
rect 60056 520628 106832 520656
rect 60056 520616 60062 520628
rect 106826 520616 106832 520628
rect 106884 520616 106890 520668
rect 291838 520616 291844 520668
rect 291896 520656 291902 520668
rect 495406 520656 495434 520764
rect 504266 520752 504272 520764
rect 504324 520752 504330 520804
rect 498102 520684 498108 520736
rect 498160 520724 498166 520736
rect 515030 520724 515036 520736
rect 498160 520696 515036 520724
rect 498160 520684 498166 520696
rect 515030 520684 515036 520696
rect 515088 520684 515094 520736
rect 291896 520628 495434 520656
rect 496096 520628 504404 520656
rect 291896 520616 291902 520628
rect 59446 520548 59452 520600
rect 59504 520588 59510 520600
rect 119890 520588 119896 520600
rect 59504 520560 119896 520588
rect 59504 520548 59510 520560
rect 119890 520548 119896 520560
rect 119948 520548 119954 520600
rect 288342 520548 288348 520600
rect 288400 520588 288406 520600
rect 496096 520588 496124 520628
rect 504376 520600 504404 520628
rect 288400 520560 496124 520588
rect 288400 520548 288406 520560
rect 496170 520548 496176 520600
rect 496228 520588 496234 520600
rect 500402 520588 500408 520600
rect 496228 520560 500408 520588
rect 496228 520548 496234 520560
rect 500402 520548 500408 520560
rect 500460 520548 500466 520600
rect 504358 520548 504364 520600
rect 504416 520548 504422 520600
rect 52362 520480 52368 520532
rect 52420 520520 52426 520532
rect 113910 520520 113916 520532
rect 52420 520492 113916 520520
rect 52420 520480 52426 520492
rect 113910 520480 113916 520492
rect 113968 520480 113974 520532
rect 207198 520480 207204 520532
rect 207256 520520 207262 520532
rect 521838 520520 521844 520532
rect 207256 520492 521844 520520
rect 207256 520480 207262 520492
rect 521838 520480 521844 520492
rect 521896 520480 521902 520532
rect 57974 520412 57980 520464
rect 58032 520452 58038 520464
rect 60182 520452 60188 520464
rect 58032 520424 60188 520452
rect 58032 520412 58038 520424
rect 60182 520412 60188 520424
rect 60240 520412 60246 520464
rect 61654 520452 61660 520464
rect 60384 520424 61660 520452
rect 59722 520344 59728 520396
rect 59780 520384 59786 520396
rect 60384 520384 60412 520424
rect 61654 520412 61660 520424
rect 61712 520412 61718 520464
rect 62114 520412 62120 520464
rect 62172 520452 62178 520464
rect 127986 520452 127992 520464
rect 62172 520424 127992 520452
rect 62172 520412 62178 520424
rect 127986 520412 127992 520424
rect 128044 520412 128050 520464
rect 164694 520412 164700 520464
rect 164752 520452 164758 520464
rect 498010 520452 498016 520464
rect 164752 520424 498016 520452
rect 164752 520412 164758 520424
rect 498010 520412 498016 520424
rect 498068 520412 498074 520464
rect 498102 520412 498108 520464
rect 498160 520452 498166 520464
rect 537202 520452 537208 520464
rect 498160 520424 537208 520452
rect 498160 520412 498166 520424
rect 537202 520412 537208 520424
rect 537260 520412 537266 520464
rect 59780 520356 60412 520384
rect 59780 520344 59786 520356
rect 60550 520344 60556 520396
rect 60608 520384 60614 520396
rect 134058 520384 134064 520396
rect 60608 520356 134064 520384
rect 60608 520344 60614 520356
rect 134058 520344 134064 520356
rect 134116 520344 134122 520396
rect 188982 520344 188988 520396
rect 189040 520384 189046 520396
rect 545298 520384 545304 520396
rect 189040 520356 545304 520384
rect 189040 520344 189046 520356
rect 545298 520344 545304 520356
rect 545356 520344 545362 520396
rect 43530 520276 43536 520328
rect 43588 520316 43594 520328
rect 72326 520316 72332 520328
rect 43588 520288 72332 520316
rect 43588 520276 43594 520288
rect 72326 520276 72332 520288
rect 72384 520276 72390 520328
rect 86678 520276 86684 520328
rect 86736 520316 86742 520328
rect 516410 520316 516416 520328
rect 86736 520288 516416 520316
rect 86736 520276 86742 520288
rect 516410 520276 516416 520288
rect 516468 520276 516474 520328
rect 56134 520208 56140 520260
rect 56192 520248 56198 520260
rect 61102 520248 61108 520260
rect 56192 520220 61108 520248
rect 56192 520208 56198 520220
rect 61102 520208 61108 520220
rect 61160 520208 61166 520260
rect 61194 520208 61200 520260
rect 61252 520248 61258 520260
rect 61838 520248 61844 520260
rect 61252 520220 61844 520248
rect 61252 520208 61258 520220
rect 61838 520208 61844 520220
rect 61896 520208 61902 520260
rect 498194 520208 498200 520260
rect 498252 520248 498258 520260
rect 498252 520220 500632 520248
rect 498252 520208 498258 520220
rect 53282 520140 53288 520192
rect 53340 520180 53346 520192
rect 59630 520180 59636 520192
rect 53340 520152 59636 520180
rect 53340 520140 53346 520152
rect 59630 520140 59636 520152
rect 59688 520140 59694 520192
rect 59814 520140 59820 520192
rect 59872 520140 59878 520192
rect 60458 520140 60464 520192
rect 60516 520180 60522 520192
rect 62022 520180 62028 520192
rect 60516 520152 62028 520180
rect 60516 520140 60522 520152
rect 62022 520140 62028 520152
rect 62080 520140 62086 520192
rect 499298 520140 499304 520192
rect 499356 520180 499362 520192
rect 500604 520180 500632 520220
rect 500678 520208 500684 520260
rect 500736 520248 500742 520260
rect 507946 520248 507952 520260
rect 500736 520220 507952 520248
rect 500736 520208 500742 520220
rect 507946 520208 507952 520220
rect 508004 520208 508010 520260
rect 506014 520180 506020 520192
rect 499356 520152 500540 520180
rect 500604 520152 506020 520180
rect 499356 520140 499362 520152
rect 52730 520072 52736 520124
rect 52788 520112 52794 520124
rect 59832 520112 59860 520140
rect 52788 520084 59860 520112
rect 52788 520072 52794 520084
rect 60182 520072 60188 520124
rect 60240 520112 60246 520124
rect 61746 520112 61752 520124
rect 60240 520084 61752 520112
rect 60240 520072 60246 520084
rect 61746 520072 61752 520084
rect 61804 520072 61810 520124
rect 498010 520072 498016 520124
rect 498068 520112 498074 520124
rect 500512 520112 500540 520152
rect 506014 520140 506020 520152
rect 506072 520140 506078 520192
rect 505922 520112 505928 520124
rect 498068 520084 499574 520112
rect 500512 520084 505928 520112
rect 498068 520072 498074 520084
rect 56502 520004 56508 520056
rect 56560 520044 56566 520056
rect 60642 520044 60648 520056
rect 56560 520016 60648 520044
rect 56560 520004 56566 520016
rect 60642 520004 60648 520016
rect 60700 520004 60706 520056
rect 499546 520044 499574 520084
rect 505922 520072 505928 520084
rect 505980 520072 505986 520124
rect 509234 520112 509240 520124
rect 509206 520072 509240 520112
rect 509292 520072 509298 520124
rect 509206 520044 509234 520072
rect 499546 520016 509234 520044
rect 502242 519868 502248 519920
rect 502300 519908 502306 519920
rect 510614 519908 510620 519920
rect 502300 519880 510620 519908
rect 502300 519868 502306 519880
rect 510614 519868 510620 519880
rect 510672 519868 510678 519920
rect 501230 519800 501236 519852
rect 501288 519800 501294 519852
rect 501322 519800 501328 519852
rect 501380 519840 501386 519852
rect 501380 519812 505094 519840
rect 501380 519800 501386 519812
rect 501248 519772 501276 519800
rect 502242 519772 502248 519784
rect 501248 519744 502248 519772
rect 502242 519732 502248 519744
rect 502300 519732 502306 519784
rect 52362 519664 52368 519716
rect 52420 519704 52426 519716
rect 52420 519676 60872 519704
rect 52420 519664 52426 519676
rect 43714 519596 43720 519648
rect 43772 519636 43778 519648
rect 52546 519636 52552 519648
rect 43772 519608 52552 519636
rect 43772 519596 43778 519608
rect 52546 519596 52552 519608
rect 52604 519596 52610 519648
rect 28902 519528 28908 519580
rect 28960 519568 28966 519580
rect 59998 519568 60004 519580
rect 28960 519540 60004 519568
rect 28960 519528 28966 519540
rect 59998 519528 60004 519540
rect 60056 519528 60062 519580
rect 60844 519512 60872 519676
rect 501322 519664 501328 519716
rect 501380 519704 501386 519716
rect 502150 519704 502156 519716
rect 501380 519676 502156 519704
rect 501380 519664 501386 519676
rect 502150 519664 502156 519676
rect 502208 519664 502214 519716
rect 501874 519596 501880 519648
rect 501932 519636 501938 519648
rect 503714 519636 503720 519648
rect 501932 519608 503720 519636
rect 501932 519596 501938 519608
rect 503714 519596 503720 519608
rect 503772 519596 503778 519648
rect 505066 519636 505094 519812
rect 509510 519636 509516 519648
rect 505066 519608 509516 519636
rect 509510 519596 509516 519608
rect 509568 519596 509574 519648
rect 60918 519528 60924 519580
rect 60976 519528 60982 519580
rect 501322 519528 501328 519580
rect 501380 519568 501386 519580
rect 501690 519568 501696 519580
rect 501380 519540 501696 519568
rect 501380 519528 501386 519540
rect 501690 519528 501696 519540
rect 501748 519528 501754 519580
rect 60826 519460 60832 519512
rect 60884 519460 60890 519512
rect 60642 519052 60648 519104
rect 60700 519092 60706 519104
rect 60936 519092 60964 519528
rect 60700 519064 60964 519092
rect 60700 519052 60706 519064
rect 58710 518984 58716 519036
rect 58768 519024 58774 519036
rect 60918 519024 60924 519036
rect 58768 518996 60924 519024
rect 58768 518984 58774 518996
rect 60918 518984 60924 518996
rect 60976 518984 60982 519036
rect 49510 518916 49516 518968
rect 49568 518956 49574 518968
rect 55858 518956 55864 518968
rect 49568 518928 55864 518956
rect 49568 518916 49574 518928
rect 55858 518916 55864 518928
rect 55916 518916 55922 518968
rect 57698 516128 57704 516180
rect 57756 516168 57762 516180
rect 59354 516168 59360 516180
rect 57756 516140 59360 516168
rect 57756 516128 57762 516140
rect 59354 516128 59360 516140
rect 59412 516128 59418 516180
rect 53742 514836 53748 514888
rect 53800 514876 53806 514888
rect 54570 514876 54576 514888
rect 53800 514848 54576 514876
rect 53800 514836 53806 514848
rect 54570 514836 54576 514848
rect 54628 514836 54634 514888
rect 53466 514768 53472 514820
rect 53524 514808 53530 514820
rect 54478 514808 54484 514820
rect 53524 514780 54484 514808
rect 53524 514768 53530 514780
rect 54478 514768 54484 514780
rect 54536 514768 54542 514820
rect 53650 514700 53656 514752
rect 53708 514740 53714 514752
rect 55858 514740 55864 514752
rect 53708 514712 55864 514740
rect 53708 514700 53714 514712
rect 55858 514700 55864 514712
rect 55916 514700 55922 514752
rect 53282 514020 53288 514072
rect 53340 514060 53346 514072
rect 53650 514060 53656 514072
rect 53340 514032 53656 514060
rect 53340 514020 53346 514032
rect 53650 514020 53656 514032
rect 53708 514020 53714 514072
rect 57974 513272 57980 513324
rect 58032 513312 58038 513324
rect 58526 513312 58532 513324
rect 58032 513284 58532 513312
rect 58032 513272 58038 513284
rect 58526 513272 58532 513284
rect 58584 513272 58590 513324
rect 500310 513272 500316 513324
rect 500368 513312 500374 513324
rect 500954 513312 500960 513324
rect 500368 513284 500960 513312
rect 500368 513272 500374 513284
rect 500954 513272 500960 513284
rect 501012 513272 501018 513324
rect 500494 512592 500500 512644
rect 500552 512632 500558 512644
rect 509326 512632 509332 512644
rect 500552 512604 509332 512632
rect 500552 512592 500558 512604
rect 509326 512592 509332 512604
rect 509384 512592 509390 512644
rect 57882 511912 57888 511964
rect 57940 511952 57946 511964
rect 59446 511952 59452 511964
rect 57940 511924 59452 511952
rect 57940 511912 57946 511924
rect 59446 511912 59452 511924
rect 59504 511912 59510 511964
rect 510522 511912 510528 511964
rect 510580 511952 510586 511964
rect 580166 511952 580172 511964
rect 510580 511924 580172 511952
rect 510580 511912 510586 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 53282 511232 53288 511284
rect 53340 511272 53346 511284
rect 58618 511272 58624 511284
rect 53340 511244 58624 511272
rect 53340 511232 53346 511244
rect 58618 511232 58624 511244
rect 58676 511232 58682 511284
rect 500402 511232 500408 511284
rect 500460 511272 500466 511284
rect 510522 511272 510528 511284
rect 500460 511244 510528 511272
rect 500460 511232 500466 511244
rect 510522 511232 510528 511244
rect 510580 511232 510586 511284
rect 55030 510620 55036 510672
rect 55088 510660 55094 510672
rect 56594 510660 56600 510672
rect 55088 510632 56600 510660
rect 55088 510620 55094 510632
rect 56594 510620 56600 510632
rect 56652 510620 56658 510672
rect 511442 510008 511448 510060
rect 511500 510048 511506 510060
rect 511626 510048 511632 510060
rect 511500 510020 511632 510048
rect 511500 510008 511506 510020
rect 511626 510008 511632 510020
rect 511684 510008 511690 510060
rect 53742 509872 53748 509924
rect 53800 509912 53806 509924
rect 57974 509912 57980 509924
rect 53800 509884 57980 509912
rect 53800 509872 53806 509884
rect 57974 509872 57980 509884
rect 58032 509872 58038 509924
rect 49510 507832 49516 507884
rect 49568 507872 49574 507884
rect 57146 507872 57152 507884
rect 49568 507844 57152 507872
rect 49568 507832 49574 507844
rect 57146 507832 57152 507844
rect 57204 507832 57210 507884
rect 57790 507832 57796 507884
rect 57848 507872 57854 507884
rect 58710 507872 58716 507884
rect 57848 507844 58716 507872
rect 57848 507832 57854 507844
rect 58710 507832 58716 507844
rect 58768 507832 58774 507884
rect 55858 505112 55864 505164
rect 55916 505152 55922 505164
rect 59354 505152 59360 505164
rect 55916 505124 59360 505152
rect 55916 505112 55922 505124
rect 59354 505112 59360 505124
rect 59412 505112 59418 505164
rect 58526 504364 58532 504416
rect 58584 504404 58590 504416
rect 60182 504404 60188 504416
rect 58584 504376 60188 504404
rect 58584 504364 58590 504376
rect 60182 504364 60188 504376
rect 60240 504364 60246 504416
rect 55122 503616 55128 503668
rect 55180 503656 55186 503668
rect 56594 503656 56600 503668
rect 55180 503628 56600 503656
rect 55180 503616 55186 503628
rect 56594 503616 56600 503628
rect 56652 503616 56658 503668
rect 58434 503616 58440 503668
rect 58492 503656 58498 503668
rect 59814 503656 59820 503668
rect 58492 503628 59820 503656
rect 58492 503616 58498 503628
rect 59814 503616 59820 503628
rect 59872 503616 59878 503668
rect 52822 503072 52828 503124
rect 52880 503112 52886 503124
rect 58618 503112 58624 503124
rect 52880 503084 58624 503112
rect 52880 503072 52886 503084
rect 58618 503072 58624 503084
rect 58676 503072 58682 503124
rect 53650 501576 53656 501628
rect 53708 501616 53714 501628
rect 60090 501616 60096 501628
rect 53708 501588 60096 501616
rect 53708 501576 53714 501588
rect 60090 501576 60096 501588
rect 60148 501576 60154 501628
rect 57698 500896 57704 500948
rect 57756 500936 57762 500948
rect 58066 500936 58072 500948
rect 57756 500908 58072 500936
rect 57756 500896 57762 500908
rect 58066 500896 58072 500908
rect 58124 500896 58130 500948
rect 59814 500148 59820 500200
rect 59872 500188 59878 500200
rect 60182 500188 60188 500200
rect 59872 500160 60188 500188
rect 59872 500148 59878 500160
rect 60182 500148 60188 500160
rect 60240 500148 60246 500200
rect 55122 499536 55128 499588
rect 55180 499576 55186 499588
rect 57238 499576 57244 499588
rect 55180 499548 57244 499576
rect 55180 499536 55186 499548
rect 57238 499536 57244 499548
rect 57296 499536 57302 499588
rect 57606 498992 57612 499044
rect 57664 498992 57670 499044
rect 57624 498840 57652 498992
rect 57606 498788 57612 498840
rect 57664 498788 57670 498840
rect 27522 497428 27528 497480
rect 27580 497468 27586 497480
rect 43346 497468 43352 497480
rect 27580 497440 43352 497468
rect 27580 497428 27586 497440
rect 43346 497428 43352 497440
rect 43404 497428 43410 497480
rect 28902 496748 28908 496800
rect 28960 496788 28966 496800
rect 31846 496788 31852 496800
rect 28960 496760 31852 496788
rect 28960 496748 28966 496760
rect 31846 496748 31852 496760
rect 31904 496748 31910 496800
rect 57698 496272 57704 496324
rect 57756 496312 57762 496324
rect 60274 496312 60280 496324
rect 57756 496284 60280 496312
rect 57756 496272 57762 496284
rect 60274 496272 60280 496284
rect 60332 496272 60338 496324
rect 34422 495456 34428 495508
rect 34480 495496 34486 495508
rect 35066 495496 35072 495508
rect 34480 495468 35072 495496
rect 34480 495456 34486 495468
rect 35066 495456 35072 495468
rect 35124 495456 35130 495508
rect 57146 494708 57152 494760
rect 57204 494748 57210 494760
rect 58710 494748 58716 494760
rect 57204 494720 58716 494748
rect 57204 494708 57210 494720
rect 58710 494708 58716 494720
rect 58768 494708 58774 494760
rect 31846 493960 31852 494012
rect 31904 494000 31910 494012
rect 38102 494000 38108 494012
rect 31904 493972 38108 494000
rect 31904 493960 31910 493972
rect 38102 493960 38108 493972
rect 38160 493960 38166 494012
rect 46474 493280 46480 493332
rect 46532 493320 46538 493332
rect 57974 493320 57980 493332
rect 46532 493292 57980 493320
rect 46532 493280 46538 493292
rect 57974 493280 57980 493292
rect 58032 493280 58038 493332
rect 57146 491580 57152 491632
rect 57204 491620 57210 491632
rect 57514 491620 57520 491632
rect 57204 491592 57520 491620
rect 57204 491580 57210 491592
rect 57514 491580 57520 491592
rect 57572 491580 57578 491632
rect 57790 488588 57796 488640
rect 57848 488628 57854 488640
rect 58802 488628 58808 488640
rect 57848 488600 58808 488628
rect 57848 488588 57854 488600
rect 58802 488588 58808 488600
rect 58860 488588 58866 488640
rect 57698 488520 57704 488572
rect 57756 488560 57762 488572
rect 58066 488560 58072 488572
rect 57756 488532 58072 488560
rect 57756 488520 57762 488532
rect 58066 488520 58072 488532
rect 58124 488520 58130 488572
rect 503622 488452 503628 488504
rect 503680 488492 503686 488504
rect 511166 488492 511172 488504
rect 503680 488464 511172 488492
rect 503680 488452 503686 488464
rect 511166 488452 511172 488464
rect 511224 488452 511230 488504
rect 500034 486072 500040 486124
rect 500092 486112 500098 486124
rect 500494 486112 500500 486124
rect 500092 486084 500500 486112
rect 500092 486072 500098 486084
rect 500494 486072 500500 486084
rect 500552 486072 500558 486124
rect 502334 485392 502340 485444
rect 502392 485432 502398 485444
rect 502392 485404 502472 485432
rect 502392 485392 502398 485404
rect 502444 485240 502472 485404
rect 502426 485188 502432 485240
rect 502484 485188 502490 485240
rect 502978 485052 502984 485104
rect 503036 485092 503042 485104
rect 541434 485092 541440 485104
rect 503036 485064 541440 485092
rect 503036 485052 503042 485064
rect 541434 485052 541440 485064
rect 541492 485052 541498 485104
rect 501598 483624 501604 483676
rect 501656 483664 501662 483676
rect 517698 483664 517704 483676
rect 501656 483636 517704 483664
rect 501656 483624 501662 483636
rect 517698 483624 517704 483636
rect 517756 483624 517762 483676
rect 503530 482944 503536 482996
rect 503588 482984 503594 482996
rect 505830 482984 505836 482996
rect 503588 482956 505836 482984
rect 503588 482944 503594 482956
rect 505830 482944 505836 482956
rect 505888 482944 505894 482996
rect 508590 482400 508596 482452
rect 508648 482440 508654 482452
rect 517698 482440 517704 482452
rect 508648 482412 517704 482440
rect 508648 482400 508654 482412
rect 517698 482400 517704 482412
rect 517756 482400 517762 482452
rect 503438 482332 503444 482384
rect 503496 482372 503502 482384
rect 515582 482372 515588 482384
rect 503496 482344 515588 482372
rect 503496 482332 503502 482344
rect 515582 482332 515588 482344
rect 515640 482332 515646 482384
rect 503162 482264 503168 482316
rect 503220 482304 503226 482316
rect 516870 482304 516876 482316
rect 503220 482276 516876 482304
rect 503220 482264 503226 482276
rect 516870 482264 516876 482276
rect 516928 482264 516934 482316
rect 503070 481720 503076 481772
rect 503128 481760 503134 481772
rect 509878 481760 509884 481772
rect 503128 481732 509884 481760
rect 503128 481720 503134 481732
rect 509878 481720 509884 481732
rect 509936 481720 509942 481772
rect 502978 480836 502984 480888
rect 503036 480876 503042 480888
rect 503254 480876 503260 480888
rect 503036 480848 503260 480876
rect 503036 480836 503042 480848
rect 503254 480836 503260 480848
rect 503312 480836 503318 480888
rect 26878 479476 26884 479528
rect 26936 479516 26942 479528
rect 37918 479516 37924 479528
rect 26936 479488 37924 479516
rect 26936 479476 26942 479488
rect 37918 479476 37924 479488
rect 37976 479476 37982 479528
rect 503254 478864 503260 478916
rect 503312 478904 503318 478916
rect 511258 478904 511264 478916
rect 503312 478876 511264 478904
rect 503312 478864 503318 478876
rect 511258 478864 511264 478876
rect 511316 478864 511322 478916
rect 38102 478116 38108 478168
rect 38160 478156 38166 478168
rect 51810 478156 51816 478168
rect 38160 478128 51816 478156
rect 38160 478116 38166 478128
rect 51810 478116 51816 478128
rect 51868 478116 51874 478168
rect 503530 478116 503536 478168
rect 503588 478156 503594 478168
rect 538674 478156 538680 478168
rect 503588 478128 538680 478156
rect 503588 478116 503594 478128
rect 538674 478116 538680 478128
rect 538732 478116 538738 478168
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 11698 474756 11704 474768
rect 3476 474728 11704 474756
rect 3476 474716 3482 474728
rect 11698 474716 11704 474728
rect 11756 474716 11762 474768
rect 502886 470500 502892 470552
rect 502944 470540 502950 470552
rect 536282 470540 536288 470552
rect 502944 470512 536288 470540
rect 502944 470500 502950 470512
rect 536282 470500 536288 470512
rect 536340 470500 536346 470552
rect 502886 469140 502892 469192
rect 502944 469180 502950 469192
rect 534902 469180 534908 469192
rect 502944 469152 534908 469180
rect 502944 469140 502950 469152
rect 534902 469140 534908 469152
rect 534960 469140 534966 469192
rect 502794 469072 502800 469124
rect 502852 469112 502858 469124
rect 522390 469112 522396 469124
rect 502852 469084 522396 469112
rect 502852 469072 502858 469084
rect 522390 469072 522396 469084
rect 522448 469072 522454 469124
rect 502702 467780 502708 467832
rect 502760 467820 502766 467832
rect 534718 467820 534724 467832
rect 502760 467792 534724 467820
rect 502760 467780 502766 467792
rect 534718 467780 534724 467792
rect 534776 467780 534782 467832
rect 502794 467712 502800 467764
rect 502852 467752 502858 467764
rect 530670 467752 530676 467764
rect 502852 467724 530676 467752
rect 502852 467712 502858 467724
rect 530670 467712 530676 467724
rect 530728 467712 530734 467764
rect 502886 467644 502892 467696
rect 502944 467684 502950 467696
rect 527910 467684 527916 467696
rect 502944 467656 527916 467684
rect 502944 467644 502950 467656
rect 527910 467644 527916 467656
rect 527968 467644 527974 467696
rect 35066 467100 35072 467152
rect 35124 467140 35130 467152
rect 51074 467140 51080 467152
rect 35124 467112 51080 467140
rect 35124 467100 35130 467112
rect 51074 467100 51080 467112
rect 51132 467100 51138 467152
rect 502702 466352 502708 466404
rect 502760 466392 502766 466404
rect 534626 466392 534632 466404
rect 502760 466364 534632 466392
rect 502760 466352 502766 466364
rect 534626 466352 534632 466364
rect 534684 466352 534690 466404
rect 502610 466284 502616 466336
rect 502668 466324 502674 466336
rect 534534 466324 534540 466336
rect 502668 466296 534540 466324
rect 502668 466284 502674 466296
rect 534534 466284 534540 466296
rect 534592 466284 534598 466336
rect 502794 466216 502800 466268
rect 502852 466256 502858 466268
rect 533246 466256 533252 466268
rect 502852 466228 533252 466256
rect 502852 466216 502858 466228
rect 533246 466216 533252 466228
rect 533304 466216 533310 466268
rect 502886 466148 502892 466200
rect 502944 466188 502950 466200
rect 533338 466188 533344 466200
rect 502944 466160 533344 466188
rect 502944 466148 502950 466160
rect 533338 466148 533344 466160
rect 533396 466148 533402 466200
rect 502886 464992 502892 465044
rect 502944 465032 502950 465044
rect 520918 465032 520924 465044
rect 502944 465004 520924 465032
rect 502944 464992 502950 465004
rect 520918 464992 520924 465004
rect 520976 464992 520982 465044
rect 502610 463632 502616 463684
rect 502668 463672 502674 463684
rect 527818 463672 527824 463684
rect 502668 463644 527824 463672
rect 502668 463632 502674 463644
rect 527818 463632 527824 463644
rect 527876 463632 527882 463684
rect 502702 463564 502708 463616
rect 502760 463604 502766 463616
rect 524966 463604 524972 463616
rect 502760 463576 524972 463604
rect 502760 463564 502766 463576
rect 524966 463564 524972 463576
rect 525024 463564 525030 463616
rect 502794 463496 502800 463548
rect 502852 463536 502858 463548
rect 518250 463536 518256 463548
rect 502852 463508 518256 463536
rect 502852 463496 502858 463508
rect 518250 463496 518256 463508
rect 518308 463496 518314 463548
rect 502886 463428 502892 463480
rect 502944 463468 502950 463480
rect 516778 463468 516784 463480
rect 502944 463440 516784 463468
rect 502944 463428 502950 463440
rect 516778 463428 516784 463440
rect 516836 463428 516842 463480
rect 51074 462272 51080 462324
rect 51132 462312 51138 462324
rect 54754 462312 54760 462324
rect 51132 462284 54760 462312
rect 51132 462272 51138 462284
rect 54754 462272 54760 462284
rect 54812 462272 54818 462324
rect 502518 462272 502524 462324
rect 502576 462312 502582 462324
rect 529290 462312 529296 462324
rect 502576 462284 529296 462312
rect 502576 462272 502582 462284
rect 529290 462272 529296 462284
rect 529348 462272 529354 462324
rect 502886 462204 502892 462256
rect 502944 462244 502950 462256
rect 529106 462244 529112 462256
rect 502944 462216 529112 462244
rect 502944 462204 502950 462216
rect 529106 462204 529112 462216
rect 529164 462204 529170 462256
rect 502610 462136 502616 462188
rect 502668 462176 502674 462188
rect 526530 462176 526536 462188
rect 502668 462148 526536 462176
rect 502668 462136 502674 462148
rect 526530 462136 526536 462148
rect 526588 462136 526594 462188
rect 502886 462068 502892 462120
rect 502944 462108 502950 462120
rect 525058 462108 525064 462120
rect 502944 462080 525064 462108
rect 502944 462068 502950 462080
rect 525058 462068 525064 462080
rect 525116 462068 525122 462120
rect 502794 462000 502800 462052
rect 502852 462040 502858 462052
rect 521010 462040 521016 462052
rect 502852 462012 521016 462040
rect 502852 462000 502858 462012
rect 521010 462000 521016 462012
rect 521068 462000 521074 462052
rect 502794 460844 502800 460896
rect 502852 460884 502858 460896
rect 544470 460884 544476 460896
rect 502852 460856 544476 460884
rect 502852 460844 502858 460856
rect 544470 460844 544476 460856
rect 544528 460844 544534 460896
rect 502886 460776 502892 460828
rect 502944 460816 502950 460828
rect 538582 460816 538588 460828
rect 502944 460788 538588 460816
rect 502944 460776 502950 460788
rect 538582 460776 538588 460788
rect 538640 460776 538646 460828
rect 502610 459484 502616 459536
rect 502668 459524 502674 459536
rect 531682 459524 531688 459536
rect 502668 459496 531688 459524
rect 502668 459484 502674 459496
rect 531682 459484 531688 459496
rect 531740 459484 531746 459536
rect 502886 459416 502892 459468
rect 502944 459456 502950 459468
rect 530486 459456 530492 459468
rect 502944 459428 530492 459456
rect 502944 459416 502950 459428
rect 530486 459416 530492 459428
rect 530544 459416 530550 459468
rect 502794 459348 502800 459400
rect 502852 459388 502858 459400
rect 529014 459388 529020 459400
rect 502852 459360 529020 459388
rect 502852 459348 502858 459360
rect 529014 459348 529020 459360
rect 529072 459348 529078 459400
rect 502702 459280 502708 459332
rect 502760 459320 502766 459332
rect 522206 459320 522212 459332
rect 502760 459292 522212 459320
rect 502760 459280 502766 459292
rect 522206 459280 522212 459292
rect 522264 459280 522270 459332
rect 502794 458124 502800 458176
rect 502852 458164 502858 458176
rect 534442 458164 534448 458176
rect 502852 458136 534448 458164
rect 502852 458124 502858 458136
rect 534442 458124 534448 458136
rect 534500 458124 534506 458176
rect 535730 458124 535736 458176
rect 535788 458164 535794 458176
rect 580166 458164 580172 458176
rect 535788 458136 580172 458164
rect 535788 458124 535794 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 502610 458056 502616 458108
rect 502668 458096 502674 458108
rect 537294 458096 537300 458108
rect 502668 458068 537300 458096
rect 502668 458056 502674 458068
rect 537294 458056 537300 458068
rect 537352 458056 537358 458108
rect 502702 457988 502708 458040
rect 502760 458028 502766 458040
rect 526346 458028 526352 458040
rect 502760 458000 526352 458028
rect 502760 457988 502766 458000
rect 526346 457988 526352 458000
rect 526404 457988 526410 458040
rect 502886 457920 502892 457972
rect 502944 457960 502950 457972
rect 518066 457960 518072 457972
rect 502944 457932 518072 457960
rect 502944 457920 502950 457932
rect 518066 457920 518072 457932
rect 518124 457920 518130 457972
rect 501690 457444 501696 457496
rect 501748 457484 501754 457496
rect 535730 457484 535736 457496
rect 501748 457456 535736 457484
rect 501748 457444 501754 457456
rect 535730 457444 535736 457456
rect 535788 457444 535794 457496
rect 502610 456696 502616 456748
rect 502668 456736 502674 456748
rect 536006 456736 536012 456748
rect 502668 456708 536012 456736
rect 502668 456696 502674 456708
rect 536006 456696 536012 456708
rect 536064 456696 536070 456748
rect 502886 456628 502892 456680
rect 502944 456668 502950 456680
rect 533154 456668 533160 456680
rect 502944 456640 533160 456668
rect 502944 456628 502950 456640
rect 533154 456628 533160 456640
rect 533212 456628 533218 456680
rect 502794 456560 502800 456612
rect 502852 456600 502858 456612
rect 530394 456600 530400 456612
rect 502852 456572 530400 456600
rect 502852 456560 502858 456572
rect 530394 456560 530400 456572
rect 530452 456560 530458 456612
rect 502886 456492 502892 456544
rect 502944 456532 502950 456544
rect 513926 456532 513932 456544
rect 502944 456504 513932 456532
rect 502944 456492 502950 456504
rect 513926 456492 513932 456504
rect 513984 456492 513990 456544
rect 502702 455336 502708 455388
rect 502760 455376 502766 455388
rect 531590 455376 531596 455388
rect 502760 455348 531596 455376
rect 502760 455336 502766 455348
rect 531590 455336 531596 455348
rect 531648 455336 531654 455388
rect 502518 455268 502524 455320
rect 502576 455308 502582 455320
rect 523310 455308 523316 455320
rect 502576 455280 523316 455308
rect 502576 455268 502582 455280
rect 523310 455268 523316 455280
rect 523368 455268 523374 455320
rect 502610 455200 502616 455252
rect 502668 455240 502674 455252
rect 522114 455240 522120 455252
rect 502668 455212 522120 455240
rect 502668 455200 502674 455212
rect 522114 455200 522120 455212
rect 522172 455200 522178 455252
rect 502794 455132 502800 455184
rect 502852 455172 502858 455184
rect 512178 455172 512184 455184
rect 502852 455144 512184 455172
rect 502852 455132 502858 455144
rect 512178 455132 512184 455144
rect 512236 455132 512242 455184
rect 502886 455064 502892 455116
rect 502944 455104 502950 455116
rect 509786 455104 509792 455116
rect 502944 455076 509792 455104
rect 502944 455064 502950 455076
rect 509786 455064 509792 455076
rect 509844 455064 509850 455116
rect 502886 453908 502892 453960
rect 502944 453948 502950 453960
rect 519630 453948 519636 453960
rect 502944 453920 519636 453948
rect 502944 453908 502950 453920
rect 519630 453908 519636 453920
rect 519688 453908 519694 453960
rect 502702 453840 502708 453892
rect 502760 453880 502766 453892
rect 514846 453880 514852 453892
rect 502760 453852 514852 453880
rect 502760 453840 502766 453852
rect 514846 453840 514852 453852
rect 514904 453840 514910 453892
rect 502794 453772 502800 453824
rect 502852 453812 502858 453824
rect 541618 453812 541624 453824
rect 502852 453784 541624 453812
rect 502852 453772 502858 453784
rect 541618 453772 541624 453784
rect 541676 453772 541682 453824
rect 502702 452548 502708 452600
rect 502760 452588 502766 452600
rect 515306 452588 515312 452600
rect 502760 452560 515312 452588
rect 502760 452548 502766 452560
rect 515306 452548 515312 452560
rect 515364 452548 515370 452600
rect 502610 452480 502616 452532
rect 502668 452520 502674 452532
rect 515122 452520 515128 452532
rect 502668 452492 515128 452520
rect 502668 452480 502674 452492
rect 515122 452480 515128 452492
rect 515180 452480 515186 452532
rect 502886 452412 502892 452464
rect 502944 452452 502950 452464
rect 514938 452452 514944 452464
rect 502944 452424 514944 452452
rect 502944 452412 502950 452424
rect 514938 452412 514944 452424
rect 514996 452412 515002 452464
rect 502794 452344 502800 452396
rect 502852 452384 502858 452396
rect 513834 452384 513840 452396
rect 502852 452356 513840 452384
rect 502852 452344 502858 452356
rect 513834 452344 513840 452356
rect 513892 452344 513898 452396
rect 502610 451188 502616 451240
rect 502668 451228 502674 451240
rect 526254 451228 526260 451240
rect 502668 451200 526260 451228
rect 502668 451188 502674 451200
rect 526254 451188 526260 451200
rect 526312 451188 526318 451240
rect 502702 451120 502708 451172
rect 502760 451160 502766 451172
rect 520734 451160 520740 451172
rect 502760 451132 520740 451160
rect 502760 451120 502766 451132
rect 520734 451120 520740 451132
rect 520792 451120 520798 451172
rect 503622 451052 503628 451104
rect 503680 451092 503686 451104
rect 513742 451092 513748 451104
rect 503680 451064 513748 451092
rect 503680 451052 503686 451064
rect 513742 451052 513748 451064
rect 513800 451052 513806 451104
rect 502886 450984 502892 451036
rect 502944 451024 502950 451036
rect 512822 451024 512828 451036
rect 502944 450996 512828 451024
rect 502944 450984 502950 450996
rect 512822 450984 512828 450996
rect 512880 450984 512886 451036
rect 503622 450916 503628 450968
rect 503680 450956 503686 450968
rect 507210 450956 507216 450968
rect 503680 450928 507216 450956
rect 503680 450916 503686 450928
rect 507210 450916 507216 450928
rect 507268 450916 507274 450968
rect 503622 449828 503628 449880
rect 503680 449868 503686 449880
rect 537110 449868 537116 449880
rect 503680 449840 537116 449868
rect 503680 449828 503686 449840
rect 537110 449828 537116 449840
rect 537168 449828 537174 449880
rect 502702 449760 502708 449812
rect 502760 449800 502766 449812
rect 537018 449800 537024 449812
rect 502760 449772 537024 449800
rect 502760 449760 502766 449772
rect 537018 449760 537024 449772
rect 537076 449760 537082 449812
rect 502794 449692 502800 449744
rect 502852 449732 502858 449744
rect 527634 449732 527640 449744
rect 502852 449704 527640 449732
rect 502852 449692 502858 449704
rect 527634 449692 527640 449704
rect 527692 449692 527698 449744
rect 502886 449624 502892 449676
rect 502944 449664 502950 449676
rect 524690 449664 524696 449676
rect 502944 449636 524696 449664
rect 502944 449624 502950 449636
rect 524690 449624 524696 449636
rect 524748 449624 524754 449676
rect 503622 449556 503628 449608
rect 503680 449596 503686 449608
rect 517974 449596 517980 449608
rect 503680 449568 517980 449596
rect 503680 449556 503686 449568
rect 517974 449556 517980 449568
rect 518032 449556 518038 449608
rect 502702 448468 502708 448520
rect 502760 448508 502766 448520
rect 540330 448508 540336 448520
rect 502760 448480 540336 448508
rect 502760 448468 502766 448480
rect 540330 448468 540336 448480
rect 540388 448468 540394 448520
rect 502610 448400 502616 448452
rect 502668 448440 502674 448452
rect 538490 448440 538496 448452
rect 502668 448412 538496 448440
rect 502668 448400 502674 448412
rect 538490 448400 538496 448412
rect 538548 448400 538554 448452
rect 503622 448332 503628 448384
rect 503680 448372 503686 448384
rect 516594 448372 516600 448384
rect 503680 448344 516600 448372
rect 503680 448332 503686 448344
rect 516594 448332 516600 448344
rect 516652 448332 516658 448384
rect 502886 448264 502892 448316
rect 502944 448304 502950 448316
rect 513558 448304 513564 448316
rect 502944 448276 513564 448304
rect 502944 448264 502950 448276
rect 513558 448264 513564 448276
rect 513616 448264 513622 448316
rect 503622 445680 503628 445732
rect 503680 445720 503686 445732
rect 538398 445720 538404 445732
rect 503680 445692 538404 445720
rect 503680 445680 503686 445692
rect 538398 445680 538404 445692
rect 538456 445680 538462 445732
rect 499850 444456 499856 444508
rect 499908 444496 499914 444508
rect 500126 444496 500132 444508
rect 499908 444468 500132 444496
rect 499908 444456 499914 444468
rect 500126 444456 500132 444468
rect 500184 444456 500190 444508
rect 503622 442892 503628 442944
rect 503680 442932 503686 442944
rect 545758 442932 545764 442944
rect 503680 442904 545764 442932
rect 503680 442892 503686 442904
rect 545758 442892 545764 442904
rect 545816 442892 545822 442944
rect 500218 441940 500224 441992
rect 500276 441980 500282 441992
rect 500862 441980 500868 441992
rect 500276 441952 500868 441980
rect 500276 441940 500282 441952
rect 500862 441940 500868 441952
rect 500920 441940 500926 441992
rect 503622 441124 503628 441176
rect 503680 441164 503686 441176
rect 508498 441164 508504 441176
rect 503680 441136 508504 441164
rect 503680 441124 503686 441136
rect 508498 441124 508504 441136
rect 508556 441124 508562 441176
rect 501874 440308 501880 440360
rect 501932 440348 501938 440360
rect 503530 440348 503536 440360
rect 501932 440320 503536 440348
rect 501932 440308 501938 440320
rect 503530 440308 503536 440320
rect 503588 440308 503594 440360
rect 501782 440240 501788 440292
rect 501840 440280 501846 440292
rect 502426 440280 502432 440292
rect 501840 440252 502432 440280
rect 501840 440240 501846 440252
rect 502426 440240 502432 440252
rect 502484 440240 502490 440292
rect 503622 440172 503628 440224
rect 503680 440212 503686 440224
rect 512914 440212 512920 440224
rect 503680 440184 512920 440212
rect 503680 440172 503686 440184
rect 512914 440172 512920 440184
rect 512972 440172 512978 440224
rect 503622 440036 503628 440088
rect 503680 440076 503686 440088
rect 510798 440076 510804 440088
rect 503680 440048 510804 440076
rect 503680 440036 503686 440048
rect 510798 440036 510804 440048
rect 510856 440036 510862 440088
rect 503530 438812 503536 438864
rect 503588 438852 503594 438864
rect 526162 438852 526168 438864
rect 503588 438824 526168 438852
rect 503588 438812 503594 438824
rect 526162 438812 526168 438824
rect 526220 438812 526226 438864
rect 503622 438744 503628 438796
rect 503680 438784 503686 438796
rect 524874 438784 524880 438796
rect 503680 438756 524880 438784
rect 503680 438744 503686 438756
rect 524874 438744 524880 438756
rect 524932 438744 524938 438796
rect 503622 437384 503628 437436
rect 503680 437424 503686 437436
rect 515214 437424 515220 437436
rect 503680 437396 515220 437424
rect 503680 437384 503686 437396
rect 515214 437384 515220 437396
rect 515272 437384 515278 437436
rect 503622 437044 503628 437096
rect 503680 437084 503686 437096
rect 511074 437084 511080 437096
rect 503680 437056 511080 437084
rect 503680 437044 503686 437056
rect 511074 437044 511080 437056
rect 511132 437044 511138 437096
rect 502886 436772 502892 436824
rect 502944 436812 502950 436824
rect 503438 436812 503444 436824
rect 502944 436784 503444 436812
rect 502944 436772 502950 436784
rect 503438 436772 503444 436784
rect 503496 436772 503502 436824
rect 503622 436024 503628 436076
rect 503680 436064 503686 436076
rect 541526 436064 541532 436076
rect 503680 436036 541532 436064
rect 503680 436024 503686 436036
rect 541526 436024 541532 436036
rect 541584 436024 541590 436076
rect 503438 435956 503444 436008
rect 503496 435996 503502 436008
rect 506934 435996 506940 436008
rect 503496 435968 506940 435996
rect 503496 435956 503502 435968
rect 506934 435956 506940 435968
rect 506992 435956 506998 436008
rect 502794 434664 502800 434716
rect 502852 434704 502858 434716
rect 506566 434704 506572 434716
rect 502852 434676 506572 434704
rect 502852 434664 502858 434676
rect 506566 434664 506572 434676
rect 506624 434664 506630 434716
rect 503530 434596 503536 434648
rect 503588 434636 503594 434648
rect 530210 434636 530216 434648
rect 503588 434608 530216 434636
rect 503588 434596 503594 434608
rect 530210 434596 530216 434608
rect 530268 434596 530274 434648
rect 503622 434528 503628 434580
rect 503680 434568 503686 434580
rect 526070 434568 526076 434580
rect 503680 434540 526076 434568
rect 503680 434528 503686 434540
rect 526070 434528 526076 434540
rect 526128 434528 526134 434580
rect 503438 434460 503444 434512
rect 503496 434500 503502 434512
rect 530026 434500 530032 434512
rect 503496 434472 530032 434500
rect 503496 434460 503502 434472
rect 530026 434460 530032 434472
rect 530084 434460 530090 434512
rect 502610 433236 502616 433288
rect 502668 433276 502674 433288
rect 505554 433276 505560 433288
rect 502668 433248 505560 433276
rect 502668 433236 502674 433248
rect 505554 433236 505560 433248
rect 505612 433236 505618 433288
rect 503438 433168 503444 433220
rect 503496 433208 503502 433220
rect 506842 433208 506848 433220
rect 503496 433180 506848 433208
rect 503496 433168 503502 433180
rect 506842 433168 506848 433180
rect 506900 433168 506906 433220
rect 503530 433100 503536 433152
rect 503588 433140 503594 433152
rect 506750 433140 506756 433152
rect 503588 433112 506756 433140
rect 503588 433100 503594 433112
rect 506750 433100 506756 433112
rect 506808 433100 506814 433152
rect 503622 433032 503628 433084
rect 503680 433072 503686 433084
rect 507394 433072 507400 433084
rect 503680 433044 507400 433072
rect 503680 433032 503686 433044
rect 507394 433032 507400 433044
rect 507452 433032 507458 433084
rect 503438 432964 503444 433016
rect 503496 433004 503502 433016
rect 506658 433004 506664 433016
rect 503496 432976 506664 433004
rect 503496 432964 503502 432976
rect 506658 432964 506664 432976
rect 506716 432964 506722 433016
rect 503438 431876 503444 431928
rect 503496 431916 503502 431928
rect 545666 431916 545672 431928
rect 503496 431888 545672 431916
rect 503496 431876 503502 431888
rect 545666 431876 545672 431888
rect 545724 431876 545730 431928
rect 503622 431740 503628 431792
rect 503680 431780 503686 431792
rect 521930 431780 521936 431792
rect 503680 431752 521936 431780
rect 503680 431740 503686 431752
rect 521930 431740 521936 431752
rect 521988 431740 521994 431792
rect 503530 431672 503536 431724
rect 503588 431712 503594 431724
rect 523494 431712 523500 431724
rect 503588 431684 523500 431712
rect 503588 431672 503594 431684
rect 523494 431672 523500 431684
rect 523552 431672 523558 431724
rect 502518 431400 502524 431452
rect 502576 431440 502582 431452
rect 505370 431440 505376 431452
rect 502576 431412 505376 431440
rect 502576 431400 502582 431412
rect 505370 431400 505376 431412
rect 505428 431400 505434 431452
rect 502702 431264 502708 431316
rect 502760 431304 502766 431316
rect 505738 431304 505744 431316
rect 502760 431276 505744 431304
rect 502760 431264 502766 431276
rect 505738 431264 505744 431276
rect 505796 431264 505802 431316
rect 502610 430516 502616 430568
rect 502668 430556 502674 430568
rect 505646 430556 505652 430568
rect 502668 430528 505652 430556
rect 502668 430516 502674 430528
rect 505646 430516 505652 430528
rect 505704 430516 505710 430568
rect 503622 430448 503628 430500
rect 503680 430488 503686 430500
rect 528922 430488 528928 430500
rect 503680 430460 528928 430488
rect 503680 430448 503686 430460
rect 528922 430448 528928 430460
rect 528980 430448 528986 430500
rect 503438 430380 503444 430432
rect 503496 430420 503502 430432
rect 525978 430420 525984 430432
rect 503496 430392 525984 430420
rect 503496 430380 503502 430392
rect 525978 430380 525984 430392
rect 526036 430380 526042 430432
rect 503530 430312 503536 430364
rect 503588 430352 503594 430364
rect 532970 430352 532976 430364
rect 503588 430324 532976 430352
rect 503588 430312 503594 430324
rect 532970 430312 532976 430324
rect 533028 430312 533034 430364
rect 57698 429156 57704 429208
rect 57756 429196 57762 429208
rect 58526 429196 58532 429208
rect 57756 429168 58532 429196
rect 57756 429156 57762 429168
rect 58526 429156 58532 429168
rect 58584 429156 58590 429208
rect 502518 429088 502524 429140
rect 502576 429128 502582 429140
rect 505462 429128 505468 429140
rect 502576 429100 505468 429128
rect 502576 429088 502582 429100
rect 505462 429088 505468 429100
rect 505520 429088 505526 429140
rect 503622 429020 503628 429072
rect 503680 429060 503686 429072
rect 529934 429060 529940 429072
rect 503680 429032 529940 429060
rect 503680 429020 503686 429032
rect 529934 429020 529940 429032
rect 529992 429020 529998 429072
rect 503622 428816 503628 428868
rect 503680 428856 503686 428868
rect 530118 428856 530124 428868
rect 503680 428828 530124 428856
rect 503680 428816 503686 428828
rect 530118 428816 530124 428828
rect 530176 428816 530182 428868
rect 503622 428612 503628 428664
rect 503680 428652 503686 428664
rect 508038 428652 508044 428664
rect 503680 428624 508044 428652
rect 503680 428612 503686 428624
rect 508038 428612 508044 428624
rect 508096 428612 508102 428664
rect 503622 428340 503628 428392
rect 503680 428380 503686 428392
rect 508222 428380 508228 428392
rect 503680 428352 508228 428380
rect 503680 428340 503686 428352
rect 508222 428340 508228 428352
rect 508280 428340 508286 428392
rect 503438 427728 503444 427780
rect 503496 427768 503502 427780
rect 528830 427768 528836 427780
rect 503496 427740 528836 427768
rect 503496 427728 503502 427740
rect 528830 427728 528836 427740
rect 528888 427728 528894 427780
rect 503530 427660 503536 427712
rect 503588 427700 503594 427712
rect 527358 427700 527364 427712
rect 503588 427672 527364 427700
rect 503588 427660 503594 427672
rect 527358 427660 527364 427672
rect 527416 427660 527422 427712
rect 503622 427592 503628 427644
rect 503680 427632 503686 427644
rect 519354 427632 519360 427644
rect 503680 427604 519360 427632
rect 503680 427592 503686 427604
rect 519354 427592 519360 427604
rect 519412 427592 519418 427644
rect 502794 427524 502800 427576
rect 502852 427564 502858 427576
rect 508130 427564 508136 427576
rect 502852 427536 508136 427564
rect 502852 427524 502858 427536
rect 508130 427524 508136 427536
rect 508188 427524 508194 427576
rect 502702 427456 502708 427508
rect 502760 427496 502766 427508
rect 508314 427496 508320 427508
rect 502760 427468 508320 427496
rect 502760 427456 502766 427468
rect 508314 427456 508320 427468
rect 508372 427456 508378 427508
rect 503438 426368 503444 426420
rect 503496 426408 503502 426420
rect 530302 426408 530308 426420
rect 503496 426380 530308 426408
rect 503496 426368 503502 426380
rect 530302 426368 530308 426380
rect 530360 426368 530366 426420
rect 503622 426300 503628 426352
rect 503680 426340 503686 426352
rect 527450 426340 527456 426352
rect 503680 426312 527456 426340
rect 503680 426300 503686 426312
rect 527450 426300 527456 426312
rect 527508 426300 527514 426352
rect 503530 426232 503536 426284
rect 503588 426272 503594 426284
rect 515030 426272 515036 426284
rect 503588 426244 515036 426272
rect 503588 426232 503594 426244
rect 515030 426232 515036 426244
rect 515088 426232 515094 426284
rect 503622 425008 503628 425060
rect 503680 425048 503686 425060
rect 537202 425048 537208 425060
rect 503680 425020 537208 425048
rect 503680 425008 503686 425020
rect 537202 425008 537208 425020
rect 537260 425008 537266 425060
rect 503438 424940 503444 424992
rect 503496 424980 503502 424992
rect 535822 424980 535828 424992
rect 503496 424952 535828 424980
rect 503496 424940 503502 424952
rect 535822 424940 535828 424952
rect 535880 424940 535886 424992
rect 503530 424872 503536 424924
rect 503588 424912 503594 424924
rect 527542 424912 527548 424924
rect 503588 424884 527548 424912
rect 503588 424872 503594 424884
rect 527542 424872 527548 424884
rect 527600 424872 527606 424924
rect 503622 424804 503628 424856
rect 503680 424844 503686 424856
rect 513650 424844 513656 424856
rect 503680 424816 513656 424844
rect 503680 424804 503686 424816
rect 513650 424804 513656 424816
rect 513708 424804 513714 424856
rect 503622 423580 503628 423632
rect 503680 423620 503686 423632
rect 524598 423620 524604 423632
rect 503680 423592 524604 423620
rect 503680 423580 503686 423592
rect 524598 423580 524604 423592
rect 524656 423580 524662 423632
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 14458 422328 14464 422340
rect 3476 422300 14464 422328
rect 3476 422288 3482 422300
rect 14458 422288 14464 422300
rect 14516 422288 14522 422340
rect 43346 420180 43352 420232
rect 43404 420220 43410 420232
rect 46198 420220 46204 420232
rect 43404 420192 46204 420220
rect 43404 420180 43410 420192
rect 46198 420180 46204 420192
rect 46256 420180 46262 420232
rect 54754 400868 54760 400920
rect 54812 400908 54818 400920
rect 57514 400908 57520 400920
rect 54812 400880 57520 400908
rect 54812 400868 54818 400880
rect 57514 400868 57520 400880
rect 57572 400868 57578 400920
rect 37918 392572 37924 392624
rect 37976 392612 37982 392624
rect 51074 392612 51080 392624
rect 37976 392584 51080 392612
rect 37976 392572 37982 392584
rect 51074 392572 51080 392584
rect 51132 392572 51138 392624
rect 60366 391620 60372 391672
rect 60424 391660 60430 391672
rect 62022 391660 62028 391672
rect 60424 391632 62028 391660
rect 60424 391620 60430 391632
rect 62022 391620 62028 391632
rect 62080 391620 62086 391672
rect 498194 390600 498200 390652
rect 498252 390640 498258 390652
rect 500310 390640 500316 390652
rect 498252 390612 500316 390640
rect 498252 390600 498258 390612
rect 500310 390600 500316 390612
rect 500368 390600 500374 390652
rect 325510 390260 325516 390312
rect 325568 390300 325574 390312
rect 503346 390300 503352 390312
rect 325568 390272 503352 390300
rect 325568 390260 325574 390272
rect 503346 390260 503352 390272
rect 503404 390260 503410 390312
rect 14458 390192 14464 390244
rect 14516 390232 14522 390244
rect 96522 390232 96528 390244
rect 14516 390204 96528 390232
rect 14516 390192 14522 390204
rect 96522 390192 96528 390204
rect 96580 390192 96586 390244
rect 306282 390192 306288 390244
rect 306340 390232 306346 390244
rect 501690 390232 501696 390244
rect 306340 390204 501696 390232
rect 306340 390192 306346 390204
rect 501690 390192 501696 390204
rect 501748 390192 501754 390244
rect 58526 390124 58532 390176
rect 58584 390164 58590 390176
rect 144178 390164 144184 390176
rect 58584 390136 144184 390164
rect 58584 390124 58590 390136
rect 144178 390124 144184 390136
rect 144236 390124 144242 390176
rect 343082 390124 343088 390176
rect 343140 390164 343146 390176
rect 544194 390164 544200 390176
rect 343140 390136 544200 390164
rect 343140 390124 343146 390136
rect 544194 390124 544200 390136
rect 544252 390124 544258 390176
rect 57514 390056 57520 390108
rect 57572 390096 57578 390108
rect 220722 390096 220728 390108
rect 57572 390068 220728 390096
rect 57572 390056 57578 390068
rect 220722 390056 220728 390068
rect 220780 390056 220786 390108
rect 346210 390056 346216 390108
rect 346268 390096 346274 390108
rect 545482 390096 545488 390108
rect 346268 390068 545488 390096
rect 346268 390056 346274 390068
rect 545482 390056 545488 390068
rect 545540 390056 545546 390108
rect 62022 389988 62028 390040
rect 62080 390028 62086 390040
rect 273898 390028 273904 390040
rect 62080 390000 273904 390028
rect 62080 389988 62086 390000
rect 273898 389988 273904 390000
rect 273956 389988 273962 390040
rect 308122 389988 308128 390040
rect 308180 390028 308186 390040
rect 500402 390028 500408 390040
rect 308180 390000 500408 390028
rect 308180 389988 308186 390000
rect 500402 389988 500408 390000
rect 500460 389988 500466 390040
rect 51810 389920 51816 389972
rect 51868 389960 51874 389972
rect 274726 389960 274732 389972
rect 51868 389932 274732 389960
rect 51868 389920 51874 389932
rect 274726 389920 274732 389932
rect 274784 389920 274790 389972
rect 485774 389920 485780 389972
rect 485832 389960 485838 389972
rect 501874 389960 501880 389972
rect 485832 389932 501880 389960
rect 485832 389920 485838 389932
rect 501874 389920 501880 389932
rect 501932 389920 501938 389972
rect 46198 389852 46204 389904
rect 46256 389892 46262 389904
rect 294598 389892 294604 389904
rect 46256 389864 294604 389892
rect 46256 389852 46262 389864
rect 294598 389852 294604 389864
rect 294656 389852 294662 389904
rect 398098 389852 398104 389904
rect 398156 389892 398162 389904
rect 498194 389892 498200 389904
rect 398156 389864 498200 389892
rect 398156 389852 398162 389864
rect 498194 389852 498200 389864
rect 498252 389852 498258 389904
rect 51074 389784 51080 389836
rect 51132 389824 51138 389836
rect 326338 389824 326344 389836
rect 51132 389796 326344 389824
rect 51132 389784 51138 389796
rect 326338 389784 326344 389796
rect 326396 389784 326402 389836
rect 360470 389784 360476 389836
rect 360528 389824 360534 389836
rect 525886 389824 525892 389836
rect 360528 389796 525892 389824
rect 360528 389784 360534 389796
rect 525886 389784 525892 389796
rect 525944 389784 525950 389836
rect 309778 389104 309784 389156
rect 309836 389144 309842 389156
rect 537754 389144 537760 389156
rect 309836 389116 537760 389144
rect 309836 389104 309842 389116
rect 537754 389104 537760 389116
rect 537812 389104 537818 389156
rect 311158 389036 311164 389088
rect 311216 389076 311222 389088
rect 537570 389076 537576 389088
rect 311216 389048 537576 389076
rect 311216 389036 311222 389048
rect 537570 389036 537576 389048
rect 537628 389036 537634 389088
rect 346302 388968 346308 389020
rect 346360 389008 346366 389020
rect 543918 389008 543924 389020
rect 346360 388980 543924 389008
rect 346360 388968 346366 388980
rect 543918 388968 543924 388980
rect 543976 388968 543982 389020
rect 349798 388900 349804 388952
rect 349856 388940 349862 388952
rect 505830 388940 505836 388952
rect 349856 388912 505836 388940
rect 349856 388900 349862 388912
rect 505830 388900 505836 388912
rect 505888 388900 505894 388952
rect 319714 388832 319720 388884
rect 319772 388872 319778 388884
rect 398098 388872 398104 388884
rect 319772 388844 398104 388872
rect 319772 388832 319778 388844
rect 398098 388832 398104 388844
rect 398156 388832 398162 388884
rect 400306 388832 400312 388884
rect 400364 388872 400370 388884
rect 545574 388872 545580 388884
rect 400364 388844 545580 388872
rect 400364 388832 400370 388844
rect 545574 388832 545580 388844
rect 545632 388832 545638 388884
rect 398834 388492 398840 388544
rect 398892 388532 398898 388544
rect 499942 388532 499948 388544
rect 398892 388504 499948 388532
rect 398892 388492 398898 388504
rect 499942 388492 499948 388504
rect 500000 388492 500006 388544
rect 11698 388424 11704 388476
rect 11756 388464 11762 388476
rect 95142 388464 95148 388476
rect 11756 388436 95148 388464
rect 11756 388424 11762 388436
rect 95142 388424 95148 388436
rect 95200 388424 95206 388476
rect 359642 388424 359648 388476
rect 359700 388464 359706 388476
rect 509510 388464 509516 388476
rect 359700 388436 509516 388464
rect 359700 388424 359706 388436
rect 509510 388424 509516 388436
rect 509568 388424 509574 388476
rect 96522 387744 96528 387796
rect 96580 387784 96586 387796
rect 339310 387784 339316 387796
rect 96580 387756 339316 387784
rect 96580 387744 96586 387756
rect 339310 387744 339316 387756
rect 339368 387744 339374 387796
rect 343634 387744 343640 387796
rect 343692 387784 343698 387796
rect 344554 387784 344560 387796
rect 343692 387756 344560 387784
rect 343692 387744 343698 387756
rect 344554 387744 344560 387756
rect 344612 387784 344618 387796
rect 546586 387784 546592 387796
rect 344612 387756 546592 387784
rect 344612 387744 344618 387756
rect 546586 387744 546592 387756
rect 546644 387744 546650 387796
rect 95142 387676 95148 387728
rect 95200 387716 95206 387728
rect 337562 387716 337568 387728
rect 95200 387688 337568 387716
rect 95200 387676 95206 387688
rect 337562 387676 337568 387688
rect 337620 387716 337626 387728
rect 544102 387716 544108 387728
rect 337620 387688 544108 387716
rect 337620 387676 337626 387688
rect 544102 387676 544108 387688
rect 544160 387676 544166 387728
rect 314838 387608 314844 387660
rect 314896 387648 314902 387660
rect 315298 387648 315304 387660
rect 314896 387620 315304 387648
rect 314896 387608 314902 387620
rect 315298 387608 315304 387620
rect 315356 387648 315362 387660
rect 539226 387648 539232 387660
rect 315356 387620 539232 387648
rect 315356 387608 315362 387620
rect 539226 387608 539232 387620
rect 539284 387608 539290 387660
rect 37090 387540 37096 387592
rect 37148 387580 37154 387592
rect 89714 387580 89720 387592
rect 37148 387552 89720 387580
rect 37148 387540 37154 387552
rect 89714 387540 89720 387552
rect 89772 387540 89778 387592
rect 292114 387540 292120 387592
rect 292172 387580 292178 387592
rect 359642 387580 359648 387592
rect 292172 387552 359648 387580
rect 292172 387540 292178 387552
rect 359642 387540 359648 387552
rect 359700 387540 359706 387592
rect 32766 387472 32772 387524
rect 32824 387512 32830 387524
rect 91186 387512 91192 387524
rect 32824 387484 91192 387512
rect 32824 387472 32830 387484
rect 91186 387472 91192 387484
rect 91244 387472 91250 387524
rect 221826 387472 221832 387524
rect 221884 387512 221890 387524
rect 343634 387512 343640 387524
rect 221884 387484 343640 387512
rect 221884 387472 221890 387484
rect 343634 387472 343640 387484
rect 343692 387472 343698 387524
rect 348418 387472 348424 387524
rect 348476 387512 348482 387524
rect 547966 387512 547972 387524
rect 348476 387484 547972 387512
rect 348476 387472 348482 387484
rect 547966 387472 547972 387484
rect 548024 387472 548030 387524
rect 45462 387404 45468 387456
rect 45520 387444 45526 387456
rect 106182 387444 106188 387456
rect 45520 387416 106188 387444
rect 45520 387404 45526 387416
rect 106182 387404 106188 387416
rect 106240 387444 106246 387456
rect 327074 387444 327080 387456
rect 106240 387416 327080 387444
rect 106240 387404 106246 387416
rect 327074 387404 327080 387416
rect 327132 387404 327138 387456
rect 85574 387336 85580 387388
rect 85632 387376 85638 387388
rect 86862 387376 86868 387388
rect 85632 387348 86868 387376
rect 85632 387336 85638 387348
rect 86862 387336 86868 387348
rect 86920 387376 86926 387388
rect 328822 387376 328828 387388
rect 86920 387348 328828 387376
rect 86920 387336 86926 387348
rect 328822 387336 328828 387348
rect 328880 387336 328886 387388
rect 86954 387268 86960 387320
rect 87012 387308 87018 387320
rect 88242 387308 88248 387320
rect 87012 387280 88248 387308
rect 87012 387268 87018 387280
rect 88242 387268 88248 387280
rect 88300 387308 88306 387320
rect 330570 387308 330576 387320
rect 88300 387280 330576 387308
rect 88300 387268 88306 387280
rect 330570 387268 330576 387280
rect 330628 387268 330634 387320
rect 31570 387200 31576 387252
rect 31628 387240 31634 387252
rect 89622 387240 89628 387252
rect 31628 387212 89628 387240
rect 31628 387200 31634 387212
rect 89622 387200 89628 387212
rect 89680 387240 89686 387252
rect 332318 387240 332324 387252
rect 89680 387212 332324 387240
rect 89680 387200 89686 387212
rect 332318 387200 332324 387212
rect 332376 387200 332382 387252
rect 341518 387200 341524 387252
rect 341576 387240 341582 387252
rect 360194 387240 360200 387252
rect 341576 387212 360200 387240
rect 341576 387200 341582 387212
rect 360194 387200 360200 387212
rect 360252 387200 360258 387252
rect 27154 387132 27160 387184
rect 27212 387172 27218 387184
rect 85574 387172 85580 387184
rect 27212 387144 85580 387172
rect 27212 387132 27218 387144
rect 85574 387132 85580 387144
rect 85632 387132 85638 387184
rect 89714 387132 89720 387184
rect 89772 387172 89778 387184
rect 91002 387172 91008 387184
rect 89772 387144 91008 387172
rect 89772 387132 89778 387144
rect 91002 387132 91008 387144
rect 91060 387172 91066 387184
rect 334066 387172 334072 387184
rect 91060 387144 334072 387172
rect 91060 387132 91066 387144
rect 334066 387132 334072 387144
rect 334124 387132 334130 387184
rect 359734 387132 359740 387184
rect 359792 387172 359798 387184
rect 403986 387172 403992 387184
rect 359792 387144 403992 387172
rect 359792 387132 359798 387144
rect 403986 387132 403992 387144
rect 404044 387132 404050 387184
rect 26142 387064 26148 387116
rect 26200 387104 26206 387116
rect 86954 387104 86960 387116
rect 26200 387076 86960 387104
rect 26200 387064 26206 387076
rect 86954 387064 86960 387076
rect 87012 387064 87018 387116
rect 91186 387064 91192 387116
rect 91244 387104 91250 387116
rect 92382 387104 92388 387116
rect 91244 387076 92388 387104
rect 91244 387064 91250 387076
rect 92382 387064 92388 387076
rect 92440 387104 92446 387116
rect 335814 387104 335820 387116
rect 92440 387076 335820 387104
rect 92440 387064 92446 387076
rect 335814 387064 335820 387076
rect 335872 387064 335878 387116
rect 339310 387064 339316 387116
rect 339368 387104 339374 387116
rect 360102 387104 360108 387116
rect 339368 387076 360108 387104
rect 339368 387064 339374 387076
rect 360102 387064 360108 387076
rect 360160 387064 360166 387116
rect 360378 387064 360384 387116
rect 360436 387104 360442 387116
rect 419718 387104 419724 387116
rect 360436 387076 419724 387104
rect 360436 387064 360442 387076
rect 419718 387064 419724 387076
rect 419776 387064 419782 387116
rect 293862 386996 293868 387048
rect 293920 387036 293926 387048
rect 355962 387036 355968 387048
rect 293920 387008 355968 387036
rect 293920 386996 293926 387008
rect 355962 386996 355968 387008
rect 356020 387036 356026 387048
rect 360470 387036 360476 387048
rect 356020 387008 360476 387036
rect 356020 386996 356026 387008
rect 360470 386996 360476 387008
rect 360528 386996 360534 387048
rect 360102 386520 360108 386572
rect 360160 386560 360166 386572
rect 394602 386560 394608 386572
rect 360160 386532 394608 386560
rect 360160 386520 360166 386532
rect 394602 386520 394608 386532
rect 394660 386520 394666 386572
rect 360194 386452 360200 386504
rect 360252 386492 360258 386504
rect 395982 386492 395988 386504
rect 360252 386464 395988 386492
rect 360252 386452 360258 386464
rect 395982 386452 395988 386464
rect 396040 386452 396046 386504
rect 302878 386384 302884 386436
rect 302936 386424 302942 386436
rect 498194 386424 498200 386436
rect 302936 386396 498200 386424
rect 302936 386384 302942 386396
rect 498194 386384 498200 386396
rect 498252 386384 498258 386436
rect 220722 386316 220728 386368
rect 220780 386356 220786 386368
rect 227714 386356 227720 386368
rect 220780 386328 227720 386356
rect 220780 386316 220786 386328
rect 227714 386316 227720 386328
rect 227772 386316 227778 386368
rect 394602 386316 394608 386368
rect 394660 386356 394666 386368
rect 544010 386356 544016 386368
rect 394660 386328 544016 386356
rect 394660 386316 394666 386328
rect 544010 386316 544016 386328
rect 544068 386316 544074 386368
rect 395982 386248 395988 386300
rect 396040 386288 396046 386300
rect 545390 386288 545396 386300
rect 396040 386260 545396 386288
rect 396040 386248 396046 386260
rect 545390 386248 545396 386260
rect 545448 386248 545454 386300
rect 466362 385636 466368 385688
rect 466420 385676 466426 385688
rect 485774 385676 485780 385688
rect 466420 385648 485780 385676
rect 466420 385636 466426 385648
rect 485774 385636 485780 385648
rect 485832 385636 485838 385688
rect 282086 384956 282092 385008
rect 282144 384996 282150 385008
rect 491386 384996 491392 385008
rect 282144 384968 491392 384996
rect 282144 384956 282150 384968
rect 491386 384956 491392 384968
rect 491444 384956 491450 385008
rect 355962 384888 355968 384940
rect 356020 384928 356026 384940
rect 542722 384928 542728 384940
rect 356020 384900 542728 384928
rect 356020 384888 356026 384900
rect 542722 384888 542728 384900
rect 542780 384888 542786 384940
rect 357342 384820 357348 384872
rect 357400 384860 357406 384872
rect 542814 384860 542820 384872
rect 357400 384832 542820 384860
rect 357400 384820 357406 384832
rect 542814 384820 542820 384832
rect 542872 384820 542878 384872
rect 274726 384344 274732 384396
rect 274784 384384 274790 384396
rect 287698 384384 287704 384396
rect 274784 384356 287704 384384
rect 274784 384344 274790 384356
rect 287698 384344 287704 384356
rect 287756 384344 287762 384396
rect 498194 384344 498200 384396
rect 498252 384384 498258 384396
rect 529934 384384 529940 384396
rect 498252 384356 529940 384384
rect 498252 384344 498258 384356
rect 529934 384344 529940 384356
rect 529992 384344 529998 384396
rect 239950 384276 239956 384328
rect 240008 384316 240014 384328
rect 580350 384316 580356 384328
rect 240008 384288 580356 384316
rect 240008 384276 240014 384288
rect 580350 384276 580356 384288
rect 580408 384276 580414 384328
rect 234614 383664 234620 383716
rect 234672 383704 234678 383716
rect 313918 383704 313924 383716
rect 234672 383676 313924 383704
rect 234672 383664 234678 383676
rect 313918 383664 313924 383676
rect 313976 383664 313982 383716
rect 498838 383664 498844 383716
rect 498896 383704 498902 383716
rect 501782 383704 501788 383716
rect 498896 383676 501788 383704
rect 498896 383664 498902 383676
rect 501782 383664 501788 383676
rect 501840 383664 501846 383716
rect 294598 382916 294604 382968
rect 294656 382956 294662 382968
rect 308490 382956 308496 382968
rect 294656 382928 308496 382956
rect 294656 382916 294662 382928
rect 308490 382916 308496 382928
rect 308548 382916 308554 382968
rect 445662 382916 445668 382968
rect 445720 382956 445726 382968
rect 466362 382956 466368 382968
rect 445720 382928 466368 382956
rect 445720 382916 445726 382928
rect 466362 382916 466368 382928
rect 466420 382916 466426 382968
rect 273898 382236 273904 382288
rect 273956 382276 273962 382288
rect 276658 382276 276664 382288
rect 273956 382248 276664 382276
rect 273956 382236 273962 382248
rect 276658 382236 276664 382248
rect 276716 382236 276722 382288
rect 529934 382236 529940 382288
rect 529992 382276 529998 382288
rect 531222 382276 531228 382288
rect 529992 382248 531228 382276
rect 529992 382236 529998 382248
rect 531222 382236 531228 382248
rect 531280 382276 531286 382288
rect 532786 382276 532792 382288
rect 531280 382248 532792 382276
rect 531280 382236 531286 382248
rect 532786 382236 532792 382248
rect 532844 382236 532850 382288
rect 240042 382168 240048 382220
rect 240100 382208 240106 382220
rect 535546 382208 535552 382220
rect 240100 382180 535552 382208
rect 240100 382168 240106 382180
rect 535546 382168 535552 382180
rect 535604 382168 535610 382220
rect 266354 382100 266360 382152
rect 266412 382140 266418 382152
rect 527266 382140 527272 382152
rect 266412 382112 527272 382140
rect 266412 382100 266418 382112
rect 527266 382100 527272 382112
rect 527324 382100 527330 382152
rect 227714 380128 227720 380180
rect 227772 380168 227778 380180
rect 235994 380168 236000 380180
rect 227772 380140 236000 380168
rect 227772 380128 227778 380140
rect 235994 380128 236000 380140
rect 236052 380128 236058 380180
rect 282546 378836 282552 378888
rect 282604 378876 282610 378888
rect 541250 378876 541256 378888
rect 282604 378848 541256 378876
rect 282604 378836 282610 378848
rect 541250 378836 541256 378848
rect 541308 378836 541314 378888
rect 144178 378768 144184 378820
rect 144236 378808 144242 378820
rect 146938 378808 146944 378820
rect 144236 378780 146944 378808
rect 144236 378768 144242 378780
rect 146938 378768 146944 378780
rect 146996 378768 147002 378820
rect 282270 378768 282276 378820
rect 282328 378808 282334 378820
rect 541342 378808 541348 378820
rect 282328 378780 541348 378808
rect 282328 378768 282334 378780
rect 541342 378768 541348 378780
rect 541400 378768 541406 378820
rect 239306 378156 239312 378208
rect 239364 378196 239370 378208
rect 580166 378196 580172 378208
rect 239364 378168 580172 378196
rect 239364 378156 239370 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 436738 377408 436744 377460
rect 436796 377448 436802 377460
rect 445662 377448 445668 377460
rect 436796 377420 445668 377448
rect 436796 377408 436802 377420
rect 445662 377408 445668 377420
rect 445720 377408 445726 377460
rect 234614 376660 234620 376712
rect 234672 376700 234678 376712
rect 530762 376700 530768 376712
rect 234672 376672 530768 376700
rect 234672 376660 234678 376672
rect 530762 376660 530768 376672
rect 530820 376660 530826 376712
rect 485958 376592 485964 376644
rect 486016 376632 486022 376644
rect 549254 376632 549260 376644
rect 486016 376604 549260 376632
rect 486016 376592 486022 376604
rect 549254 376592 549260 376604
rect 549312 376592 549318 376644
rect 282454 376048 282460 376100
rect 282512 376088 282518 376100
rect 539962 376088 539968 376100
rect 282512 376060 539968 376088
rect 282512 376048 282518 376060
rect 539962 376048 539968 376060
rect 540020 376048 540026 376100
rect 231210 375980 231216 376032
rect 231268 376020 231274 376032
rect 537662 376020 537668 376032
rect 231268 375992 537668 376020
rect 231268 375980 231274 375992
rect 537662 375980 537668 375992
rect 537720 375980 537726 376032
rect 235994 375368 236000 375420
rect 236052 375408 236058 375420
rect 238846 375408 238852 375420
rect 236052 375380 238852 375408
rect 236052 375368 236058 375380
rect 238846 375368 238852 375380
rect 238904 375368 238910 375420
rect 287698 375300 287704 375352
rect 287756 375340 287762 375352
rect 294598 375340 294604 375352
rect 287756 375312 294604 375340
rect 287756 375300 287762 375312
rect 294598 375300 294604 375312
rect 294656 375300 294662 375352
rect 276014 373940 276020 373992
rect 276072 373980 276078 373992
rect 511442 373980 511448 373992
rect 276072 373952 511448 373980
rect 276072 373940 276078 373952
rect 511442 373940 511448 373952
rect 511500 373940 511506 373992
rect 238846 373260 238852 373312
rect 238904 373300 238910 373312
rect 264974 373300 264980 373312
rect 238904 373272 264980 373300
rect 238904 373260 238910 373272
rect 264974 373260 264980 373272
rect 265032 373260 265038 373312
rect 97902 371832 97908 371884
rect 97960 371872 97966 371884
rect 341518 371872 341524 371884
rect 97960 371844 341524 371872
rect 97960 371832 97966 371844
rect 341518 371832 341524 371844
rect 341576 371832 341582 371884
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 97902 371260 97908 371272
rect 3476 371232 97908 371260
rect 3476 371220 3482 371232
rect 97902 371220 97908 371232
rect 97960 371220 97966 371272
rect 264974 369112 264980 369164
rect 265032 369152 265038 369164
rect 276014 369152 276020 369164
rect 265032 369124 276020 369152
rect 265032 369112 265038 369124
rect 276014 369112 276020 369124
rect 276072 369112 276078 369164
rect 359366 369112 359372 369164
rect 359424 369152 359430 369164
rect 435450 369152 435456 369164
rect 359424 369124 435456 369152
rect 359424 369112 359430 369124
rect 435450 369112 435456 369124
rect 435508 369112 435514 369164
rect 495434 368772 495440 368824
rect 495492 368812 495498 368824
rect 498838 368812 498844 368824
rect 495492 368784 498844 368812
rect 495492 368772 495498 368784
rect 498838 368772 498844 368784
rect 498896 368772 498902 368824
rect 358354 367752 358360 367804
rect 358412 367792 358418 367804
rect 479150 367792 479156 367804
rect 358412 367764 479156 367792
rect 358412 367752 358418 367764
rect 479150 367752 479156 367764
rect 479208 367752 479214 367804
rect 276014 366664 276020 366716
rect 276072 366704 276078 366716
rect 293586 366704 293592 366716
rect 276072 366676 293592 366704
rect 276072 366664 276078 366676
rect 293586 366664 293592 366676
rect 293644 366664 293650 366716
rect 294598 366664 294604 366716
rect 294656 366704 294662 366716
rect 306006 366704 306012 366716
rect 294656 366676 306012 366704
rect 294656 366664 294662 366676
rect 306006 366664 306012 366676
rect 306064 366664 306070 366716
rect 57422 366596 57428 366648
rect 57480 366636 57486 366648
rect 341518 366636 341524 366648
rect 57480 366608 341524 366636
rect 57480 366596 57486 366608
rect 341518 366596 341524 366608
rect 341576 366596 341582 366648
rect 29730 366528 29736 366580
rect 29788 366568 29794 366580
rect 333238 366568 333244 366580
rect 29788 366540 333244 366568
rect 29788 366528 29794 366540
rect 333238 366528 333244 366540
rect 333296 366528 333302 366580
rect 356698 366528 356704 366580
rect 356756 366568 356762 366580
rect 452930 366568 452936 366580
rect 356756 366540 452936 366568
rect 356756 366528 356762 366540
rect 452930 366528 452936 366540
rect 452988 366528 452994 366580
rect 29822 366460 29828 366512
rect 29880 366500 29886 366512
rect 358078 366500 358084 366512
rect 29880 366472 358084 366500
rect 29880 366460 29886 366472
rect 358078 366460 358084 366472
rect 358136 366460 358142 366512
rect 487798 366460 487804 366512
rect 487856 366500 487862 366512
rect 495434 366500 495440 366512
rect 487856 366472 495440 366500
rect 487856 366460 487862 366472
rect 495434 366460 495440 366472
rect 495492 366460 495498 366512
rect 43530 366392 43536 366444
rect 43588 366432 43594 366444
rect 502334 366432 502340 366444
rect 43588 366404 502340 366432
rect 43588 366392 43594 366404
rect 502334 366392 502340 366404
rect 502392 366392 502398 366444
rect 42242 366324 42248 366376
rect 42300 366364 42306 366376
rect 501138 366364 501144 366376
rect 42300 366336 501144 366364
rect 42300 366324 42306 366336
rect 501138 366324 501144 366336
rect 501196 366324 501202 366376
rect 420914 365032 420920 365084
rect 420972 365072 420978 365084
rect 436738 365072 436744 365084
rect 420972 365044 436744 365072
rect 420972 365032 420978 365044
rect 436738 365032 436744 365044
rect 436796 365032 436802 365084
rect 43622 364964 43628 365016
rect 43680 365004 43686 365016
rect 502426 365004 502432 365016
rect 43680 364976 502432 365004
rect 43680 364964 43686 364976
rect 502426 364964 502432 364976
rect 502484 364964 502490 365016
rect 146938 364352 146944 364404
rect 146996 364392 147002 364404
rect 153838 364392 153844 364404
rect 146996 364364 153844 364392
rect 146996 364352 147002 364364
rect 153838 364352 153844 364364
rect 153896 364352 153902 364404
rect 60274 364216 60280 364268
rect 60332 364256 60338 364268
rect 341702 364256 341708 364268
rect 60332 364228 341708 364256
rect 60332 364216 60338 364228
rect 341702 364216 341708 364228
rect 341760 364216 341766 364268
rect 46658 364148 46664 364200
rect 46716 364188 46722 364200
rect 333422 364188 333428 364200
rect 46716 364160 333428 364188
rect 46716 364148 46722 364160
rect 333422 364148 333428 364160
rect 333480 364148 333486 364200
rect 42426 364080 42432 364132
rect 42484 364120 42490 364132
rect 335998 364120 336004 364132
rect 42484 364092 336004 364120
rect 42484 364080 42490 364092
rect 335998 364080 336004 364092
rect 336056 364080 336062 364132
rect 40954 364012 40960 364064
rect 41012 364052 41018 364064
rect 338758 364052 338764 364064
rect 41012 364024 338764 364052
rect 41012 364012 41018 364024
rect 338758 364012 338764 364024
rect 338816 364012 338822 364064
rect 47394 363944 47400 363996
rect 47452 363984 47458 363996
rect 347038 363984 347044 363996
rect 47452 363956 347044 363984
rect 47452 363944 47458 363956
rect 347038 363944 347044 363956
rect 347096 363944 347102 363996
rect 29914 363876 29920 363928
rect 29972 363916 29978 363928
rect 333330 363916 333336 363928
rect 29972 363888 333336 363916
rect 29972 363876 29978 363888
rect 333330 363876 333336 363888
rect 333388 363876 333394 363928
rect 39942 363808 39948 363860
rect 40000 363848 40006 363860
rect 347130 363848 347136 363860
rect 40000 363820 347136 363848
rect 40000 363808 40006 363820
rect 347130 363808 347136 363820
rect 347188 363808 347194 363860
rect 43714 363740 43720 363792
rect 43772 363780 43778 363792
rect 359458 363780 359464 363792
rect 43772 363752 359464 363780
rect 43772 363740 43778 363752
rect 359458 363740 359464 363752
rect 359516 363740 359522 363792
rect 477494 363740 477500 363792
rect 477552 363780 477558 363792
rect 487798 363780 487804 363792
rect 477552 363752 487804 363780
rect 477552 363740 477558 363752
rect 487798 363740 487804 363752
rect 487856 363740 487862 363792
rect 42334 363672 42340 363724
rect 42392 363712 42398 363724
rect 499666 363712 499672 363724
rect 42392 363684 499672 363712
rect 42392 363672 42398 363684
rect 499666 363672 499672 363684
rect 499724 363672 499730 363724
rect 45094 363604 45100 363656
rect 45152 363644 45158 363656
rect 505094 363644 505100 363656
rect 45152 363616 505100 363644
rect 45152 363604 45158 363616
rect 505094 363604 505100 363616
rect 505152 363604 505158 363656
rect 45186 362176 45192 362228
rect 45244 362216 45250 362228
rect 503898 362216 503904 362228
rect 45244 362188 503904 362216
rect 45244 362176 45250 362188
rect 503898 362176 503904 362188
rect 503956 362176 503962 362228
rect 60458 361360 60464 361412
rect 60516 361400 60522 361412
rect 336366 361400 336372 361412
rect 60516 361372 336372 361400
rect 60516 361360 60522 361372
rect 336366 361360 336372 361372
rect 336424 361360 336430 361412
rect 59262 361292 59268 361344
rect 59320 361332 59326 361344
rect 336182 361332 336188 361344
rect 59320 361304 336188 361332
rect 59320 361292 59326 361304
rect 336182 361292 336188 361304
rect 336240 361292 336246 361344
rect 58618 361224 58624 361276
rect 58676 361264 58682 361276
rect 336274 361264 336280 361276
rect 58676 361236 336280 361264
rect 58676 361224 58682 361236
rect 336274 361224 336280 361236
rect 336332 361224 336338 361276
rect 57882 361156 57888 361208
rect 57940 361196 57946 361208
rect 338850 361196 338856 361208
rect 57940 361168 338856 361196
rect 57940 361156 57946 361168
rect 338850 361156 338856 361168
rect 338908 361156 338914 361208
rect 41046 361088 41052 361140
rect 41104 361128 41110 361140
rect 336090 361128 336096 361140
rect 41104 361100 336096 361128
rect 41104 361088 41110 361100
rect 336090 361088 336096 361100
rect 336148 361088 336154 361140
rect 25774 361020 25780 361072
rect 25832 361060 25838 361072
rect 347222 361060 347228 361072
rect 25832 361032 347228 361060
rect 25832 361020 25838 361032
rect 347222 361020 347228 361032
rect 347280 361020 347286 361072
rect 25958 360952 25964 361004
rect 26016 360992 26022 361004
rect 355318 360992 355324 361004
rect 26016 360964 355324 360992
rect 26016 360952 26022 360964
rect 355318 360952 355324 360964
rect 355376 360952 355382 361004
rect 25590 360884 25596 360936
rect 25648 360924 25654 360936
rect 359550 360924 359556 360936
rect 25648 360896 359556 360924
rect 25648 360884 25654 360896
rect 359550 360884 359556 360896
rect 359608 360884 359614 360936
rect 408494 360884 408500 360936
rect 408552 360924 408558 360936
rect 420914 360924 420920 360936
rect 408552 360896 420920 360924
rect 408552 360884 408558 360896
rect 420914 360884 420920 360896
rect 420972 360884 420978 360936
rect 45278 360816 45284 360868
rect 45336 360856 45342 360868
rect 503806 360856 503812 360868
rect 45336 360828 503812 360856
rect 45336 360816 45342 360828
rect 503806 360816 503812 360828
rect 503864 360816 503870 360868
rect 253198 359524 253204 359576
rect 253256 359564 253262 359576
rect 430206 359564 430212 359576
rect 253256 359536 430212 359564
rect 253256 359524 253262 359536
rect 430206 359524 430212 359536
rect 430264 359524 430270 359576
rect 40862 359456 40868 359508
rect 40920 359496 40926 359508
rect 502518 359496 502524 359508
rect 40920 359468 502524 359496
rect 40920 359456 40926 359468
rect 502518 359456 502524 359468
rect 502576 359456 502582 359508
rect 252462 358844 252468 358896
rect 252520 358884 252526 358896
rect 289078 358884 289084 358896
rect 252520 358856 289084 358884
rect 252520 358844 252526 358856
rect 289078 358844 289084 358856
rect 289136 358844 289142 358896
rect 252370 358776 252376 358828
rect 252428 358816 252434 358828
rect 294598 358816 294604 358828
rect 252428 358788 294604 358816
rect 252428 358776 252434 358788
rect 294598 358776 294604 358788
rect 294656 358776 294662 358828
rect 271782 358640 271788 358692
rect 271840 358680 271846 358692
rect 282914 358680 282920 358692
rect 271840 358652 282920 358680
rect 271840 358640 271846 358652
rect 282914 358640 282920 358652
rect 282972 358640 282978 358692
rect 272426 358572 272432 358624
rect 272484 358612 272490 358624
rect 472158 358612 472164 358624
rect 272484 358584 472164 358612
rect 272484 358572 272490 358584
rect 472158 358572 472164 358584
rect 472216 358572 472222 358624
rect 273346 358504 273352 358556
rect 273404 358544 273410 358556
rect 473906 358544 473912 358556
rect 273404 358516 473912 358544
rect 273404 358504 273410 358516
rect 473906 358504 473912 358516
rect 473964 358504 473970 358556
rect 274266 358436 274272 358488
rect 274324 358476 274330 358488
rect 475654 358476 475660 358488
rect 274324 358448 475660 358476
rect 274324 358436 274330 358448
rect 475654 358436 475660 358448
rect 475712 358436 475718 358488
rect 275186 358368 275192 358420
rect 275244 358408 275250 358420
rect 477402 358408 477408 358420
rect 275244 358380 477408 358408
rect 275244 358368 275250 358380
rect 477402 358368 477408 358380
rect 477460 358368 477466 358420
rect 60182 358300 60188 358352
rect 60240 358340 60246 358352
rect 302234 358340 302240 358352
rect 60240 358312 302240 358340
rect 60240 358300 60246 358312
rect 302234 358300 302240 358312
rect 302292 358300 302298 358352
rect 57330 358232 57336 358284
rect 57388 358272 57394 358284
rect 338942 358272 338948 358284
rect 57388 358244 338948 358272
rect 57388 358232 57394 358244
rect 338942 358232 338948 358244
rect 339000 358232 339006 358284
rect 56226 358164 56232 358216
rect 56284 358204 56290 358216
rect 347314 358204 347320 358216
rect 56284 358176 347320 358204
rect 56284 358164 56290 358176
rect 347314 358164 347320 358176
rect 347372 358164 347378 358216
rect 54570 358096 54576 358148
rect 54628 358136 54634 358148
rect 349890 358136 349896 358148
rect 54628 358108 349896 358136
rect 54628 358096 54634 358108
rect 349890 358096 349896 358108
rect 349948 358096 349954 358148
rect 53282 358028 53288 358080
rect 53340 358068 53346 358080
rect 349798 358068 349804 358080
rect 53340 358040 349804 358068
rect 53340 358028 53346 358040
rect 349798 358028 349804 358040
rect 349856 358028 349862 358080
rect 402238 358028 402244 358080
rect 402296 358068 402302 358080
rect 408494 358068 408500 358080
rect 402296 358040 408500 358068
rect 402296 358028 402302 358040
rect 408494 358028 408500 358040
rect 408552 358028 408558 358080
rect 474642 357620 474648 357672
rect 474700 357660 474706 357672
rect 477494 357660 477500 357672
rect 474700 357632 477500 357660
rect 474700 357620 474706 357632
rect 477494 357620 477500 357632
rect 477552 357620 477558 357672
rect 271782 357416 271788 357468
rect 271840 357456 271846 357468
rect 303614 357456 303620 357468
rect 271840 357428 303620 357456
rect 271840 357416 271846 357428
rect 303614 357416 303620 357428
rect 303672 357416 303678 357468
rect 260466 356804 260472 356856
rect 260524 356844 260530 356856
rect 449434 356844 449440 356856
rect 260524 356816 449440 356844
rect 260524 356804 260530 356816
rect 449434 356804 449440 356816
rect 449492 356804 449498 356856
rect 261386 356736 261392 356788
rect 261444 356776 261450 356788
rect 451182 356776 451188 356788
rect 261444 356748 451188 356776
rect 261444 356736 261450 356748
rect 451182 356736 451188 356748
rect 451240 356736 451246 356788
rect 45370 356668 45376 356720
rect 45428 356708 45434 356720
rect 502702 356708 502708 356720
rect 45428 356680 502708 356708
rect 45428 356668 45434 356680
rect 502702 356668 502708 356680
rect 502760 356668 502766 356720
rect 238386 355920 238392 355972
rect 238444 355960 238450 355972
rect 284294 355960 284300 355972
rect 238444 355932 284300 355960
rect 238444 355920 238450 355932
rect 284294 355920 284300 355932
rect 284352 355920 284358 355972
rect 276014 355852 276020 355904
rect 276072 355892 276078 355904
rect 532694 355892 532700 355904
rect 276072 355864 532700 355892
rect 276072 355852 276078 355864
rect 532694 355852 532700 355864
rect 532752 355852 532758 355904
rect 269022 355784 269028 355836
rect 269080 355824 269086 355836
rect 534074 355824 534080 355836
rect 269080 355796 534080 355824
rect 269080 355784 269086 355796
rect 534074 355784 534080 355796
rect 534132 355784 534138 355836
rect 60090 355716 60096 355768
rect 60148 355756 60154 355768
rect 341886 355756 341892 355768
rect 60148 355728 341892 355756
rect 60148 355716 60154 355728
rect 341886 355716 341892 355728
rect 341944 355716 341950 355768
rect 58710 355648 58716 355700
rect 58768 355688 58774 355700
rect 341794 355688 341800 355700
rect 58768 355660 341800 355688
rect 58768 355648 58774 355660
rect 341794 355648 341800 355660
rect 341852 355648 341858 355700
rect 57238 355580 57244 355632
rect 57296 355620 57302 355632
rect 344370 355620 344376 355632
rect 57296 355592 344376 355620
rect 57296 355580 57302 355592
rect 344370 355580 344376 355592
rect 344428 355580 344434 355632
rect 238202 355512 238208 355564
rect 238260 355552 238266 355564
rect 529934 355552 529940 355564
rect 238260 355524 529940 355552
rect 238260 355512 238266 355524
rect 529934 355512 529940 355524
rect 529992 355512 529998 355564
rect 53098 355444 53104 355496
rect 53156 355484 53162 355496
rect 344278 355484 344284 355496
rect 53156 355456 344284 355484
rect 53156 355444 53162 355456
rect 344278 355444 344284 355456
rect 344336 355444 344342 355496
rect 58802 355376 58808 355428
rect 58860 355416 58866 355428
rect 355410 355416 355416 355428
rect 58860 355388 355416 355416
rect 58860 355376 58866 355388
rect 355410 355376 355416 355388
rect 355468 355376 355474 355428
rect 452654 355376 452660 355428
rect 452712 355416 452718 355428
rect 474642 355416 474648 355428
rect 452712 355388 474648 355416
rect 452712 355376 452718 355388
rect 474642 355376 474648 355388
rect 474700 355376 474706 355428
rect 237742 355308 237748 355360
rect 237800 355348 237806 355360
rect 536098 355348 536104 355360
rect 237800 355320 536104 355348
rect 237800 355308 237806 355320
rect 536098 355308 536104 355320
rect 536156 355308 536162 355360
rect 240042 354628 240048 354680
rect 240100 354668 240106 354680
rect 580442 354668 580448 354680
rect 240100 354640 580448 354668
rect 240100 354628 240106 354640
rect 580442 354628 580448 354640
rect 580500 354628 580506 354680
rect 237834 353948 237840 354000
rect 237892 353988 237898 354000
rect 452654 353988 452660 354000
rect 237892 353960 452660 353988
rect 237892 353948 237898 353960
rect 452654 353948 452660 353960
rect 452712 353948 452718 354000
rect 239398 353404 239404 353456
rect 239456 353444 239462 353456
rect 296806 353444 296812 353456
rect 239456 353416 296812 353444
rect 239456 353404 239462 353416
rect 296806 353404 296812 353416
rect 296864 353404 296870 353456
rect 237098 353336 237104 353388
rect 237156 353376 237162 353388
rect 295334 353376 295340 353388
rect 237156 353348 295340 353376
rect 237156 353336 237162 353348
rect 295334 353336 295340 353348
rect 295392 353336 295398 353388
rect 237006 353268 237012 353320
rect 237064 353308 237070 353320
rect 296714 353308 296720 353320
rect 237064 353280 296720 353308
rect 237064 353268 237070 353280
rect 296714 353268 296720 353280
rect 296772 353268 296778 353320
rect 240042 353200 240048 353252
rect 240100 353240 240106 353252
rect 402238 353240 402244 353252
rect 240100 353212 402244 353240
rect 240100 353200 240106 353212
rect 402238 353200 402244 353212
rect 402296 353200 402302 353252
rect 531222 353200 531228 353252
rect 531280 353240 531286 353252
rect 580166 353240 580172 353252
rect 531280 353212 580172 353240
rect 531280 353200 531286 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 282086 353132 282092 353184
rect 282144 353172 282150 353184
rect 539594 353172 539600 353184
rect 282144 353144 539600 353172
rect 282144 353132 282150 353144
rect 539594 353132 539600 353144
rect 539652 353132 539658 353184
rect 60550 353064 60556 353116
rect 60608 353104 60614 353116
rect 350074 353104 350080 353116
rect 60608 353076 350080 353104
rect 60608 353064 60614 353076
rect 350074 353064 350080 353076
rect 350132 353064 350138 353116
rect 52730 352996 52736 353048
rect 52788 353036 52794 353048
rect 347498 353036 347504 353048
rect 52788 353008 347504 353036
rect 52788 352996 52794 353008
rect 347498 352996 347504 353008
rect 347556 352996 347562 353048
rect 52362 352928 52368 352980
rect 52420 352968 52426 352980
rect 347406 352968 347412 352980
rect 52420 352940 347412 352968
rect 52420 352928 52426 352940
rect 347406 352928 347412 352940
rect 347464 352928 347470 352980
rect 56134 352860 56140 352912
rect 56192 352900 56198 352912
rect 352650 352900 352656 352912
rect 56192 352872 352656 352900
rect 56192 352860 56198 352872
rect 352650 352860 352656 352872
rect 352708 352860 352714 352912
rect 54478 352792 54484 352844
rect 54536 352832 54542 352844
rect 352742 352832 352748 352844
rect 54536 352804 352748 352832
rect 54536 352792 54542 352804
rect 352742 352792 352748 352804
rect 352800 352792 352806 352844
rect 46474 352724 46480 352776
rect 46532 352764 46538 352776
rect 349982 352764 349988 352776
rect 46532 352736 349988 352764
rect 46532 352724 46538 352736
rect 349982 352724 349988 352736
rect 350040 352724 350046 352776
rect 46750 352656 46756 352708
rect 46808 352696 46814 352708
rect 352558 352696 352564 352708
rect 46808 352668 352564 352696
rect 46808 352656 46814 352668
rect 352558 352656 352564 352668
rect 352616 352656 352622 352708
rect 28626 352588 28632 352640
rect 28684 352628 28690 352640
rect 355502 352628 355508 352640
rect 28684 352600 355508 352628
rect 28684 352588 28690 352600
rect 355502 352588 355508 352600
rect 355560 352588 355566 352640
rect 27338 352520 27344 352572
rect 27396 352560 27402 352572
rect 355594 352560 355600 352572
rect 27396 352532 355600 352560
rect 27396 352520 27402 352532
rect 355594 352520 355600 352532
rect 355652 352520 355658 352572
rect 235350 351908 235356 351960
rect 235408 351948 235414 351960
rect 288434 351948 288440 351960
rect 235408 351920 288440 351948
rect 235408 351908 235414 351920
rect 288434 351908 288440 351920
rect 288492 351908 288498 351960
rect 234982 351772 234988 351824
rect 235040 351812 235046 351824
rect 235350 351812 235356 351824
rect 235040 351784 235356 351812
rect 235040 351772 235046 351784
rect 235350 351772 235356 351784
rect 235408 351772 235414 351824
rect 359918 351432 359924 351484
rect 359976 351472 359982 351484
rect 503254 351472 503260 351484
rect 359976 351444 503260 351472
rect 359976 351432 359982 351444
rect 503254 351432 503260 351444
rect 503312 351432 503318 351484
rect 281994 351364 282000 351416
rect 282052 351404 282058 351416
rect 541158 351404 541164 351416
rect 282052 351376 541164 351404
rect 282052 351364 282058 351376
rect 541158 351364 541164 351376
rect 541216 351364 541222 351416
rect 239582 351296 239588 351348
rect 239640 351336 239646 351348
rect 510062 351336 510068 351348
rect 239640 351308 510068 351336
rect 239640 351296 239646 351308
rect 510062 351296 510068 351308
rect 510120 351296 510126 351348
rect 239858 351228 239864 351280
rect 239916 351268 239922 351280
rect 580258 351268 580264 351280
rect 239916 351240 580264 351268
rect 239916 351228 239922 351240
rect 580258 351228 580264 351240
rect 580316 351228 580322 351280
rect 43254 351160 43260 351212
rect 43312 351200 43318 351212
rect 503714 351200 503720 351212
rect 43312 351172 503720 351200
rect 43312 351160 43318 351172
rect 503714 351160 503720 351172
rect 503772 351160 503778 351212
rect 229922 351092 229928 351144
rect 229980 351132 229986 351144
rect 280246 351132 280252 351144
rect 229980 351104 280252 351132
rect 229980 351092 229986 351104
rect 280246 351092 280252 351104
rect 280304 351092 280310 351144
rect 230290 351024 230296 351076
rect 230348 351064 230354 351076
rect 283006 351064 283012 351076
rect 230348 351036 283012 351064
rect 230348 351024 230354 351036
rect 283006 351024 283012 351036
rect 283064 351024 283070 351076
rect 224678 350956 224684 351008
rect 224736 350996 224742 351008
rect 280338 350996 280344 351008
rect 224736 350968 280344 350996
rect 224736 350956 224742 350968
rect 280338 350956 280344 350968
rect 280396 350956 280402 351008
rect 221458 350888 221464 350940
rect 221516 350928 221522 350940
rect 277946 350928 277952 350940
rect 221516 350900 277952 350928
rect 221516 350888 221522 350900
rect 277946 350888 277952 350900
rect 278004 350888 278010 350940
rect 224218 350820 224224 350872
rect 224276 350860 224282 350872
rect 290550 350860 290556 350872
rect 224276 350832 290556 350860
rect 224276 350820 224282 350832
rect 290550 350820 290556 350832
rect 290608 350820 290614 350872
rect 217410 350752 217416 350804
rect 217468 350792 217474 350804
rect 288710 350792 288716 350804
rect 217468 350764 288716 350792
rect 217468 350752 217474 350764
rect 288710 350752 288716 350764
rect 288768 350752 288774 350804
rect 217318 350684 217324 350736
rect 217376 350724 217382 350736
rect 291562 350724 291568 350736
rect 217376 350696 291568 350724
rect 217376 350684 217382 350696
rect 291562 350684 291568 350696
rect 291620 350684 291626 350736
rect 237926 350616 237932 350668
rect 237984 350656 237990 350668
rect 318058 350656 318064 350668
rect 237984 350628 318064 350656
rect 237984 350616 237990 350628
rect 318058 350616 318064 350628
rect 318116 350616 318122 350668
rect 222102 350548 222108 350600
rect 222160 350588 222166 350600
rect 311250 350588 311256 350600
rect 222160 350560 311256 350588
rect 222160 350548 222166 350560
rect 311250 350548 311256 350560
rect 311308 350548 311314 350600
rect 232498 350480 232504 350532
rect 232556 350520 232562 350532
rect 240042 350520 240048 350532
rect 232556 350492 240048 350520
rect 232556 350480 232562 350492
rect 240042 350480 240048 350492
rect 240100 350480 240106 350532
rect 226334 350344 226340 350396
rect 226392 350384 226398 350396
rect 298094 350384 298100 350396
rect 226392 350356 298100 350384
rect 226392 350344 226398 350356
rect 298094 350344 298100 350356
rect 298152 350344 298158 350396
rect 282730 350276 282736 350328
rect 282788 350316 282794 350328
rect 539778 350316 539784 350328
rect 282788 350288 539784 350316
rect 282788 350276 282794 350288
rect 539778 350276 539784 350288
rect 539836 350276 539842 350328
rect 50798 350208 50804 350260
rect 50856 350248 50862 350260
rect 336458 350248 336464 350260
rect 50856 350220 336464 350248
rect 50856 350208 50862 350220
rect 336458 350208 336464 350220
rect 336516 350208 336522 350260
rect 55858 350140 55864 350192
rect 55916 350180 55922 350192
rect 344462 350180 344468 350192
rect 55916 350152 344468 350180
rect 55916 350140 55922 350152
rect 344462 350140 344468 350152
rect 344520 350140 344526 350192
rect 42610 350072 42616 350124
rect 42668 350112 42674 350124
rect 339034 350112 339040 350124
rect 42668 350084 339040 350112
rect 42668 350072 42674 350084
rect 339034 350072 339040 350084
rect 339092 350072 339098 350124
rect 43806 350004 43812 350056
rect 43864 350044 43870 350056
rect 352834 350044 352840 350056
rect 43864 350016 352840 350044
rect 43864 350004 43870 350016
rect 352834 350004 352840 350016
rect 352892 350004 352898 350056
rect 48774 349936 48780 349988
rect 48832 349976 48838 349988
rect 359642 349976 359648 349988
rect 48832 349948 359648 349976
rect 48832 349936 48838 349948
rect 359642 349936 359648 349948
rect 359700 349936 359706 349988
rect 43898 349868 43904 349920
rect 43956 349908 43962 349920
rect 501230 349908 501236 349920
rect 43956 349880 501236 349908
rect 43956 349868 43962 349880
rect 501230 349868 501236 349880
rect 501288 349868 501294 349920
rect 41138 349800 41144 349852
rect 41196 349840 41202 349852
rect 502610 349840 502616 349852
rect 41196 349812 502616 349840
rect 41196 349800 41202 349812
rect 502610 349800 502616 349812
rect 502668 349800 502674 349852
rect 153838 349732 153844 349784
rect 153896 349772 153902 349784
rect 158714 349772 158720 349784
rect 153896 349744 158720 349772
rect 153896 349732 153902 349744
rect 158714 349732 158720 349744
rect 158772 349732 158778 349784
rect 254578 349324 254584 349376
rect 254636 349364 254642 349376
rect 292574 349364 292580 349376
rect 254636 349336 292580 349364
rect 254636 349324 254642 349336
rect 292574 349324 292580 349336
rect 292632 349324 292638 349376
rect 234982 349256 234988 349308
rect 235040 349296 235046 349308
rect 580258 349296 580264 349308
rect 235040 349268 580264 349296
rect 235040 349256 235046 349268
rect 580258 349256 580264 349268
rect 580316 349256 580322 349308
rect 220170 349188 220176 349240
rect 220228 349228 220234 349240
rect 283374 349228 283380 349240
rect 220228 349200 283380 349228
rect 220228 349188 220234 349200
rect 283374 349188 283380 349200
rect 283432 349188 283438 349240
rect 221642 349120 221648 349172
rect 221700 349160 221706 349172
rect 302326 349160 302332 349172
rect 221700 349132 302332 349160
rect 221700 349120 221706 349132
rect 302326 349120 302332 349132
rect 302384 349120 302390 349172
rect 259362 348576 259368 348628
rect 259420 348616 259426 348628
rect 302510 348616 302516 348628
rect 259420 348588 302516 348616
rect 259420 348576 259426 348588
rect 302510 348576 302516 348588
rect 302568 348576 302574 348628
rect 233970 348508 233976 348560
rect 234028 348548 234034 348560
rect 282914 348548 282920 348560
rect 234028 348520 282920 348548
rect 234028 348508 234034 348520
rect 282914 348508 282920 348520
rect 282972 348508 282978 348560
rect 226518 348440 226524 348492
rect 226576 348480 226582 348492
rect 278038 348480 278044 348492
rect 226576 348452 278044 348480
rect 226576 348440 226582 348452
rect 278038 348440 278044 348452
rect 278096 348440 278102 348492
rect 212258 348372 212264 348424
rect 212316 348412 212322 348424
rect 312538 348412 312544 348424
rect 212316 348384 312544 348412
rect 212316 348372 212322 348384
rect 312538 348372 312544 348384
rect 312596 348372 312602 348424
rect 249702 348304 249708 348356
rect 249760 348344 249766 348356
rect 301038 348344 301044 348356
rect 249760 348316 301044 348344
rect 249760 348304 249766 348316
rect 301038 348304 301044 348316
rect 301096 348304 301102 348356
rect 232682 348236 232688 348288
rect 232740 348276 232746 348288
rect 284294 348276 284300 348288
rect 232740 348248 284300 348276
rect 232740 348236 232746 348248
rect 284294 348236 284300 348248
rect 284352 348236 284358 348288
rect 226426 348168 226432 348220
rect 226484 348208 226490 348220
rect 290642 348208 290648 348220
rect 226484 348180 290648 348208
rect 226484 348168 226490 348180
rect 290642 348168 290648 348180
rect 290700 348168 290706 348220
rect 226334 348100 226340 348152
rect 226392 348140 226398 348152
rect 299566 348140 299572 348152
rect 226392 348112 299572 348140
rect 226392 348100 226398 348112
rect 299566 348100 299572 348112
rect 299624 348100 299630 348152
rect 222102 348032 222108 348084
rect 222160 348072 222166 348084
rect 296070 348072 296076 348084
rect 222160 348044 296076 348072
rect 222160 348032 222166 348044
rect 296070 348032 296076 348044
rect 296128 348032 296134 348084
rect 212442 347964 212448 348016
rect 212500 348004 212506 348016
rect 287790 348004 287796 348016
rect 212500 347976 287796 348004
rect 212500 347964 212506 347976
rect 287790 347964 287796 347976
rect 287848 347964 287854 348016
rect 220722 347896 220728 347948
rect 220780 347936 220786 347948
rect 298830 347936 298836 347948
rect 220780 347908 298836 347936
rect 220780 347896 220786 347908
rect 298830 347896 298836 347908
rect 298888 347896 298894 347948
rect 211982 347828 211988 347880
rect 212040 347868 212046 347880
rect 292850 347868 292856 347880
rect 212040 347840 292856 347868
rect 212040 347828 212046 347840
rect 292850 347828 292856 347840
rect 292908 347828 292914 347880
rect 224218 347760 224224 347812
rect 224276 347800 224282 347812
rect 322290 347800 322296 347812
rect 224276 347772 322296 347800
rect 224276 347760 224282 347772
rect 322290 347760 322296 347772
rect 322348 347760 322354 347812
rect 60642 347216 60648 347268
rect 60700 347256 60706 347268
rect 350258 347256 350264 347268
rect 60700 347228 350264 347256
rect 60700 347216 60706 347228
rect 350258 347216 350264 347228
rect 350316 347216 350322 347268
rect 50614 347148 50620 347200
rect 50672 347188 50678 347200
rect 344554 347188 344560 347200
rect 50672 347160 344560 347188
rect 50672 347148 50678 347160
rect 344554 347148 344560 347160
rect 344612 347148 344618 347200
rect 47946 347080 47952 347132
rect 48004 347120 48010 347132
rect 350166 347120 350172 347132
rect 48004 347092 350172 347120
rect 48004 347080 48010 347092
rect 350166 347080 350172 347092
rect 350224 347080 350230 347132
rect 31478 347012 31484 347064
rect 31536 347052 31542 347064
rect 358170 347052 358176 347064
rect 31536 347024 358176 347052
rect 31536 347012 31542 347024
rect 358170 347012 358176 347024
rect 358228 347012 358234 347064
rect 266354 346944 266360 346996
rect 266412 346984 266418 346996
rect 285766 346984 285772 346996
rect 266412 346956 285772 346984
rect 266412 346944 266418 346956
rect 285766 346944 285772 346956
rect 285824 346944 285830 346996
rect 273254 346876 273260 346928
rect 273312 346916 273318 346928
rect 298278 346916 298284 346928
rect 273312 346888 298284 346916
rect 273312 346876 273318 346888
rect 298278 346876 298284 346888
rect 298336 346876 298342 346928
rect 243538 346808 243544 346860
rect 243596 346848 243602 346860
rect 283190 346848 283196 346860
rect 243596 346820 283196 346848
rect 243596 346808 243602 346820
rect 283190 346808 283196 346820
rect 283248 346808 283254 346860
rect 226058 346740 226064 346792
rect 226116 346780 226122 346792
rect 280522 346780 280528 346792
rect 226116 346752 280528 346780
rect 226116 346740 226122 346752
rect 280522 346740 280528 346752
rect 280580 346740 280586 346792
rect 224218 346672 224224 346724
rect 224276 346712 224282 346724
rect 291194 346712 291200 346724
rect 224276 346684 291200 346712
rect 224276 346672 224282 346684
rect 291194 346672 291200 346684
rect 291252 346672 291258 346724
rect 220722 346604 220728 346656
rect 220780 346644 220786 346656
rect 289262 346644 289268 346656
rect 220780 346616 289268 346644
rect 220780 346604 220786 346616
rect 289262 346604 289268 346616
rect 289320 346604 289326 346656
rect 223298 346536 223304 346588
rect 223356 346576 223362 346588
rect 303062 346576 303068 346588
rect 223356 346548 303068 346576
rect 223356 346536 223362 346548
rect 303062 346536 303068 346548
rect 303120 346536 303126 346588
rect 225046 346468 225052 346520
rect 225104 346508 225110 346520
rect 314102 346508 314108 346520
rect 225104 346480 314108 346508
rect 225104 346468 225110 346480
rect 314102 346468 314108 346480
rect 314160 346468 314166 346520
rect 224954 346400 224960 346452
rect 225012 346440 225018 346452
rect 325050 346440 325056 346452
rect 225012 346412 325056 346440
rect 225012 346400 225018 346412
rect 325050 346400 325056 346412
rect 325108 346400 325114 346452
rect 260742 346332 260748 346384
rect 260800 346372 260806 346384
rect 360378 346372 360384 346384
rect 260800 346344 360384 346372
rect 260800 346332 260806 346344
rect 360378 346332 360384 346344
rect 360436 346332 360442 346384
rect 503622 346332 503628 346384
rect 503680 346372 503686 346384
rect 523402 346372 523408 346384
rect 503680 346344 523408 346372
rect 503680 346332 503686 346344
rect 523402 346332 523408 346344
rect 523460 346332 523466 346384
rect 253106 346264 253112 346316
rect 253164 346304 253170 346316
rect 273254 346304 273260 346316
rect 253164 346276 273260 346304
rect 253164 346264 253170 346276
rect 273254 346264 273260 346276
rect 273312 346264 273318 346316
rect 229738 345856 229744 345908
rect 229796 345896 229802 345908
rect 280154 345896 280160 345908
rect 229796 345868 280160 345896
rect 229796 345856 229802 345868
rect 280154 345856 280160 345868
rect 280212 345856 280218 345908
rect 227714 345788 227720 345840
rect 227772 345828 227778 345840
rect 278958 345828 278964 345840
rect 227772 345800 278964 345828
rect 227772 345788 227778 345800
rect 278958 345788 278964 345800
rect 279016 345788 279022 345840
rect 225874 345720 225880 345772
rect 225932 345760 225938 345772
rect 284294 345760 284300 345772
rect 225932 345732 284300 345760
rect 225932 345720 225938 345732
rect 284294 345720 284300 345732
rect 284352 345720 284358 345772
rect 216674 345652 216680 345704
rect 216732 345692 216738 345704
rect 304350 345692 304356 345704
rect 216732 345664 304356 345692
rect 216732 345652 216738 345664
rect 304350 345652 304356 345664
rect 304408 345652 304414 345704
rect 274634 345584 274640 345636
rect 274692 345624 274698 345636
rect 295518 345624 295524 345636
rect 274692 345596 295524 345624
rect 274692 345584 274698 345596
rect 295518 345584 295524 345596
rect 295576 345584 295582 345636
rect 244274 345516 244280 345568
rect 244332 345556 244338 345568
rect 298186 345556 298192 345568
rect 244332 345528 298192 345556
rect 244332 345516 244338 345528
rect 298186 345516 298192 345528
rect 298244 345516 298250 345568
rect 223206 345448 223212 345500
rect 223264 345488 223270 345500
rect 289354 345488 289360 345500
rect 223264 345460 289360 345488
rect 223264 345448 223270 345460
rect 289354 345448 289360 345460
rect 289412 345448 289418 345500
rect 228358 345380 228364 345432
rect 228416 345420 228422 345432
rect 299474 345420 299480 345432
rect 228416 345392 299480 345420
rect 228416 345380 228422 345392
rect 299474 345380 299480 345392
rect 299532 345380 299538 345432
rect 158714 345312 158720 345364
rect 158772 345352 158778 345364
rect 161566 345352 161572 345364
rect 158772 345324 161572 345352
rect 158772 345312 158778 345324
rect 161566 345312 161572 345324
rect 161624 345312 161630 345364
rect 226334 345312 226340 345364
rect 226392 345352 226398 345364
rect 307294 345352 307300 345364
rect 226392 345324 307300 345352
rect 226392 345312 226398 345324
rect 307294 345312 307300 345324
rect 307352 345312 307358 345364
rect 223298 345244 223304 345296
rect 223356 345284 223362 345296
rect 305822 345284 305828 345296
rect 223356 345256 305828 345284
rect 223356 345244 223362 345256
rect 305822 345244 305828 345256
rect 305880 345244 305886 345296
rect 209130 345176 209136 345228
rect 209188 345216 209194 345228
rect 296898 345216 296904 345228
rect 209188 345188 296904 345216
rect 209188 345176 209194 345188
rect 296898 345176 296904 345188
rect 296956 345176 296962 345228
rect 223114 345108 223120 345160
rect 223172 345148 223178 345160
rect 327718 345148 327724 345160
rect 223172 345120 327724 345148
rect 223172 345108 223178 345120
rect 327718 345108 327724 345120
rect 327776 345108 327782 345160
rect 220722 345040 220728 345092
rect 220780 345080 220786 345092
rect 334618 345080 334624 345092
rect 220780 345052 334624 345080
rect 220780 345040 220786 345052
rect 334618 345040 334624 345052
rect 334676 345040 334682 345092
rect 243538 344972 243544 345024
rect 243596 345012 243602 345024
rect 360286 345012 360292 345024
rect 243596 344984 360292 345012
rect 243596 344972 243602 344984
rect 360286 344972 360292 344984
rect 360344 344972 360350 345024
rect 228450 344360 228456 344412
rect 228508 344400 228514 344412
rect 254578 344400 254584 344412
rect 228508 344372 254584 344400
rect 228508 344360 228514 344372
rect 254578 344360 254584 344372
rect 254636 344360 254642 344412
rect 271782 344360 271788 344412
rect 271840 344400 271846 344412
rect 287238 344400 287244 344412
rect 271840 344372 287244 344400
rect 271840 344360 271846 344372
rect 287238 344360 287244 344372
rect 287296 344360 287302 344412
rect 251082 344292 251088 344344
rect 251140 344332 251146 344344
rect 279326 344332 279332 344344
rect 251140 344304 279332 344332
rect 251140 344292 251146 344304
rect 279326 344292 279332 344304
rect 279384 344292 279390 344344
rect 293586 344292 293592 344344
rect 293644 344332 293650 344344
rect 304534 344332 304540 344344
rect 293644 344304 304540 344332
rect 293644 344292 293650 344304
rect 304534 344292 304540 344304
rect 304592 344292 304598 344344
rect 255314 344224 255320 344276
rect 255372 344264 255378 344276
rect 292758 344264 292764 344276
rect 255372 344236 292764 344264
rect 255372 344224 255378 344236
rect 292758 344224 292764 344236
rect 292816 344224 292822 344276
rect 235994 344156 236000 344208
rect 236052 344196 236058 344208
rect 285030 344196 285036 344208
rect 236052 344168 285036 344196
rect 236052 344156 236058 344168
rect 285030 344156 285036 344168
rect 285088 344156 285094 344208
rect 218054 344088 218060 344140
rect 218112 344128 218118 344140
rect 293310 344128 293316 344140
rect 218112 344100 293316 344128
rect 218112 344088 218118 344100
rect 293310 344088 293316 344100
rect 293368 344088 293374 344140
rect 231118 344020 231124 344072
rect 231176 344060 231182 344072
rect 316678 344060 316684 344072
rect 231176 344032 316684 344060
rect 231176 344020 231182 344032
rect 316678 344020 316684 344032
rect 316736 344020 316742 344072
rect 216674 343952 216680 344004
rect 216732 343992 216738 344004
rect 307110 343992 307116 344004
rect 216732 343964 307116 343992
rect 216732 343952 216738 343964
rect 307110 343952 307116 343964
rect 307168 343952 307174 344004
rect 228266 343884 228272 343936
rect 228324 343924 228330 343936
rect 319438 343924 319444 343936
rect 228324 343896 319444 343924
rect 228324 343884 228330 343896
rect 319438 343884 319444 343896
rect 319496 343884 319502 343936
rect 224218 343816 224224 343868
rect 224276 343856 224282 343868
rect 319530 343856 319536 343868
rect 224276 343828 319536 343856
rect 224276 343816 224282 343828
rect 319530 343816 319536 343828
rect 319588 343816 319594 343868
rect 214558 343748 214564 343800
rect 214616 343788 214622 343800
rect 314010 343788 314016 343800
rect 214616 343760 314016 343788
rect 214616 343748 214622 343760
rect 314010 343748 314016 343760
rect 314068 343748 314074 343800
rect 125502 343680 125508 343732
rect 125560 343720 125566 343732
rect 322198 343720 322204 343732
rect 125560 343692 322204 343720
rect 125560 343680 125566 343692
rect 322198 343680 322204 343692
rect 322256 343680 322262 343732
rect 61930 343612 61936 343664
rect 61988 343652 61994 343664
rect 302878 343652 302884 343664
rect 61988 343624 302884 343652
rect 61988 343612 61994 343624
rect 302878 343612 302884 343624
rect 302936 343612 302942 343664
rect 231118 343204 231124 343256
rect 231176 343244 231182 343256
rect 280706 343244 280712 343256
rect 231176 343216 280712 343244
rect 231176 343204 231182 343216
rect 280706 343204 280712 343216
rect 280764 343204 280770 343256
rect 276106 343136 276112 343188
rect 276164 343176 276170 343188
rect 358354 343176 358360 343188
rect 276164 343148 358360 343176
rect 276164 343136 276170 343148
rect 358354 343136 358360 343148
rect 358412 343136 358418 343188
rect 262306 343068 262312 343120
rect 262364 343108 262370 343120
rect 356698 343108 356704 343120
rect 262364 343080 356704 343108
rect 262364 343068 262370 343080
rect 356698 343068 356704 343080
rect 356756 343068 356762 343120
rect 250346 343000 250352 343052
rect 250404 343040 250410 343052
rect 253198 343040 253204 343052
rect 250404 343012 253204 343040
rect 250404 343000 250410 343012
rect 253198 343000 253204 343012
rect 253256 343000 253262 343052
rect 253474 343000 253480 343052
rect 253532 343040 253538 343052
rect 359366 343040 359372 343052
rect 253532 343012 359372 343040
rect 253532 343000 253538 343012
rect 359366 343000 359372 343012
rect 359424 343000 359430 343052
rect 161566 342932 161572 342984
rect 161624 342972 161630 342984
rect 176654 342972 176660 342984
rect 161624 342944 176660 342972
rect 161624 342932 161630 342944
rect 176654 342932 176660 342944
rect 176712 342932 176718 342984
rect 239214 342932 239220 342984
rect 239272 342972 239278 342984
rect 358538 342972 358544 342984
rect 239272 342944 358544 342972
rect 239272 342932 239278 342944
rect 358538 342932 358544 342944
rect 358596 342932 358602 342984
rect 59998 342864 60004 342916
rect 60056 342904 60062 342916
rect 350350 342904 350356 342916
rect 60056 342876 350356 342904
rect 60056 342864 60062 342876
rect 350350 342864 350356 342876
rect 350408 342864 350414 342916
rect 221734 342796 221740 342848
rect 221792 342836 221798 342848
rect 276014 342836 276020 342848
rect 221792 342808 276020 342836
rect 221792 342796 221798 342808
rect 276014 342796 276020 342808
rect 276072 342796 276078 342848
rect 224218 342728 224224 342780
rect 224276 342768 224282 342780
rect 282914 342768 282920 342780
rect 224276 342740 282920 342768
rect 224276 342728 224282 342740
rect 282914 342728 282920 342740
rect 282972 342728 282978 342780
rect 209222 342660 209228 342712
rect 209280 342700 209286 342712
rect 279418 342700 279424 342712
rect 209280 342672 279424 342700
rect 209280 342660 209286 342672
rect 279418 342660 279424 342672
rect 279476 342660 279482 342712
rect 214558 342592 214564 342644
rect 214616 342632 214622 342644
rect 286594 342632 286600 342644
rect 214616 342604 286600 342632
rect 214616 342592 214622 342604
rect 286594 342592 286600 342604
rect 286652 342592 286658 342644
rect 214466 342524 214472 342576
rect 214524 342564 214530 342576
rect 287974 342564 287980 342576
rect 214524 342536 287980 342564
rect 214524 342524 214530 342536
rect 287974 342524 287980 342536
rect 288032 342524 288038 342576
rect 220354 342456 220360 342508
rect 220412 342496 220418 342508
rect 305638 342496 305644 342508
rect 220412 342468 305644 342496
rect 220412 342456 220418 342468
rect 305638 342456 305644 342468
rect 305696 342496 305702 342508
rect 306098 342496 306104 342508
rect 305696 342468 306104 342496
rect 305696 342456 305702 342468
rect 306098 342456 306104 342468
rect 306156 342456 306162 342508
rect 244274 342388 244280 342440
rect 244332 342428 244338 342440
rect 339218 342428 339224 342440
rect 244332 342400 339224 342428
rect 244332 342388 244338 342400
rect 339218 342388 339224 342400
rect 339276 342388 339282 342440
rect 214650 342320 214656 342372
rect 214708 342360 214714 342372
rect 311342 342360 311348 342372
rect 214708 342332 311348 342360
rect 214708 342320 214714 342332
rect 311342 342320 311348 342332
rect 311400 342320 311406 342372
rect 214374 342252 214380 342304
rect 214432 342292 214438 342304
rect 320818 342292 320824 342304
rect 214432 342264 320824 342292
rect 214432 342252 214438 342264
rect 320818 342252 320824 342264
rect 320876 342252 320882 342304
rect 240042 342184 240048 342236
rect 240100 342224 240106 342236
rect 356790 342224 356796 342236
rect 240100 342196 356796 342224
rect 240100 342184 240106 342196
rect 356790 342184 356796 342196
rect 356848 342184 356854 342236
rect 270402 341708 270408 341760
rect 270460 341748 270466 341760
rect 295702 341748 295708 341760
rect 270460 341720 295708 341748
rect 270460 341708 270466 341720
rect 295702 341708 295708 341720
rect 295760 341708 295766 341760
rect 256694 341640 256700 341692
rect 256752 341680 256758 341692
rect 285858 341680 285864 341692
rect 256752 341652 285864 341680
rect 256752 341640 256758 341652
rect 285858 341640 285864 341652
rect 285916 341640 285922 341692
rect 231118 341572 231124 341624
rect 231176 341612 231182 341624
rect 280614 341612 280620 341624
rect 231176 341584 280620 341612
rect 231176 341572 231182 341584
rect 280614 341572 280620 341584
rect 280672 341572 280678 341624
rect 216674 341504 216680 341556
rect 216732 341544 216738 341556
rect 285674 341544 285680 341556
rect 216732 341516 285680 341544
rect 216732 341504 216738 341516
rect 285674 341504 285680 341516
rect 285732 341504 285738 341556
rect 224954 341436 224960 341488
rect 225012 341476 225018 341488
rect 300394 341476 300400 341488
rect 225012 341448 300400 341476
rect 225012 341436 225018 341448
rect 300394 341436 300400 341448
rect 300452 341436 300458 341488
rect 228542 341368 228548 341420
rect 228600 341408 228606 341420
rect 323578 341408 323584 341420
rect 228600 341380 323584 341408
rect 228600 341368 228606 341380
rect 323578 341368 323584 341380
rect 323636 341368 323642 341420
rect 223298 341300 223304 341352
rect 223356 341340 223362 341352
rect 321002 341340 321008 341352
rect 223356 341312 321008 341340
rect 223356 341300 223362 341312
rect 321002 341300 321008 341312
rect 321060 341300 321066 341352
rect 235994 341232 236000 341284
rect 236052 341272 236058 341284
rect 342898 341272 342904 341284
rect 236052 341244 342904 341272
rect 236052 341232 236058 341244
rect 342898 341232 342904 341244
rect 342956 341232 342962 341284
rect 220722 341164 220728 341216
rect 220780 341204 220786 341216
rect 336550 341204 336556 341216
rect 220780 341176 336556 341204
rect 220780 341164 220786 341176
rect 336550 341164 336556 341176
rect 336608 341164 336614 341216
rect 68922 341096 68928 341148
rect 68980 341136 68986 341148
rect 311158 341136 311164 341148
rect 68980 341108 311164 341136
rect 68980 341096 68986 341108
rect 311158 341096 311164 341108
rect 311216 341096 311222 341148
rect 66070 341028 66076 341080
rect 66128 341068 66134 341080
rect 307846 341068 307852 341080
rect 66128 341040 307852 341068
rect 66128 341028 66134 341040
rect 307846 341028 307852 341040
rect 307904 341068 307910 341080
rect 308398 341068 308404 341080
rect 307904 341040 308404 341068
rect 307904 341028 307910 341040
rect 308398 341028 308404 341040
rect 308456 341028 308462 341080
rect 66162 340960 66168 341012
rect 66220 341000 66226 341012
rect 309778 341000 309784 341012
rect 66220 340972 309784 341000
rect 66220 340960 66226 340972
rect 309778 340960 309784 340972
rect 309836 340960 309842 341012
rect 71590 340892 71596 340944
rect 71648 340932 71654 340944
rect 315298 340932 315304 340944
rect 71648 340904 315304 340932
rect 71648 340892 71654 340904
rect 315298 340892 315304 340904
rect 315356 340892 315362 340944
rect 216674 340824 216680 340876
rect 216732 340864 216738 340876
rect 348418 340864 348424 340876
rect 216732 340836 348424 340864
rect 216732 340824 216738 340836
rect 348418 340824 348424 340836
rect 348476 340824 348482 340876
rect 503622 340824 503628 340876
rect 503680 340864 503686 340876
rect 520642 340864 520648 340876
rect 503680 340836 520648 340864
rect 503680 340824 503686 340836
rect 520642 340824 520648 340836
rect 520700 340824 520706 340876
rect 216858 340756 216864 340808
rect 216916 340796 216922 340808
rect 342806 340796 342812 340808
rect 216916 340768 342812 340796
rect 216916 340756 216922 340768
rect 342806 340756 342812 340768
rect 342864 340756 342870 340808
rect 278038 340416 278044 340468
rect 278096 340456 278102 340468
rect 303706 340456 303712 340468
rect 278096 340428 303712 340456
rect 278096 340416 278102 340428
rect 303706 340416 303712 340428
rect 303764 340416 303770 340468
rect 276014 340348 276020 340400
rect 276072 340388 276078 340400
rect 302418 340388 302424 340400
rect 276072 340360 302424 340388
rect 276072 340348 276078 340360
rect 302418 340348 302424 340360
rect 302476 340348 302482 340400
rect 236914 340280 236920 340332
rect 236972 340320 236978 340332
rect 355042 340320 355048 340332
rect 236972 340292 355048 340320
rect 236972 340280 236978 340292
rect 355042 340280 355048 340292
rect 355100 340280 355106 340332
rect 238386 340212 238392 340264
rect 238444 340252 238450 340264
rect 359734 340252 359740 340264
rect 238444 340224 359740 340252
rect 238444 340212 238450 340224
rect 359734 340212 359740 340224
rect 359792 340212 359798 340264
rect 103422 340144 103428 340196
rect 103480 340184 103486 340196
rect 346302 340184 346308 340196
rect 103480 340156 346308 340184
rect 103480 340144 103486 340156
rect 346302 340144 346308 340156
rect 346360 340144 346366 340196
rect 279050 340076 279056 340128
rect 279108 340116 279114 340128
rect 281350 340116 281356 340128
rect 279108 340088 281356 340116
rect 279108 340076 279114 340088
rect 281350 340076 281356 340088
rect 281408 340076 281414 340128
rect 242434 340008 242440 340060
rect 242492 340048 242498 340060
rect 275738 340048 275744 340060
rect 242492 340020 275744 340048
rect 242492 340008 242498 340020
rect 275738 340008 275744 340020
rect 275796 340008 275802 340060
rect 280062 340008 280068 340060
rect 280120 340048 280126 340060
rect 281166 340048 281172 340060
rect 280120 340020 281172 340048
rect 280120 340008 280126 340020
rect 281166 340008 281172 340020
rect 281224 340008 281230 340060
rect 241422 339940 241428 339992
rect 241480 339980 241486 339992
rect 250990 339980 250996 339992
rect 241480 339952 250996 339980
rect 241480 339940 241486 339952
rect 250990 339940 250996 339952
rect 251048 339940 251054 339992
rect 279786 339940 279792 339992
rect 279844 339980 279850 339992
rect 281258 339980 281264 339992
rect 279844 339952 281264 339980
rect 279844 339940 279850 339952
rect 281258 339940 281264 339952
rect 281316 339940 281322 339992
rect 250898 339872 250904 339924
rect 250956 339912 250962 339924
rect 300946 339912 300952 339924
rect 250956 339884 300952 339912
rect 250956 339872 250962 339884
rect 300946 339872 300952 339884
rect 301004 339872 301010 339924
rect 229922 339804 229928 339856
rect 229980 339844 229986 339856
rect 289538 339844 289544 339856
rect 229980 339816 289544 339844
rect 229980 339804 229986 339816
rect 289538 339804 289544 339816
rect 289596 339804 289602 339856
rect 221918 339736 221924 339788
rect 221976 339776 221982 339788
rect 283558 339776 283564 339788
rect 221976 339748 283564 339776
rect 221976 339736 221982 339748
rect 283558 339736 283564 339748
rect 283616 339736 283622 339788
rect 222010 339668 222016 339720
rect 222068 339708 222074 339720
rect 284294 339708 284300 339720
rect 222068 339680 284300 339708
rect 222068 339668 222074 339680
rect 284294 339668 284300 339680
rect 284352 339668 284358 339720
rect 216766 339600 216772 339652
rect 216824 339640 216830 339652
rect 294782 339640 294788 339652
rect 216824 339612 294788 339640
rect 216824 339600 216830 339612
rect 294782 339600 294788 339612
rect 294840 339600 294846 339652
rect 220722 339532 220728 339584
rect 220780 339572 220786 339584
rect 309962 339572 309968 339584
rect 220780 339544 309968 339572
rect 220780 339532 220786 339544
rect 309962 339532 309968 339544
rect 310020 339532 310026 339584
rect 274634 339464 274640 339516
rect 274692 339504 274698 339516
rect 298094 339504 298100 339516
rect 274692 339476 298100 339504
rect 274692 339464 274698 339476
rect 298094 339464 298100 339476
rect 298152 339464 298158 339516
rect 176654 339396 176660 339448
rect 176712 339436 176718 339448
rect 181438 339436 181444 339448
rect 176712 339408 181444 339436
rect 176712 339396 176718 339408
rect 181438 339396 181444 339408
rect 181496 339396 181502 339448
rect 279326 339396 279332 339448
rect 279384 339396 279390 339448
rect 279418 339396 279424 339448
rect 279476 339396 279482 339448
rect 279510 339396 279516 339448
rect 279568 339396 279574 339448
rect 279602 339396 279608 339448
rect 279660 339396 279666 339448
rect 279970 339396 279976 339448
rect 280028 339436 280034 339448
rect 283742 339436 283748 339448
rect 280028 339408 283748 339436
rect 280028 339396 280034 339408
rect 283742 339396 283748 339408
rect 283800 339396 283806 339448
rect 358354 339436 358360 339448
rect 287026 339408 358360 339436
rect 279344 338824 279372 339396
rect 279436 338892 279464 339396
rect 279528 339232 279556 339396
rect 279620 339300 279648 339396
rect 287026 339300 287054 339408
rect 358354 339396 358360 339408
rect 358412 339396 358418 339448
rect 279620 339272 287054 339300
rect 284846 339232 284852 339244
rect 279528 339204 284852 339232
rect 284846 339192 284852 339204
rect 284904 339192 284910 339244
rect 280154 338920 280160 338972
rect 280212 338960 280218 338972
rect 294322 338960 294328 338972
rect 280212 338932 294328 338960
rect 280212 338920 280218 338932
rect 294322 338920 294328 338932
rect 294380 338920 294386 338972
rect 298370 338892 298376 338904
rect 279436 338864 298376 338892
rect 298370 338852 298376 338864
rect 298428 338852 298434 338904
rect 301222 338824 301228 338836
rect 279344 338796 301228 338824
rect 301222 338784 301228 338796
rect 301280 338784 301286 338836
rect 280062 338716 280068 338768
rect 280120 338756 280126 338768
rect 324958 338756 324964 338768
rect 280120 338728 324964 338756
rect 280120 338716 280126 338728
rect 324958 338716 324964 338728
rect 325016 338716 325022 338768
rect 239122 338580 239128 338632
rect 239180 338620 239186 338632
rect 239766 338620 239772 338632
rect 239180 338592 239772 338620
rect 239180 338580 239186 338592
rect 239766 338580 239772 338592
rect 239824 338580 239830 338632
rect 228634 338444 228640 338496
rect 228692 338484 228698 338496
rect 231118 338484 231124 338496
rect 228692 338456 231124 338484
rect 228692 338444 228698 338456
rect 231118 338444 231124 338456
rect 231176 338444 231182 338496
rect 217502 338308 217508 338360
rect 217560 338348 217566 338360
rect 292942 338348 292948 338360
rect 217560 338320 292948 338348
rect 217560 338308 217566 338320
rect 292942 338308 292948 338320
rect 293000 338308 293006 338360
rect 280154 338240 280160 338292
rect 280212 338280 280218 338292
rect 289906 338280 289912 338292
rect 280212 338252 289912 338280
rect 280212 338240 280218 338252
rect 289906 338240 289912 338252
rect 289964 338240 289970 338292
rect 280062 338172 280068 338224
rect 280120 338212 280126 338224
rect 291470 338212 291476 338224
rect 280120 338184 291476 338212
rect 280120 338172 280126 338184
rect 291470 338172 291476 338184
rect 291528 338172 291534 338224
rect 280154 336132 280160 336184
rect 280212 336172 280218 336184
rect 281074 336172 281080 336184
rect 280212 336144 281080 336172
rect 280212 336132 280218 336144
rect 281074 336132 281080 336144
rect 281132 336132 281138 336184
rect 503622 333888 503628 333940
rect 503680 333928 503686 333940
rect 516502 333928 516508 333940
rect 503680 333900 516508 333928
rect 503680 333888 503686 333900
rect 516502 333888 516508 333900
rect 516560 333888 516566 333940
rect 326338 330488 326344 330540
rect 326396 330528 326402 330540
rect 329190 330528 329196 330540
rect 326396 330500 329196 330528
rect 326396 330488 326402 330500
rect 329190 330488 329196 330500
rect 329248 330488 329254 330540
rect 503622 328380 503628 328432
rect 503680 328420 503686 328432
rect 517790 328420 517796 328432
rect 503680 328392 517796 328420
rect 503680 328380 503686 328392
rect 517790 328380 517796 328392
rect 517848 328380 517854 328432
rect 304534 322872 304540 322924
rect 304592 322912 304598 322924
rect 308674 322912 308680 322924
rect 304592 322884 308680 322912
rect 304592 322872 304598 322884
rect 308674 322872 308680 322884
rect 308732 322872 308738 322924
rect 503622 322872 503628 322924
rect 503680 322912 503686 322924
rect 520550 322912 520556 322924
rect 503680 322884 520556 322912
rect 503680 322872 503686 322884
rect 520550 322872 520556 322884
rect 520608 322872 520614 322924
rect 90358 320832 90364 320884
rect 90416 320872 90422 320884
rect 125594 320872 125600 320884
rect 90416 320844 125600 320872
rect 90416 320832 90422 320844
rect 125594 320832 125600 320844
rect 125652 320832 125658 320884
rect 3418 319404 3424 319456
rect 3476 319444 3482 319456
rect 98638 319444 98644 319456
rect 3476 319416 98644 319444
rect 3476 319404 3482 319416
rect 98638 319404 98644 319416
rect 98696 319404 98702 319456
rect 88978 317432 88984 317484
rect 89036 317472 89042 317484
rect 89036 317444 124904 317472
rect 89036 317432 89042 317444
rect 124876 317416 124904 317444
rect 124858 317364 124864 317416
rect 124916 317404 124922 317416
rect 228266 317404 228272 317416
rect 124916 317376 228272 317404
rect 124916 317364 124922 317376
rect 228266 317364 228272 317376
rect 228324 317364 228330 317416
rect 281810 307708 281816 307760
rect 281868 307748 281874 307760
rect 284294 307748 284300 307760
rect 281868 307720 284300 307748
rect 281868 307708 281874 307720
rect 284294 307708 284300 307720
rect 284352 307708 284358 307760
rect 329190 307708 329196 307760
rect 329248 307748 329254 307760
rect 331950 307748 331956 307760
rect 329248 307720 331956 307748
rect 329248 307708 329254 307720
rect 331950 307708 331956 307720
rect 332008 307708 332014 307760
rect 503622 304920 503628 304972
rect 503680 304960 503686 304972
rect 519262 304960 519268 304972
rect 503680 304932 519268 304960
rect 503680 304920 503686 304932
rect 519262 304920 519268 304932
rect 519320 304920 519326 304972
rect 106182 303628 106188 303680
rect 106240 303668 106246 303680
rect 129918 303668 129924 303680
rect 106240 303640 129924 303668
rect 106240 303628 106246 303640
rect 129918 303628 129924 303640
rect 129976 303628 129982 303680
rect 181438 303628 181444 303680
rect 181496 303668 181502 303680
rect 186958 303668 186964 303680
rect 181496 303640 186964 303668
rect 181496 303628 181502 303640
rect 186958 303628 186964 303640
rect 187016 303628 187022 303680
rect 306006 303560 306012 303612
rect 306064 303600 306070 303612
rect 309042 303600 309048 303612
rect 306064 303572 309048 303600
rect 306064 303560 306070 303572
rect 309042 303560 309048 303572
rect 309100 303560 309106 303612
rect 79410 303084 79416 303136
rect 79468 303124 79474 303136
rect 90358 303124 90364 303136
rect 79468 303096 90364 303124
rect 79468 303084 79474 303096
rect 90358 303084 90364 303096
rect 90416 303084 90422 303136
rect 83918 303016 83924 303068
rect 83976 303056 83982 303068
rect 106182 303056 106188 303068
rect 83976 303028 106188 303056
rect 83976 303016 83982 303028
rect 106182 303016 106188 303028
rect 106240 303016 106246 303068
rect 77846 302948 77852 303000
rect 77904 302988 77910 303000
rect 88978 302988 88984 303000
rect 77904 302960 88984 302988
rect 77904 302948 77910 302960
rect 88978 302948 88984 302960
rect 89036 302948 89042 303000
rect 126790 302948 126796 303000
rect 126848 302988 126854 303000
rect 221826 302988 221832 303000
rect 126848 302960 221832 302988
rect 126848 302948 126854 302960
rect 221826 302948 221832 302960
rect 221884 302948 221890 303000
rect 63494 302880 63500 302932
rect 63552 302920 63558 302932
rect 64322 302920 64328 302932
rect 63552 302892 64328 302920
rect 63552 302880 63558 302892
rect 64322 302880 64328 302892
rect 64380 302920 64386 302932
rect 220354 302920 220360 302932
rect 64380 302892 220360 302920
rect 64380 302880 64386 302892
rect 220354 302880 220360 302892
rect 220412 302880 220418 302932
rect 66162 302812 66168 302864
rect 66220 302852 66226 302864
rect 67174 302852 67180 302864
rect 66220 302824 67180 302852
rect 66220 302812 66226 302824
rect 67174 302812 67180 302824
rect 67232 302812 67238 302864
rect 71590 302812 71596 302864
rect 71648 302852 71654 302864
rect 72142 302852 72148 302864
rect 71648 302824 72148 302852
rect 71648 302812 71654 302824
rect 72142 302812 72148 302824
rect 72200 302812 72206 302864
rect 94314 302744 94320 302796
rect 94372 302784 94378 302796
rect 95142 302784 95148 302796
rect 94372 302756 95148 302784
rect 94372 302744 94378 302756
rect 95142 302744 95148 302756
rect 95200 302784 95206 302796
rect 95200 302756 103514 302784
rect 95200 302744 95206 302756
rect 103486 302648 103514 302756
rect 132494 302648 132500 302660
rect 103486 302620 132500 302648
rect 132494 302608 132500 302620
rect 132552 302608 132558 302660
rect 102594 302540 102600 302592
rect 102652 302580 102658 302592
rect 103422 302580 103428 302592
rect 102652 302552 103428 302580
rect 102652 302540 102658 302552
rect 103422 302540 103428 302552
rect 103480 302580 103486 302592
rect 111794 302580 111800 302592
rect 103480 302552 111800 302580
rect 103480 302540 103486 302552
rect 111794 302540 111800 302552
rect 111852 302540 111858 302592
rect 104802 302472 104808 302524
rect 104860 302512 104866 302524
rect 124214 302512 124220 302524
rect 104860 302484 124220 302512
rect 104860 302472 104866 302484
rect 124214 302472 124220 302484
rect 124272 302472 124278 302524
rect 89622 302404 89628 302456
rect 89680 302444 89686 302456
rect 124306 302444 124312 302456
rect 89680 302416 124312 302444
rect 89680 302404 89686 302416
rect 124306 302404 124312 302416
rect 124364 302404 124370 302456
rect 46842 302336 46848 302388
rect 46900 302376 46906 302388
rect 57146 302376 57152 302388
rect 46900 302348 57152 302376
rect 46900 302336 46906 302348
rect 57146 302336 57152 302348
rect 57204 302336 57210 302388
rect 92382 302336 92388 302388
rect 92440 302376 92446 302388
rect 129826 302376 129832 302388
rect 92440 302348 129832 302376
rect 92440 302336 92446 302348
rect 129826 302336 129832 302348
rect 129884 302336 129890 302388
rect 45370 302268 45376 302320
rect 45428 302308 45434 302320
rect 55582 302308 55588 302320
rect 45428 302280 55588 302308
rect 45428 302268 45434 302280
rect 55582 302268 55588 302280
rect 55640 302268 55646 302320
rect 82722 302268 82728 302320
rect 82780 302308 82786 302320
rect 95142 302308 95148 302320
rect 82780 302280 95148 302308
rect 82780 302268 82786 302280
rect 95142 302268 95148 302280
rect 95200 302268 95206 302320
rect 88242 302200 88248 302252
rect 88300 302240 88306 302252
rect 131114 302240 131120 302252
rect 88300 302212 131120 302240
rect 88300 302200 88306 302212
rect 131114 302200 131120 302212
rect 131172 302200 131178 302252
rect 95142 301452 95148 301504
rect 95200 301492 95206 301504
rect 128446 301492 128452 301504
rect 95200 301464 128452 301492
rect 95200 301452 95206 301464
rect 128446 301452 128452 301464
rect 128504 301452 128510 301504
rect 100478 301044 100484 301096
rect 100536 301084 100542 301096
rect 125778 301084 125784 301096
rect 100536 301056 125784 301084
rect 100536 301044 100542 301056
rect 125778 301044 125784 301056
rect 125836 301084 125842 301096
rect 126790 301084 126796 301096
rect 125836 301056 126796 301084
rect 125836 301044 125842 301056
rect 126790 301044 126796 301056
rect 126848 301044 126854 301096
rect 98638 300976 98644 301028
rect 98696 301016 98702 301028
rect 131298 301016 131304 301028
rect 98696 300988 131304 301016
rect 98696 300976 98702 300988
rect 131298 300976 131304 300988
rect 131356 300976 131362 301028
rect 46750 300908 46756 300960
rect 46808 300948 46814 300960
rect 53926 300948 53932 300960
rect 46808 300920 53932 300948
rect 46808 300908 46814 300920
rect 53926 300908 53932 300920
rect 53984 300908 53990 300960
rect 91002 300908 91008 300960
rect 91060 300948 91066 300960
rect 128354 300948 128360 300960
rect 91060 300920 128360 300948
rect 91060 300908 91066 300920
rect 128354 300908 128360 300920
rect 128412 300908 128418 300960
rect 47854 300840 47860 300892
rect 47912 300880 47918 300892
rect 58894 300880 58900 300892
rect 47912 300852 58900 300880
rect 47912 300840 47918 300852
rect 58894 300840 58900 300852
rect 58952 300840 58958 300892
rect 86126 300840 86132 300892
rect 86184 300880 86190 300892
rect 86862 300880 86868 300892
rect 86184 300852 86868 300880
rect 86184 300840 86190 300852
rect 86862 300840 86868 300852
rect 86920 300880 86926 300892
rect 129734 300880 129740 300892
rect 86920 300852 129740 300880
rect 86920 300840 86926 300852
rect 129734 300840 129740 300852
rect 129792 300840 129798 300892
rect 128446 300772 128452 300824
rect 128504 300812 128510 300824
rect 128998 300812 129004 300824
rect 128504 300784 129004 300812
rect 128504 300772 128510 300784
rect 128998 300772 129004 300784
rect 129056 300812 129062 300824
rect 228634 300812 228640 300824
rect 129056 300784 228640 300812
rect 129056 300772 129062 300784
rect 228634 300772 228640 300784
rect 228692 300772 228698 300824
rect 47578 299548 47584 299600
rect 47636 299588 47642 299600
rect 47636 299560 55214 299588
rect 47636 299548 47642 299560
rect 50246 299480 50252 299532
rect 50304 299520 50310 299532
rect 52454 299520 52460 299532
rect 50304 299492 52460 299520
rect 50304 299480 50310 299492
rect 52454 299480 52460 299492
rect 52512 299480 52518 299532
rect 55186 299520 55214 299560
rect 100294 299520 100300 299532
rect 55186 299492 100300 299520
rect 100294 299480 100300 299492
rect 100352 299480 100358 299532
rect 357342 299480 357348 299532
rect 357400 299480 357406 299532
rect 357360 299328 357388 299480
rect 531958 299412 531964 299464
rect 532016 299452 532022 299464
rect 580166 299452 580172 299464
rect 532016 299424 580172 299452
rect 532016 299412 532022 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 357342 299276 357348 299328
rect 357400 299276 357406 299328
rect 281902 298120 281908 298172
rect 281960 298160 281966 298172
rect 292666 298160 292672 298172
rect 281960 298132 292672 298160
rect 281960 298120 281966 298132
rect 292666 298120 292672 298132
rect 292724 298120 292730 298172
rect 309042 298052 309048 298104
rect 309100 298092 309106 298104
rect 315574 298092 315580 298104
rect 309100 298064 315580 298092
rect 309100 298052 309106 298064
rect 315574 298052 315580 298064
rect 315632 298052 315638 298104
rect 503622 298052 503628 298104
rect 503680 298092 503686 298104
rect 516410 298092 516416 298104
rect 503680 298064 516416 298092
rect 503680 298052 503686 298064
rect 516410 298052 516416 298064
rect 516468 298052 516474 298104
rect 331950 295332 331956 295384
rect 332008 295372 332014 295384
rect 337378 295372 337384 295384
rect 332008 295344 337384 295372
rect 332008 295332 332014 295344
rect 337378 295332 337384 295344
rect 337436 295332 337442 295384
rect 281810 292544 281816 292596
rect 281868 292584 281874 292596
rect 284294 292584 284300 292596
rect 281868 292556 284300 292584
rect 281868 292544 281874 292556
rect 284294 292544 284300 292556
rect 284352 292544 284358 292596
rect 503622 292476 503628 292528
rect 503680 292516 503686 292528
rect 519170 292516 519176 292528
rect 503680 292488 519176 292516
rect 503680 292476 503686 292488
rect 519170 292476 519176 292488
rect 519228 292476 519234 292528
rect 281902 291184 281908 291236
rect 281960 291224 281966 291236
rect 284478 291224 284484 291236
rect 281960 291196 284484 291224
rect 281960 291184 281966 291196
rect 284478 291184 284484 291196
rect 284536 291184 284542 291236
rect 281902 289824 281908 289876
rect 281960 289864 281966 289876
rect 284570 289864 284576 289876
rect 281960 289836 284576 289864
rect 281960 289824 281966 289836
rect 284570 289824 284576 289836
rect 284628 289824 284634 289876
rect 281902 288396 281908 288448
rect 281960 288436 281966 288448
rect 294046 288436 294052 288448
rect 281960 288408 294052 288436
rect 281960 288396 281966 288408
rect 294046 288396 294052 288408
rect 294104 288396 294110 288448
rect 339218 288328 339224 288380
rect 339276 288368 339282 288380
rect 357526 288368 357532 288380
rect 339276 288340 357532 288368
rect 339276 288328 339282 288340
rect 357526 288328 357532 288340
rect 357584 288328 357590 288380
rect 503622 286968 503628 287020
rect 503680 287008 503686 287020
rect 520458 287008 520464 287020
rect 503680 286980 520464 287008
rect 503680 286968 503686 286980
rect 520458 286968 520464 286980
rect 520516 286968 520522 287020
rect 337378 285676 337384 285728
rect 337436 285716 337442 285728
rect 342254 285716 342260 285728
rect 337436 285688 342260 285716
rect 337436 285676 337442 285688
rect 342254 285676 342260 285688
rect 342312 285676 342318 285728
rect 342898 282820 342904 282872
rect 342956 282860 342962 282872
rect 357526 282860 357532 282872
rect 342956 282832 357532 282860
rect 342956 282820 342962 282832
rect 357526 282820 357532 282832
rect 357584 282820 357590 282872
rect 342254 279420 342260 279472
rect 342312 279460 342318 279472
rect 351178 279460 351184 279472
rect 342312 279432 351184 279460
rect 342312 279420 342318 279432
rect 351178 279420 351184 279432
rect 351236 279420 351242 279472
rect 285030 277312 285036 277364
rect 285088 277352 285094 277364
rect 357526 277352 357532 277364
rect 285088 277324 357532 277352
rect 285088 277312 285094 277324
rect 357526 277312 357532 277324
rect 357584 277312 357590 277364
rect 315574 275272 315580 275324
rect 315632 275312 315638 275324
rect 318242 275312 318248 275324
rect 315632 275284 318248 275312
rect 315632 275272 315638 275284
rect 318242 275272 318248 275284
rect 318300 275272 318306 275324
rect 503622 274592 503628 274644
rect 503680 274632 503686 274644
rect 516318 274632 516324 274644
rect 503680 274604 516324 274632
rect 503680 274592 503686 274604
rect 516318 274592 516324 274604
rect 516376 274592 516382 274644
rect 289538 273164 289544 273216
rect 289596 273204 289602 273216
rect 357526 273204 357532 273216
rect 289596 273176 357532 273204
rect 289596 273164 289602 273176
rect 357526 273164 357532 273176
rect 357584 273164 357590 273216
rect 307294 271804 307300 271856
rect 307352 271844 307358 271856
rect 357526 271844 357532 271856
rect 307352 271816 357532 271844
rect 307352 271804 307358 271816
rect 357526 271804 357532 271816
rect 357584 271804 357590 271856
rect 290642 270444 290648 270496
rect 290700 270484 290706 270496
rect 357526 270484 357532 270496
rect 290700 270456 357532 270484
rect 290700 270444 290706 270456
rect 357526 270444 357532 270456
rect 357584 270444 357590 270496
rect 282086 269016 282092 269068
rect 282144 269056 282150 269068
rect 284846 269056 284852 269068
rect 282144 269028 284852 269056
rect 282144 269016 282150 269028
rect 284846 269016 284852 269028
rect 284904 269016 284910 269068
rect 282822 268948 282828 269000
rect 282880 268988 282886 269000
rect 287238 268988 287244 269000
rect 282880 268960 287244 268988
rect 282880 268948 282886 268960
rect 287238 268948 287244 268960
rect 287296 268948 287302 269000
rect 3418 267656 3424 267708
rect 3476 267696 3482 267708
rect 47578 267696 47584 267708
rect 3476 267668 47584 267696
rect 3476 267656 3482 267668
rect 47578 267656 47584 267668
rect 47636 267656 47642 267708
rect 282822 266296 282828 266348
rect 282880 266336 282886 266348
rect 295702 266336 295708 266348
rect 282880 266308 295708 266336
rect 282880 266296 282886 266308
rect 295702 266296 295708 266308
rect 295760 266296 295766 266348
rect 282822 264868 282828 264920
rect 282880 264908 282886 264920
rect 294322 264908 294328 264920
rect 282880 264880 294328 264908
rect 282880 264868 282886 264880
rect 294322 264868 294328 264880
rect 294380 264868 294386 264920
rect 282730 263508 282736 263560
rect 282788 263548 282794 263560
rect 292942 263548 292948 263560
rect 282788 263520 292948 263548
rect 282788 263508 282794 263520
rect 292942 263508 292948 263520
rect 293000 263508 293006 263560
rect 282822 263440 282828 263492
rect 282880 263480 282886 263492
rect 291562 263480 291568 263492
rect 282880 263452 291568 263480
rect 282880 263440 282886 263452
rect 291562 263440 291568 263452
rect 291620 263440 291626 263492
rect 282822 262148 282828 262200
rect 282880 262188 282886 262200
rect 288710 262188 288716 262200
rect 282880 262160 288716 262188
rect 282880 262148 282886 262160
rect 288710 262148 288716 262160
rect 288768 262148 288774 262200
rect 325050 262148 325056 262200
rect 325108 262188 325114 262200
rect 357526 262188 357532 262200
rect 325108 262160 357532 262188
rect 325108 262148 325114 262160
rect 357526 262148 357532 262160
rect 357584 262148 357590 262200
rect 282822 260788 282828 260840
rect 282880 260828 282886 260840
rect 301038 260828 301044 260840
rect 282880 260800 301044 260828
rect 282880 260788 282886 260800
rect 301038 260788 301044 260800
rect 301096 260788 301102 260840
rect 318242 260788 318248 260840
rect 318300 260828 318306 260840
rect 323762 260828 323768 260840
rect 318300 260800 323768 260828
rect 318300 260788 318306 260800
rect 323762 260788 323768 260800
rect 323820 260788 323826 260840
rect 186958 259360 186964 259412
rect 187016 259400 187022 259412
rect 189718 259400 189724 259412
rect 187016 259372 189724 259400
rect 187016 259360 187022 259372
rect 189718 259360 189724 259372
rect 189776 259360 189782 259412
rect 282822 259360 282828 259412
rect 282880 259400 282886 259412
rect 302510 259400 302516 259412
rect 282880 259372 302516 259400
rect 282880 259360 282886 259372
rect 302510 259360 302516 259372
rect 302568 259360 302574 259412
rect 282638 259292 282644 259344
rect 282696 259332 282702 259344
rect 299566 259332 299572 259344
rect 282696 259304 299572 259332
rect 282696 259292 282702 259304
rect 299566 259292 299572 259304
rect 299624 259292 299630 259344
rect 282730 259224 282736 259276
rect 282788 259264 282794 259276
rect 292850 259264 292856 259276
rect 282788 259236 292856 259264
rect 282788 259224 282794 259236
rect 292850 259224 292856 259236
rect 292908 259224 292914 259276
rect 282730 258000 282736 258052
rect 282788 258040 282794 258052
rect 299658 258040 299664 258052
rect 282788 258012 299664 258040
rect 282788 258000 282794 258012
rect 299658 258000 299664 258012
rect 299716 258000 299722 258052
rect 282822 257932 282828 257984
rect 282880 257972 282886 257984
rect 298278 257972 298284 257984
rect 282880 257944 298284 257972
rect 282880 257932 282886 257944
rect 298278 257932 298284 257944
rect 298336 257932 298342 257984
rect 282638 256640 282644 256692
rect 282696 256680 282702 256692
rect 299474 256680 299480 256692
rect 282696 256652 299480 256680
rect 282696 256640 282702 256652
rect 299474 256640 299480 256652
rect 299532 256640 299538 256692
rect 300394 256640 300400 256692
rect 300452 256680 300458 256692
rect 357526 256680 357532 256692
rect 300452 256652 357532 256680
rect 300452 256640 300458 256652
rect 357526 256640 357532 256652
rect 357584 256640 357590 256692
rect 282822 256572 282828 256624
rect 282880 256612 282886 256624
rect 298186 256612 298192 256624
rect 282880 256584 298192 256612
rect 282880 256572 282886 256584
rect 298186 256572 298192 256584
rect 298244 256572 298250 256624
rect 282730 256504 282736 256556
rect 282788 256544 282794 256556
rect 296898 256544 296904 256556
rect 282788 256516 296904 256544
rect 282788 256504 282794 256516
rect 296898 256504 296904 256516
rect 296956 256504 296962 256556
rect 286594 255212 286600 255264
rect 286652 255252 286658 255264
rect 357526 255252 357532 255264
rect 286652 255224 357532 255252
rect 286652 255212 286658 255224
rect 357526 255212 357532 255224
rect 357584 255212 357590 255264
rect 282822 255144 282828 255196
rect 282880 255184 282886 255196
rect 301222 255184 301228 255196
rect 282880 255156 301228 255184
rect 282880 255144 282886 255156
rect 301222 255144 301228 255156
rect 301280 255144 301286 255196
rect 282638 253852 282644 253904
rect 282696 253892 282702 253904
rect 302326 253892 302332 253904
rect 282696 253864 302332 253892
rect 282696 253852 282702 253864
rect 302326 253852 302332 253864
rect 302384 253852 302390 253904
rect 282730 253784 282736 253836
rect 282788 253824 282794 253836
rect 298370 253824 298376 253836
rect 282788 253796 298376 253824
rect 282788 253784 282794 253796
rect 298370 253784 298376 253796
rect 298428 253784 298434 253836
rect 282822 253716 282828 253768
rect 282880 253756 282886 253768
rect 292574 253756 292580 253768
rect 282880 253728 292580 253756
rect 282880 253716 282886 253728
rect 292574 253716 292580 253728
rect 292632 253716 292638 253768
rect 282730 252492 282736 252544
rect 282788 252532 282794 252544
rect 303706 252532 303712 252544
rect 282788 252504 303712 252532
rect 282788 252492 282794 252504
rect 303706 252492 303712 252504
rect 303764 252492 303770 252544
rect 282822 252424 282828 252476
rect 282880 252464 282886 252476
rect 300946 252464 300952 252476
rect 282880 252436 300952 252464
rect 282880 252424 282886 252436
rect 300946 252424 300952 252436
rect 301004 252424 301010 252476
rect 282822 251132 282828 251184
rect 282880 251172 282886 251184
rect 302418 251172 302424 251184
rect 282880 251144 302424 251172
rect 282880 251132 282886 251144
rect 302418 251132 302424 251144
rect 302476 251132 302482 251184
rect 309962 251132 309968 251184
rect 310020 251172 310026 251184
rect 357526 251172 357532 251184
rect 310020 251144 357532 251172
rect 310020 251132 310026 251144
rect 357526 251132 357532 251144
rect 357584 251132 357590 251184
rect 502794 251132 502800 251184
rect 502852 251172 502858 251184
rect 505094 251172 505100 251184
rect 502852 251144 505100 251172
rect 502852 251132 502858 251144
rect 505094 251132 505100 251144
rect 505152 251132 505158 251184
rect 282730 251064 282736 251116
rect 282788 251104 282794 251116
rect 298094 251104 298100 251116
rect 282788 251076 298100 251104
rect 282788 251064 282794 251076
rect 298094 251064 298100 251076
rect 298152 251064 298158 251116
rect 282546 250996 282552 251048
rect 282604 251036 282610 251048
rect 285674 251036 285680 251048
rect 282604 251008 285680 251036
rect 282604 250996 282610 251008
rect 285674 250996 285680 251008
rect 285732 250996 285738 251048
rect 308674 250452 308680 250504
rect 308732 250492 308738 250504
rect 319714 250492 319720 250504
rect 308732 250464 319720 250492
rect 308732 250452 308738 250464
rect 319714 250452 319720 250464
rect 319772 250452 319778 250504
rect 282822 249704 282828 249756
rect 282880 249744 282886 249756
rect 295518 249744 295524 249756
rect 282880 249716 295524 249744
rect 282880 249704 282886 249716
rect 295518 249704 295524 249716
rect 295576 249704 295582 249756
rect 282730 249636 282736 249688
rect 282788 249676 282794 249688
rect 292758 249676 292764 249688
rect 282788 249648 292764 249676
rect 282788 249636 282794 249648
rect 292758 249636 292764 249648
rect 292816 249636 292822 249688
rect 282638 248072 282644 248124
rect 282696 248112 282702 248124
rect 285858 248112 285864 248124
rect 282696 248084 285864 248112
rect 282696 248072 282702 248084
rect 285858 248072 285864 248084
rect 285916 248072 285922 248124
rect 282822 246984 282828 247036
rect 282880 247024 282886 247036
rect 289906 247024 289912 247036
rect 282880 246996 289912 247024
rect 282880 246984 282886 246996
rect 289906 246984 289912 246996
rect 289964 246984 289970 247036
rect 322290 246984 322296 247036
rect 322348 247024 322354 247036
rect 357526 247024 357532 247036
rect 322348 246996 357532 247024
rect 322348 246984 322354 246996
rect 357526 246984 357532 246996
rect 357584 246984 357590 247036
rect 321002 245556 321008 245608
rect 321060 245596 321066 245608
rect 357526 245596 357532 245608
rect 321060 245568 357532 245596
rect 321060 245556 321066 245568
rect 357526 245556 357532 245568
rect 357584 245556 357590 245608
rect 299106 244876 299112 244928
rect 299164 244916 299170 244928
rect 355686 244916 355692 244928
rect 299164 244888 355692 244916
rect 299164 244876 299170 244888
rect 355686 244876 355692 244888
rect 355744 244876 355750 244928
rect 530578 244876 530584 244928
rect 530636 244916 530642 244928
rect 580166 244916 580172 244928
rect 530636 244888 580172 244916
rect 530636 244876 530642 244888
rect 580166 244876 580172 244888
rect 580224 244876 580230 244928
rect 50338 244196 50344 244248
rect 50396 244236 50402 244248
rect 50706 244236 50712 244248
rect 50396 244208 50712 244236
rect 50396 244196 50402 244208
rect 50706 244196 50712 244208
rect 50764 244196 50770 244248
rect 323762 244196 323768 244248
rect 323820 244236 323826 244248
rect 326338 244236 326344 244248
rect 323820 244208 326344 244236
rect 323820 244196 323826 244208
rect 326338 244196 326344 244208
rect 326396 244196 326402 244248
rect 357526 244236 357532 244248
rect 335326 244208 357532 244236
rect 319530 244128 319536 244180
rect 319588 244168 319594 244180
rect 335326 244168 335354 244208
rect 357526 244196 357532 244208
rect 357584 244196 357590 244248
rect 319588 244140 335354 244168
rect 319588 244128 319594 244140
rect 305822 240048 305828 240100
rect 305880 240088 305886 240100
rect 357526 240088 357532 240100
rect 305880 240060 357532 240088
rect 305880 240048 305886 240060
rect 357526 240048 357532 240060
rect 357584 240048 357590 240100
rect 81434 238688 81440 238740
rect 81492 238728 81498 238740
rect 221734 238728 221740 238740
rect 81492 238700 221740 238728
rect 81492 238688 81498 238700
rect 221734 238688 221740 238700
rect 221792 238688 221798 238740
rect 282822 238688 282828 238740
rect 282880 238728 282886 238740
rect 291470 238728 291476 238740
rect 282880 238700 291476 238728
rect 282880 238688 282886 238700
rect 291470 238688 291476 238700
rect 291528 238688 291534 238740
rect 88978 238620 88984 238672
rect 89036 238660 89042 238672
rect 221642 238660 221648 238672
rect 89036 238632 221648 238660
rect 89036 238620 89042 238632
rect 221642 238620 221648 238632
rect 221700 238620 221706 238672
rect 97902 238552 97908 238604
rect 97960 238592 97966 238604
rect 228450 238592 228456 238604
rect 97960 238564 228456 238592
rect 97960 238552 97966 238564
rect 228450 238552 228456 238564
rect 228508 238552 228514 238604
rect 86862 238484 86868 238536
rect 86920 238524 86926 238536
rect 209222 238524 209228 238536
rect 86920 238496 209228 238524
rect 86920 238484 86926 238496
rect 209222 238484 209228 238496
rect 209280 238484 209286 238536
rect 88242 238416 88248 238468
rect 88300 238456 88306 238468
rect 209314 238456 209320 238468
rect 88300 238428 209320 238456
rect 88300 238416 88306 238428
rect 209314 238416 209320 238428
rect 209372 238416 209378 238468
rect 102134 238348 102140 238400
rect 102192 238388 102198 238400
rect 220170 238388 220176 238400
rect 102192 238360 220176 238388
rect 102192 238348 102198 238360
rect 220170 238348 220176 238360
rect 220228 238348 220234 238400
rect 104802 238280 104808 238332
rect 104860 238320 104866 238332
rect 217502 238320 217508 238332
rect 104860 238292 217508 238320
rect 104860 238280 104866 238292
rect 217502 238280 217508 238292
rect 217560 238280 217566 238332
rect 99374 238212 99380 238264
rect 99432 238252 99438 238264
rect 211982 238252 211988 238264
rect 99432 238224 211988 238252
rect 99432 238212 99438 238224
rect 211982 238212 211988 238224
rect 212040 238212 212046 238264
rect 106182 238144 106188 238196
rect 106240 238184 106246 238196
rect 217410 238184 217416 238196
rect 106240 238156 217416 238184
rect 106240 238144 106246 238156
rect 217410 238144 217416 238156
rect 217468 238144 217474 238196
rect 98638 238076 98644 238128
rect 98696 238116 98702 238128
rect 209130 238116 209136 238128
rect 98696 238088 209136 238116
rect 98696 238076 98702 238088
rect 209130 238076 209136 238088
rect 209188 238076 209194 238128
rect 108298 238008 108304 238060
rect 108356 238048 108362 238060
rect 217318 238048 217324 238060
rect 108356 238020 217324 238048
rect 108356 238008 108362 238020
rect 217318 238008 217324 238020
rect 217376 238008 217382 238060
rect 281534 235900 281540 235952
rect 281592 235940 281598 235952
rect 283742 235940 283748 235952
rect 281592 235912 283748 235940
rect 281592 235900 281598 235912
rect 283742 235900 283748 235912
rect 283800 235900 283806 235952
rect 293310 235900 293316 235952
rect 293368 235940 293374 235952
rect 357526 235940 357532 235952
rect 293368 235912 357532 235940
rect 293368 235900 293374 235912
rect 357526 235900 357532 235912
rect 357584 235900 357590 235952
rect 189718 234540 189724 234592
rect 189776 234580 189782 234592
rect 192478 234580 192484 234592
rect 189776 234552 192484 234580
rect 189776 234540 189782 234552
rect 192478 234540 192484 234552
rect 192536 234540 192542 234592
rect 314102 231752 314108 231804
rect 314160 231792 314166 231804
rect 357526 231792 357532 231804
rect 314160 231764 357532 231792
rect 314160 231752 314166 231764
rect 357526 231752 357532 231764
rect 357584 231752 357590 231804
rect 294782 226244 294788 226296
rect 294840 226284 294846 226296
rect 357710 226284 357716 226296
rect 294840 226256 357716 226284
rect 294840 226244 294846 226256
rect 357710 226244 357716 226256
rect 357768 226244 357774 226296
rect 311342 226176 311348 226228
rect 311400 226216 311406 226228
rect 357526 226216 357532 226228
rect 311400 226188 357532 226216
rect 311400 226176 311406 226188
rect 357526 226176 357532 226188
rect 357584 226176 357590 226228
rect 296070 224884 296076 224936
rect 296128 224924 296134 224936
rect 357526 224924 357532 224936
rect 296128 224896 357532 224924
rect 296128 224884 296134 224896
rect 357526 224884 357532 224896
rect 357584 224884 357590 224936
rect 290550 223524 290556 223576
rect 290608 223564 290614 223576
rect 357526 223564 357532 223576
rect 290608 223536 357532 223564
rect 290608 223524 290614 223536
rect 357526 223524 357532 223536
rect 357584 223524 357590 223576
rect 307110 222096 307116 222148
rect 307168 222136 307174 222148
rect 357710 222136 357716 222148
rect 307168 222108 357716 222136
rect 307168 222096 307174 222108
rect 357710 222096 357716 222108
rect 357768 222096 357774 222148
rect 336550 222028 336556 222080
rect 336608 222068 336614 222080
rect 357526 222068 357532 222080
rect 336608 222040 357532 222068
rect 336608 222028 336614 222040
rect 357526 222028 357532 222040
rect 357584 222028 357590 222080
rect 308490 218016 308496 218068
rect 308548 218056 308554 218068
rect 314654 218056 314660 218068
rect 308548 218028 314660 218056
rect 308548 218016 308554 218028
rect 314654 218016 314660 218028
rect 314712 218016 314718 218068
rect 287974 217948 287980 218000
rect 288032 217988 288038 218000
rect 357526 217988 357532 218000
rect 288032 217960 357532 217988
rect 288032 217948 288038 217960
rect 357526 217948 357532 217960
rect 357584 217948 357590 218000
rect 327718 216588 327724 216640
rect 327776 216628 327782 216640
rect 357526 216628 357532 216640
rect 327776 216600 357532 216628
rect 327776 216588 327782 216600
rect 357526 216588 357532 216600
rect 357584 216588 357590 216640
rect 303062 215228 303068 215280
rect 303120 215268 303126 215280
rect 357526 215268 357532 215280
rect 303120 215240 357532 215268
rect 303120 215228 303126 215240
rect 357526 215228 357532 215240
rect 357584 215228 357590 215280
rect 3418 213936 3424 213988
rect 3476 213976 3482 213988
rect 102778 213976 102784 213988
rect 3476 213948 102784 213976
rect 3476 213936 3482 213948
rect 102778 213936 102784 213948
rect 102836 213936 102842 213988
rect 298830 212440 298836 212492
rect 298888 212480 298894 212492
rect 357526 212480 357532 212492
rect 298888 212452 357532 212480
rect 298888 212440 298894 212452
rect 357526 212440 357532 212452
rect 357584 212440 357590 212492
rect 319714 212372 319720 212424
rect 319772 212412 319778 212424
rect 321922 212412 321928 212424
rect 319772 212384 321928 212412
rect 319772 212372 319778 212384
rect 321922 212372 321928 212384
rect 321980 212372 321986 212424
rect 314654 211760 314660 211812
rect 314712 211800 314718 211812
rect 322382 211800 322388 211812
rect 314712 211772 322388 211800
rect 314712 211760 314718 211772
rect 322382 211760 322388 211772
rect 322440 211760 322446 211812
rect 320818 211080 320824 211132
rect 320876 211120 320882 211132
rect 357526 211120 357532 211132
rect 320876 211092 357532 211120
rect 320876 211080 320882 211092
rect 357526 211080 357532 211092
rect 357584 211080 357590 211132
rect 314010 209720 314016 209772
rect 314068 209760 314074 209772
rect 357526 209760 357532 209772
rect 314068 209732 357532 209760
rect 314068 209720 314074 209732
rect 357526 209720 357532 209732
rect 357584 209720 357590 209772
rect 102778 209040 102784 209092
rect 102836 209080 102842 209092
rect 111702 209080 111708 209092
rect 102836 209052 111708 209080
rect 102836 209040 102842 209052
rect 111702 209040 111708 209052
rect 111760 209040 111766 209092
rect 289354 208292 289360 208344
rect 289412 208332 289418 208344
rect 357526 208332 357532 208344
rect 289412 208304 357532 208332
rect 289412 208292 289418 208304
rect 357526 208292 357532 208304
rect 357584 208292 357590 208344
rect 192478 207000 192484 207052
rect 192536 207040 192542 207052
rect 197354 207040 197360 207052
rect 192536 207012 197360 207040
rect 192536 207000 192542 207012
rect 197354 207000 197360 207012
rect 197412 207000 197418 207052
rect 289262 206932 289268 206984
rect 289320 206972 289326 206984
rect 357526 206972 357532 206984
rect 289320 206944 357532 206972
rect 289320 206932 289326 206944
rect 357526 206932 357532 206944
rect 357584 206932 357590 206984
rect 334618 206864 334624 206916
rect 334676 206904 334682 206916
rect 334676 206876 354674 206904
rect 334676 206864 334682 206876
rect 354646 206700 354674 206876
rect 357526 206700 357532 206712
rect 354646 206672 357532 206700
rect 357526 206660 357532 206672
rect 357584 206660 357590 206712
rect 529198 206252 529204 206304
rect 529256 206292 529262 206304
rect 580166 206292 580172 206304
rect 529256 206264 580172 206292
rect 529256 206252 529262 206264
rect 580166 206252 580172 206264
rect 580224 206252 580230 206304
rect 289078 205572 289084 205624
rect 289136 205612 289142 205624
rect 357526 205612 357532 205624
rect 289136 205584 357532 205612
rect 289136 205572 289142 205584
rect 357526 205572 357532 205584
rect 357584 205572 357590 205624
rect 313918 204212 313924 204264
rect 313976 204252 313982 204264
rect 357526 204252 357532 204264
rect 313976 204224 357532 204252
rect 313976 204212 313982 204224
rect 357526 204212 357532 204224
rect 357584 204212 357590 204264
rect 321922 204144 321928 204196
rect 321980 204184 321986 204196
rect 326430 204184 326436 204196
rect 321980 204156 326436 204184
rect 321980 204144 321986 204156
rect 326430 204144 326436 204156
rect 326488 204144 326494 204196
rect 326338 202784 326344 202836
rect 326396 202824 326402 202836
rect 330478 202824 330484 202836
rect 326396 202796 330484 202824
rect 326396 202784 326402 202796
rect 330478 202784 330484 202796
rect 330536 202784 330542 202836
rect 197354 202104 197360 202156
rect 197412 202144 197418 202156
rect 226058 202144 226064 202156
rect 197412 202116 226064 202144
rect 197412 202104 197418 202116
rect 226058 202104 226064 202116
rect 226116 202104 226122 202156
rect 322382 202104 322388 202156
rect 322440 202144 322446 202156
rect 332502 202144 332508 202156
rect 322440 202116 332508 202144
rect 322440 202104 322446 202116
rect 332502 202104 332508 202116
rect 332560 202104 332566 202156
rect 294598 201424 294604 201476
rect 294656 201464 294662 201476
rect 357526 201464 357532 201476
rect 294656 201436 357532 201464
rect 294656 201424 294662 201436
rect 357526 201424 357532 201436
rect 357584 201424 357590 201476
rect 311250 201356 311256 201408
rect 311308 201396 311314 201408
rect 311308 201368 354674 201396
rect 311308 201356 311314 201368
rect 354646 201260 354674 201368
rect 357526 201260 357532 201272
rect 354646 201232 357532 201260
rect 357526 201220 357532 201232
rect 357584 201220 357590 201272
rect 326430 198704 326436 198756
rect 326488 198744 326494 198756
rect 329098 198744 329104 198756
rect 326488 198716 329104 198744
rect 326488 198704 326494 198716
rect 329098 198704 329104 198716
rect 329156 198704 329162 198756
rect 332502 197956 332508 198008
rect 332560 197996 332566 198008
rect 352926 197996 352932 198008
rect 332560 197968 352932 197996
rect 332560 197956 332566 197968
rect 352926 197956 352932 197968
rect 352984 197956 352990 198008
rect 287790 195916 287796 195968
rect 287848 195956 287854 195968
rect 357526 195956 357532 195968
rect 287848 195928 357532 195956
rect 287848 195916 287854 195928
rect 357526 195916 357532 195928
rect 357584 195916 357590 195968
rect 226058 194488 226064 194540
rect 226116 194528 226122 194540
rect 229922 194528 229928 194540
rect 226116 194500 229928 194528
rect 226116 194488 226122 194500
rect 229922 194488 229928 194500
rect 229980 194488 229986 194540
rect 282822 191836 282828 191888
rect 282880 191876 282886 191888
rect 292574 191876 292580 191888
rect 282880 191848 292580 191876
rect 282880 191836 282886 191848
rect 292574 191836 292580 191848
rect 292632 191836 292638 191888
rect 351178 189728 351184 189780
rect 351236 189768 351242 189780
rect 358262 189768 358268 189780
rect 351236 189740 358268 189768
rect 351236 189728 351242 189740
rect 358262 189728 358268 189740
rect 358320 189728 358326 189780
rect 329098 189048 329104 189100
rect 329156 189088 329162 189100
rect 338022 189088 338028 189100
rect 329156 189060 338028 189088
rect 329156 189048 329162 189060
rect 338022 189048 338028 189060
rect 338080 189048 338086 189100
rect 38562 186940 38568 186992
rect 38620 186980 38626 186992
rect 238386 186980 238392 186992
rect 38620 186952 238392 186980
rect 38620 186940 38626 186952
rect 238386 186940 238392 186952
rect 238444 186940 238450 186992
rect 111702 185580 111708 185632
rect 111760 185620 111766 185632
rect 129090 185620 129096 185632
rect 111760 185592 129096 185620
rect 111760 185580 111766 185592
rect 129090 185580 129096 185592
rect 129148 185580 129154 185632
rect 54478 184900 54484 184952
rect 54536 184940 54542 184952
rect 124214 184940 124220 184952
rect 54536 184912 124220 184940
rect 54536 184900 54542 184912
rect 124214 184900 124220 184912
rect 124272 184940 124278 184952
rect 124398 184940 124404 184952
rect 124272 184912 124404 184940
rect 124272 184900 124278 184912
rect 124398 184900 124404 184912
rect 124456 184900 124462 184952
rect 330478 184152 330484 184204
rect 330536 184192 330542 184204
rect 351178 184192 351184 184204
rect 330536 184164 351184 184192
rect 330536 184152 330542 184164
rect 351178 184152 351184 184164
rect 351236 184152 351242 184204
rect 352926 184152 352932 184204
rect 352984 184192 352990 184204
rect 359734 184192 359740 184204
rect 352984 184164 359740 184192
rect 352984 184152 352990 184164
rect 359734 184152 359740 184164
rect 359792 184152 359798 184204
rect 338022 181432 338028 181484
rect 338080 181472 338086 181484
rect 358630 181472 358636 181484
rect 338080 181444 358636 181472
rect 338080 181432 338086 181444
rect 358630 181432 358636 181444
rect 358688 181432 358694 181484
rect 350166 180616 350172 180668
rect 350224 180656 350230 180668
rect 379606 180656 379612 180668
rect 350224 180628 379612 180656
rect 350224 180616 350230 180628
rect 379606 180616 379612 180628
rect 379664 180616 379670 180668
rect 488442 180616 488448 180668
rect 488500 180656 488506 180668
rect 522574 180656 522580 180668
rect 488500 180628 522580 180656
rect 488500 180616 488506 180628
rect 522574 180616 522580 180628
rect 522632 180616 522638 180668
rect 347130 180548 347136 180600
rect 347188 180588 347194 180600
rect 380802 180588 380808 180600
rect 347188 180560 380808 180588
rect 347188 180548 347194 180560
rect 380802 180548 380808 180560
rect 380860 180548 380866 180600
rect 492490 180548 492496 180600
rect 492548 180588 492554 180600
rect 525794 180588 525800 180600
rect 492548 180560 525800 180588
rect 492548 180548 492554 180560
rect 525794 180548 525800 180560
rect 525852 180548 525858 180600
rect 350350 180480 350356 180532
rect 350408 180520 350414 180532
rect 384574 180520 384580 180532
rect 350408 180492 384580 180520
rect 350408 180480 350414 180492
rect 384574 180480 384580 180492
rect 384632 180480 384638 180532
rect 489546 180480 489552 180532
rect 489604 180520 489610 180532
rect 523126 180520 523132 180532
rect 489604 180492 523132 180520
rect 489604 180480 489610 180492
rect 523126 180480 523132 180492
rect 523184 180480 523190 180532
rect 344554 180412 344560 180464
rect 344612 180452 344618 180464
rect 382550 180452 382556 180464
rect 344612 180424 382556 180452
rect 344612 180412 344618 180424
rect 382550 180412 382556 180424
rect 382608 180412 382614 180464
rect 477402 180412 477408 180464
rect 477460 180452 477466 180464
rect 521838 180452 521844 180464
rect 477460 180424 521844 180452
rect 477460 180412 477466 180424
rect 521838 180412 521844 180424
rect 521896 180412 521902 180464
rect 344462 180344 344468 180396
rect 344520 180384 344526 180396
rect 383746 180384 383752 180396
rect 344520 180356 383752 180384
rect 344520 180344 344526 180356
rect 383746 180344 383752 180356
rect 383804 180344 383810 180396
rect 479426 180344 479432 180396
rect 479484 180384 479490 180396
rect 527174 180384 527180 180396
rect 479484 180356 527180 180384
rect 479484 180344 479490 180356
rect 527174 180344 527180 180356
rect 527232 180344 527238 180396
rect 336458 180276 336464 180328
rect 336516 180316 336522 180328
rect 381630 180316 381636 180328
rect 336516 180288 381636 180316
rect 336516 180276 336522 180288
rect 381630 180276 381636 180288
rect 381688 180276 381694 180328
rect 475378 180276 475384 180328
rect 475436 180316 475442 180328
rect 523218 180316 523224 180328
rect 475436 180288 523224 180316
rect 475436 180276 475442 180288
rect 523218 180276 523224 180288
rect 523276 180276 523282 180328
rect 339034 180208 339040 180260
rect 339092 180248 339098 180260
rect 385678 180248 385684 180260
rect 339092 180220 385684 180248
rect 339092 180208 339098 180220
rect 385678 180208 385684 180220
rect 385736 180208 385742 180260
rect 449066 180208 449072 180260
rect 449124 180248 449130 180260
rect 524506 180248 524512 180260
rect 449124 180220 524512 180248
rect 449124 180208 449130 180220
rect 524506 180208 524512 180220
rect 524564 180208 524570 180260
rect 338758 180140 338764 180192
rect 338816 180180 338822 180192
rect 386598 180180 386604 180192
rect 338816 180152 386604 180180
rect 338816 180140 338822 180152
rect 386598 180140 386604 180152
rect 386656 180140 386662 180192
rect 449802 180140 449808 180192
rect 449860 180180 449866 180192
rect 536834 180180 536840 180192
rect 449860 180152 536840 180180
rect 449860 180140 449866 180152
rect 536834 180140 536840 180152
rect 536892 180140 536898 180192
rect 350258 180072 350264 180124
rect 350316 180112 350322 180124
rect 377582 180112 377588 180124
rect 350316 180084 377588 180112
rect 350316 180072 350322 180084
rect 377582 180072 377588 180084
rect 377640 180072 377646 180124
rect 476114 180072 476120 180124
rect 476172 180072 476178 180124
rect 480162 180072 480168 180124
rect 480220 180112 480226 180124
rect 513466 180112 513472 180124
rect 480220 180084 513472 180112
rect 480220 180072 480226 180084
rect 513466 180072 513472 180084
rect 513524 180072 513530 180124
rect 355318 180004 355324 180056
rect 355376 180044 355382 180056
rect 375558 180044 375564 180056
rect 355376 180016 375564 180044
rect 355376 180004 355382 180016
rect 375558 180004 375564 180016
rect 375616 180004 375622 180056
rect 358078 179936 358084 179988
rect 358136 179976 358142 179988
rect 369486 179976 369492 179988
rect 358136 179948 369492 179976
rect 358136 179936 358142 179948
rect 369486 179936 369492 179948
rect 369544 179936 369550 179988
rect 476132 179976 476160 180072
rect 491110 180004 491116 180056
rect 491168 180044 491174 180056
rect 524414 180044 524420 180056
rect 491168 180016 524420 180044
rect 491168 180004 491174 180016
rect 524414 180004 524420 180016
rect 524472 180004 524478 180056
rect 503162 179976 503168 179988
rect 476132 179948 503168 179976
rect 503162 179936 503168 179948
rect 503220 179936 503226 179988
rect 351178 179868 351184 179920
rect 351236 179908 351242 179920
rect 367002 179908 367008 179920
rect 351236 179880 367008 179908
rect 351236 179868 351242 179880
rect 367002 179868 367008 179880
rect 367060 179868 367066 179920
rect 355410 179324 355416 179376
rect 355468 179364 355474 179376
rect 423398 179364 423404 179376
rect 355468 179336 423404 179364
rect 355468 179324 355474 179336
rect 423398 179324 423404 179336
rect 423456 179324 423462 179376
rect 451734 179324 451740 179376
rect 451792 179364 451798 179376
rect 539870 179364 539876 179376
rect 451792 179336 539876 179364
rect 451792 179324 451798 179336
rect 539870 179324 539876 179336
rect 539928 179324 539934 179376
rect 341794 179256 341800 179308
rect 341852 179296 341858 179308
rect 409230 179296 409236 179308
rect 341852 179268 409236 179296
rect 341852 179256 341858 179268
rect 409230 179256 409236 179268
rect 409288 179256 409294 179308
rect 455782 179256 455788 179308
rect 455840 179296 455846 179308
rect 543734 179296 543740 179308
rect 455840 179268 543740 179296
rect 455840 179256 455846 179268
rect 543734 179256 543740 179268
rect 543792 179256 543798 179308
rect 347498 179188 347504 179240
rect 347556 179228 347562 179240
rect 408218 179228 408224 179240
rect 347556 179200 408224 179228
rect 347556 179188 347562 179200
rect 408218 179188 408224 179200
rect 408276 179188 408282 179240
rect 458818 179188 458824 179240
rect 458876 179228 458882 179240
rect 545298 179228 545304 179240
rect 458876 179200 545304 179228
rect 458876 179188 458882 179200
rect 545298 179188 545304 179200
rect 545356 179188 545362 179240
rect 341518 179120 341524 179172
rect 341576 179160 341582 179172
rect 402146 179160 402152 179172
rect 341576 179132 402152 179160
rect 341576 179120 341582 179132
rect 402146 179120 402152 179132
rect 402204 179120 402210 179172
rect 459830 179120 459836 179172
rect 459888 179160 459894 179172
rect 545114 179160 545120 179172
rect 459888 179132 545120 179160
rect 459888 179120 459894 179132
rect 545114 179120 545120 179132
rect 545172 179120 545178 179172
rect 347406 179052 347412 179104
rect 347464 179092 347470 179104
rect 407206 179092 407212 179104
rect 347464 179064 407212 179092
rect 347464 179052 347470 179064
rect 407206 179052 407212 179064
rect 407264 179052 407270 179104
rect 460842 179052 460848 179104
rect 460900 179092 460906 179104
rect 543826 179092 543832 179104
rect 460900 179064 543832 179092
rect 460900 179052 460906 179064
rect 543826 179052 543832 179064
rect 543884 179052 543890 179104
rect 341702 178984 341708 179036
rect 341760 179024 341766 179036
rect 396074 179024 396080 179036
rect 341760 178996 396080 179024
rect 341760 178984 341766 178996
rect 396074 178984 396080 178996
rect 396132 178984 396138 179036
rect 463878 178984 463884 179036
rect 463936 179024 463942 179036
rect 545206 179024 545212 179036
rect 463936 178996 545212 179024
rect 463936 178984 463942 178996
rect 545206 178984 545212 178996
rect 545264 178984 545270 179036
rect 344370 178916 344376 178968
rect 344428 178956 344434 178968
rect 398098 178956 398104 178968
rect 344428 178928 398104 178956
rect 344428 178916 344434 178928
rect 398098 178916 398104 178928
rect 398156 178916 398162 178968
rect 444650 178916 444656 178968
rect 444708 178956 444714 178968
rect 520366 178956 520372 178968
rect 444708 178928 520372 178956
rect 444708 178916 444714 178928
rect 520366 178916 520372 178928
rect 520424 178916 520430 178968
rect 352742 178848 352748 178900
rect 352800 178888 352806 178900
rect 406194 178888 406200 178900
rect 352800 178860 406200 178888
rect 352800 178848 352806 178860
rect 406194 178848 406200 178860
rect 406252 178848 406258 178900
rect 443638 178848 443644 178900
rect 443696 178888 443702 178900
rect 519078 178888 519084 178900
rect 443696 178860 519084 178888
rect 443696 178848 443702 178860
rect 519078 178848 519084 178860
rect 519136 178848 519142 178900
rect 338850 178780 338856 178832
rect 338908 178820 338914 178832
rect 390002 178820 390008 178832
rect 338908 178792 390008 178820
rect 338908 178780 338914 178792
rect 390002 178780 390008 178792
rect 390060 178780 390066 178832
rect 465902 178780 465908 178832
rect 465960 178820 465966 178832
rect 541066 178820 541072 178832
rect 465960 178792 541072 178820
rect 465960 178780 465966 178792
rect 541066 178780 541072 178792
rect 541124 178780 541130 178832
rect 344278 178712 344284 178764
rect 344336 178752 344342 178764
rect 395062 178752 395068 178764
rect 344336 178724 395068 178752
rect 344336 178712 344342 178724
rect 395062 178712 395068 178724
rect 395120 178712 395126 178764
rect 446674 178712 446680 178764
rect 446732 178752 446738 178764
rect 521746 178752 521752 178764
rect 446732 178724 521752 178752
rect 446732 178712 446738 178724
rect 521746 178712 521752 178724
rect 521804 178712 521810 178764
rect 358262 178644 358268 178696
rect 358320 178684 358326 178696
rect 369118 178684 369124 178696
rect 358320 178656 369124 178684
rect 358320 178644 358326 178656
rect 369118 178644 369124 178656
rect 369176 178644 369182 178696
rect 464890 178644 464896 178696
rect 464948 178684 464954 178696
rect 538214 178684 538220 178696
rect 464948 178656 538220 178684
rect 464948 178644 464954 178656
rect 538214 178644 538220 178656
rect 538272 178644 538278 178696
rect 359734 178576 359740 178628
rect 359792 178616 359798 178628
rect 369854 178616 369860 178628
rect 359792 178588 369860 178616
rect 359792 178576 359798 178588
rect 369854 178576 369860 178588
rect 369912 178576 369918 178628
rect 442626 178576 442632 178628
rect 442684 178616 442690 178628
rect 501598 178616 501604 178628
rect 442684 178588 501604 178616
rect 442684 178576 442690 178588
rect 501598 178576 501604 178588
rect 501656 178576 501662 178628
rect 335998 178440 336004 178492
rect 336056 178480 336062 178492
rect 373810 178480 373816 178492
rect 336056 178452 373816 178480
rect 336056 178440 336062 178452
rect 373810 178440 373816 178452
rect 373868 178440 373874 178492
rect 358630 178032 358636 178084
rect 358688 178072 358694 178084
rect 358688 178044 366772 178072
rect 358688 178032 358694 178044
rect 347222 177964 347228 178016
rect 347280 178004 347286 178016
rect 347280 177976 354674 178004
rect 347280 177964 347286 177976
rect 354646 177868 354674 177976
rect 359642 177964 359648 178016
rect 359700 178004 359706 178016
rect 366358 178004 366364 178016
rect 359700 177976 366364 178004
rect 359700 177964 359706 177976
rect 366358 177964 366364 177976
rect 366416 177964 366422 178016
rect 366744 178004 366772 178044
rect 427446 178004 427452 178016
rect 366744 177976 427452 178004
rect 427446 177964 427452 177976
rect 427504 177964 427510 178016
rect 472986 177964 472992 178016
rect 473044 178004 473050 178016
rect 499574 178004 499580 178016
rect 473044 177976 499580 178004
rect 473044 177964 473050 177976
rect 499574 177964 499580 177976
rect 499632 177964 499638 178016
rect 355594 177896 355600 177948
rect 355652 177936 355658 177948
rect 370774 177936 370780 177948
rect 355652 177908 370780 177936
rect 355652 177896 355658 177908
rect 370774 177896 370780 177908
rect 370832 177896 370838 177948
rect 467926 177896 467932 177948
rect 467984 177936 467990 177948
rect 510614 177936 510620 177948
rect 467984 177908 510620 177936
rect 467984 177896 467990 177908
rect 510614 177896 510620 177908
rect 510672 177896 510678 177948
rect 365714 177868 365720 177880
rect 354646 177840 365720 177868
rect 365714 177828 365720 177840
rect 365772 177828 365778 177880
rect 367002 177828 367008 177880
rect 367060 177868 367066 177880
rect 376846 177868 376852 177880
rect 367060 177840 376852 177868
rect 367060 177828 367066 177840
rect 376846 177828 376852 177840
rect 376904 177828 376910 177880
rect 466914 177828 466920 177880
rect 466972 177868 466978 177880
rect 509326 177868 509332 177880
rect 466972 177840 509332 177868
rect 466972 177828 466978 177840
rect 509326 177828 509332 177840
rect 509384 177828 509390 177880
rect 350074 177760 350080 177812
rect 350132 177800 350138 177812
rect 404170 177800 404176 177812
rect 350132 177772 404176 177800
rect 350132 177760 350138 177772
rect 404170 177760 404176 177772
rect 404228 177760 404234 177812
rect 468938 177760 468944 177812
rect 468996 177800 469002 177812
rect 507854 177800 507860 177812
rect 468996 177772 507860 177800
rect 468996 177760 469002 177772
rect 507854 177760 507860 177772
rect 507912 177760 507918 177812
rect 349982 177692 349988 177744
rect 350040 177732 350046 177744
rect 403158 177732 403164 177744
rect 350040 177704 403164 177732
rect 350040 177692 350046 177704
rect 403158 177692 403164 177704
rect 403216 177692 403222 177744
rect 483106 177692 483112 177744
rect 483164 177732 483170 177744
rect 518434 177732 518440 177744
rect 483164 177704 518440 177732
rect 483164 177692 483170 177704
rect 518434 177692 518440 177704
rect 518492 177692 518498 177744
rect 333238 177624 333244 177676
rect 333296 177664 333302 177676
rect 368750 177664 368756 177676
rect 333296 177636 368756 177664
rect 333296 177624 333302 177636
rect 368750 177624 368756 177636
rect 368808 177624 368814 177676
rect 369854 177624 369860 177676
rect 369912 177664 369918 177676
rect 419350 177664 419356 177676
rect 369912 177636 419356 177664
rect 369912 177624 369918 177636
rect 419350 177624 419356 177636
rect 419408 177624 419414 177676
rect 486142 177624 486148 177676
rect 486200 177664 486206 177676
rect 520274 177664 520280 177676
rect 486200 177636 520280 177664
rect 486200 177624 486206 177636
rect 520274 177624 520280 177636
rect 520332 177624 520338 177676
rect 352650 177556 352656 177608
rect 352708 177596 352714 177608
rect 401134 177596 401140 177608
rect 352708 177568 401140 177596
rect 352708 177556 352714 177568
rect 401134 177556 401140 177568
rect 401192 177556 401198 177608
rect 482094 177556 482100 177608
rect 482152 177596 482158 177608
rect 516226 177596 516232 177608
rect 482152 177568 516232 177596
rect 482152 177556 482158 177568
rect 516226 177556 516232 177568
rect 516284 177556 516290 177608
rect 352558 177488 352564 177540
rect 352616 177528 352622 177540
rect 400122 177528 400128 177540
rect 352616 177500 400128 177528
rect 352616 177488 352622 177500
rect 400122 177488 400128 177500
rect 400180 177488 400186 177540
rect 485130 177488 485136 177540
rect 485188 177528 485194 177540
rect 518986 177528 518992 177540
rect 485188 177500 518992 177528
rect 485188 177488 485194 177500
rect 518986 177488 518992 177500
rect 519044 177488 519050 177540
rect 352834 177420 352840 177472
rect 352892 177460 352898 177472
rect 399110 177460 399116 177472
rect 352892 177432 399116 177460
rect 352892 177420 352898 177432
rect 399110 177420 399116 177432
rect 399168 177420 399174 177472
rect 484118 177420 484124 177472
rect 484176 177460 484182 177472
rect 517606 177460 517612 177472
rect 484176 177432 517612 177460
rect 484176 177420 484182 177432
rect 517606 177420 517612 177432
rect 517664 177420 517670 177472
rect 333330 177352 333336 177404
rect 333388 177392 333394 177404
rect 367738 177392 367744 177404
rect 333388 177364 367744 177392
rect 333388 177352 333394 177364
rect 367738 177352 367744 177364
rect 367796 177352 367802 177404
rect 369118 177352 369124 177404
rect 369176 177392 369182 177404
rect 412266 177392 412272 177404
rect 369176 177364 412272 177392
rect 369176 177352 369182 177364
rect 412266 177352 412272 177364
rect 412324 177352 412330 177404
rect 469950 177352 469956 177404
rect 470008 177392 470014 177404
rect 502978 177392 502984 177404
rect 470008 177364 502984 177392
rect 470008 177352 470014 177364
rect 502978 177352 502984 177364
rect 503036 177352 503042 177404
rect 359458 177284 359464 177336
rect 359516 177324 359522 177336
rect 388990 177324 388996 177336
rect 359516 177296 388996 177324
rect 359516 177284 359522 177296
rect 388990 177284 388996 177296
rect 389048 177284 389054 177336
rect 470962 177284 470968 177336
rect 471020 177324 471026 177336
rect 503070 177324 503076 177336
rect 471020 177296 503076 177324
rect 471020 177284 471026 177296
rect 503070 177284 503076 177296
rect 503128 177284 503134 177336
rect 333422 177216 333428 177268
rect 333480 177256 333486 177268
rect 378870 177256 378876 177268
rect 333480 177228 378876 177256
rect 333480 177216 333486 177228
rect 378870 177216 378876 177228
rect 378928 177216 378934 177268
rect 453758 177216 453764 177268
rect 453816 177256 453822 177268
rect 540974 177256 540980 177268
rect 453816 177228 540980 177256
rect 453816 177216 453822 177228
rect 540974 177216 540980 177228
rect 541032 177216 541038 177268
rect 336274 177148 336280 177200
rect 336332 177188 336338 177200
rect 394050 177188 394056 177200
rect 336332 177160 394056 177188
rect 336332 177148 336338 177160
rect 394050 177148 394056 177160
rect 394108 177148 394114 177200
rect 494238 177148 494244 177200
rect 494296 177188 494302 177200
rect 518894 177188 518900 177200
rect 494296 177160 518900 177188
rect 494296 177148 494302 177160
rect 518894 177148 518900 177160
rect 518952 177148 518958 177200
rect 336182 177080 336188 177132
rect 336240 177120 336246 177132
rect 397086 177120 397092 177132
rect 336240 177092 397092 177120
rect 336240 177080 336246 177092
rect 397086 177080 397092 177092
rect 397144 177080 397150 177132
rect 347314 176604 347320 176656
rect 347372 176644 347378 176656
rect 417326 176644 417332 176656
rect 347372 176616 417332 176644
rect 347372 176604 347378 176616
rect 417326 176604 417332 176616
rect 417384 176604 417390 176656
rect 426434 176604 426440 176656
rect 426492 176644 426498 176656
rect 513374 176644 513380 176656
rect 426492 176616 513380 176644
rect 426492 176604 426498 176616
rect 513374 176604 513380 176616
rect 513432 176604 513438 176656
rect 347038 176536 347044 176588
rect 347096 176576 347102 176588
rect 393038 176576 393044 176588
rect 347096 176548 393044 176576
rect 347096 176536 347102 176548
rect 393038 176536 393044 176548
rect 393096 176536 393102 176588
rect 445662 176536 445668 176588
rect 445720 176576 445726 176588
rect 531314 176576 531320 176588
rect 445720 176548 531320 176576
rect 445720 176536 445726 176548
rect 531314 176536 531320 176548
rect 531372 176536 531378 176588
rect 452746 176468 452752 176520
rect 452804 176508 452810 176520
rect 528554 176508 528560 176520
rect 452804 176480 528560 176508
rect 452804 176468 452810 176480
rect 528554 176468 528560 176480
rect 528612 176468 528618 176520
rect 429470 176400 429476 176452
rect 429528 176440 429534 176452
rect 505278 176440 505284 176452
rect 429528 176412 505284 176440
rect 429528 176400 429534 176412
rect 505278 176400 505284 176412
rect 505336 176400 505342 176452
rect 440602 176332 440608 176384
rect 440660 176372 440666 176384
rect 516134 176372 516140 176384
rect 440660 176344 516140 176372
rect 440660 176332 440666 176344
rect 516134 176332 516140 176344
rect 516192 176332 516198 176384
rect 434530 176264 434536 176316
rect 434588 176304 434594 176316
rect 509234 176304 509240 176316
rect 434588 176276 509240 176304
rect 434588 176264 434594 176276
rect 509234 176264 509240 176276
rect 509292 176264 509298 176316
rect 305638 175924 305644 175976
rect 305696 175964 305702 175976
rect 371050 175964 371056 175976
rect 305696 175936 371056 175964
rect 305696 175924 305702 175936
rect 371050 175924 371056 175936
rect 371108 175924 371114 175976
rect 416314 175176 416320 175228
rect 416372 175216 416378 175228
rect 505186 175216 505192 175228
rect 416372 175188 505192 175216
rect 416372 175176 416378 175188
rect 505186 175176 505192 175188
rect 505244 175176 505250 175228
rect 430482 175108 430488 175160
rect 430540 175148 430546 175160
rect 517698 175148 517704 175160
rect 430540 175120 517704 175148
rect 430540 175108 430546 175120
rect 517698 175108 517704 175120
rect 517756 175108 517762 175160
rect 447686 175040 447692 175092
rect 447744 175080 447750 175092
rect 523954 175080 523960 175092
rect 447744 175052 523960 175080
rect 447744 175040 447750 175052
rect 523954 175040 523960 175052
rect 524012 175040 524018 175092
rect 436554 174972 436560 175024
rect 436612 175012 436618 175024
rect 511350 175012 511356 175024
rect 436612 174984 511356 175012
rect 436612 174972 436618 174984
rect 511350 174972 511356 174984
rect 511408 174972 511414 175024
rect 450722 174904 450728 174956
rect 450780 174944 450786 174956
rect 512638 174944 512644 174956
rect 450780 174916 512644 174944
rect 450780 174904 450786 174916
rect 512638 174904 512644 174916
rect 512696 174904 512702 174956
rect 308398 170348 308404 170400
rect 308456 170388 308462 170400
rect 372246 170388 372252 170400
rect 308456 170360 372252 170388
rect 308456 170348 308462 170360
rect 372246 170348 372252 170360
rect 372304 170348 372310 170400
rect 282822 169736 282828 169788
rect 282880 169776 282886 169788
rect 289998 169776 290004 169788
rect 282880 169748 290004 169776
rect 282880 169736 282886 169748
rect 289998 169736 290004 169748
rect 290056 169736 290062 169788
rect 360102 169260 360108 169312
rect 360160 169300 360166 169312
rect 393774 169300 393780 169312
rect 360160 169272 393780 169300
rect 360160 169260 360166 169272
rect 393774 169260 393780 169272
rect 393832 169260 393838 169312
rect 315298 169192 315304 169244
rect 315356 169232 315362 169244
rect 377030 169232 377036 169244
rect 315356 169204 377036 169232
rect 315356 169192 315362 169204
rect 377030 169192 377036 169204
rect 377088 169192 377094 169244
rect 349982 169124 349988 169176
rect 350040 169164 350046 169176
rect 580258 169164 580264 169176
rect 350040 169136 580264 169164
rect 350040 169124 350046 169136
rect 580258 169124 580264 169136
rect 580316 169124 580322 169176
rect 349798 169056 349804 169108
rect 349856 169096 349862 169108
rect 580350 169096 580356 169108
rect 349856 169068 580356 169096
rect 349856 169056 349862 169068
rect 580350 169056 580356 169068
rect 580408 169056 580414 169108
rect 349890 168988 349896 169040
rect 349948 169028 349954 169040
rect 580534 169028 580540 169040
rect 349948 169000 580540 169028
rect 349948 168988 349954 169000
rect 580534 168988 580540 169000
rect 580592 168988 580598 169040
rect 282822 168376 282828 168428
rect 282880 168416 282886 168428
rect 290090 168416 290096 168428
rect 282880 168388 290096 168416
rect 282880 168376 282886 168388
rect 290090 168376 290096 168388
rect 290148 168376 290154 168428
rect 282454 168308 282460 168360
rect 282512 168348 282518 168360
rect 291194 168348 291200 168360
rect 282512 168320 291200 168348
rect 282512 168308 282518 168320
rect 291194 168308 291200 168320
rect 291252 168308 291258 168360
rect 282638 167016 282644 167068
rect 282696 167056 282702 167068
rect 289814 167056 289820 167068
rect 282696 167028 289820 167056
rect 282696 167016 282702 167028
rect 289814 167016 289820 167028
rect 289872 167016 289878 167068
rect 282822 166948 282828 167000
rect 282880 166988 282886 167000
rect 303614 166988 303620 167000
rect 282880 166960 303620 166988
rect 282880 166948 282886 166960
rect 303614 166948 303620 166960
rect 303672 166948 303678 167000
rect 524322 166948 524328 167000
rect 524380 166988 524386 167000
rect 580166 166988 580172 167000
rect 524380 166960 580172 166988
rect 524380 166948 524386 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 282822 165520 282828 165572
rect 282880 165560 282886 165572
rect 296806 165560 296812 165572
rect 282880 165532 296812 165560
rect 282880 165520 282886 165532
rect 296806 165520 296812 165532
rect 296864 165520 296870 165572
rect 302878 164840 302884 164892
rect 302936 164880 302942 164892
rect 368658 164880 368664 164892
rect 302936 164852 368664 164880
rect 302936 164840 302942 164852
rect 368658 164840 368664 164852
rect 368716 164840 368722 164892
rect 3418 164160 3424 164212
rect 3476 164200 3482 164212
rect 54478 164200 54484 164212
rect 3476 164172 54484 164200
rect 3476 164160 3482 164172
rect 54478 164160 54484 164172
rect 54536 164160 54542 164212
rect 282822 164160 282828 164212
rect 282880 164200 282886 164212
rect 296714 164200 296720 164212
rect 282880 164172 296720 164200
rect 282880 164160 282886 164172
rect 296714 164160 296720 164172
rect 296772 164160 296778 164212
rect 282638 164092 282644 164144
rect 282696 164132 282702 164144
rect 295334 164132 295340 164144
rect 282696 164104 295340 164132
rect 282696 164092 282702 164104
rect 295334 164092 295340 164104
rect 295392 164092 295398 164144
rect 282638 162800 282644 162852
rect 282696 162840 282702 162852
rect 302234 162840 302240 162852
rect 282696 162812 302240 162840
rect 282696 162800 282702 162812
rect 302234 162800 302240 162812
rect 302292 162800 302298 162852
rect 282822 162732 282828 162784
rect 282880 162772 282886 162784
rect 288434 162772 288440 162784
rect 282880 162744 288440 162772
rect 282880 162732 282886 162744
rect 288434 162732 288440 162744
rect 288492 162732 288498 162784
rect 324958 162120 324964 162172
rect 325016 162160 325022 162172
rect 384206 162160 384212 162172
rect 325016 162132 384212 162160
rect 325016 162120 325022 162132
rect 384206 162120 384212 162132
rect 384264 162120 384270 162172
rect 282822 161372 282828 161424
rect 282880 161412 282886 161424
rect 290182 161412 290188 161424
rect 282880 161384 290188 161412
rect 282880 161372 282886 161384
rect 290182 161372 290188 161384
rect 290240 161372 290246 161424
rect 309778 160692 309784 160744
rect 309836 160732 309842 160744
rect 373442 160732 373448 160744
rect 309836 160704 373448 160732
rect 309836 160692 309842 160704
rect 373442 160692 373448 160704
rect 373500 160692 373506 160744
rect 229830 155864 229836 155916
rect 229888 155904 229894 155916
rect 237374 155904 237380 155916
rect 229888 155876 237380 155904
rect 229888 155864 229894 155876
rect 237374 155864 237380 155876
rect 237432 155864 237438 155916
rect 229922 154504 229928 154556
rect 229980 154544 229986 154556
rect 237374 154544 237380 154556
rect 229980 154516 237380 154544
rect 229980 154504 229986 154516
rect 237374 154504 237380 154516
rect 237432 154504 237438 154556
rect 318150 151784 318156 151836
rect 318208 151824 318214 151836
rect 580166 151824 580172 151836
rect 318208 151796 580172 151824
rect 318208 151784 318214 151796
rect 580166 151784 580172 151796
rect 580224 151784 580230 151836
rect 311158 149676 311164 149728
rect 311216 149716 311222 149728
rect 374638 149716 374644 149728
rect 311216 149688 374644 149716
rect 311216 149676 311222 149688
rect 374638 149676 374644 149688
rect 374696 149676 374702 149728
rect 322198 148384 322204 148436
rect 322256 148424 322262 148436
rect 381814 148424 381820 148436
rect 322256 148396 381820 148424
rect 322256 148384 322262 148396
rect 381814 148384 381820 148396
rect 381872 148384 381878 148436
rect 319438 148316 319444 148368
rect 319496 148356 319502 148368
rect 380618 148356 380624 148368
rect 319496 148328 380624 148356
rect 319496 148316 319502 148328
rect 380618 148316 380624 148328
rect 380676 148316 380682 148368
rect 358722 146956 358728 147008
rect 358780 146996 358786 147008
rect 363598 146996 363604 147008
rect 358780 146968 363604 146996
rect 358780 146956 358786 146968
rect 363598 146956 363604 146968
rect 363656 146956 363662 147008
rect 355962 146888 355968 146940
rect 356020 146928 356026 146940
rect 364978 146928 364984 146940
rect 356020 146900 364984 146928
rect 356020 146888 356026 146900
rect 364978 146888 364984 146900
rect 365036 146888 365042 146940
rect 355410 146752 355416 146804
rect 355468 146792 355474 146804
rect 362862 146792 362868 146804
rect 355468 146764 362868 146792
rect 355468 146752 355474 146764
rect 362862 146752 362868 146764
rect 362920 146752 362926 146804
rect 352650 146684 352656 146736
rect 352708 146724 352714 146736
rect 365898 146724 365904 146736
rect 352708 146696 365904 146724
rect 352708 146684 352714 146696
rect 365898 146684 365904 146696
rect 365956 146684 365962 146736
rect 358170 146616 358176 146668
rect 358228 146656 358234 146668
rect 388990 146656 388996 146668
rect 358228 146628 388996 146656
rect 358228 146616 358234 146628
rect 388990 146616 388996 146628
rect 389048 146616 389054 146668
rect 358262 146548 358268 146600
rect 358320 146588 358326 146600
rect 390186 146588 390192 146600
rect 358320 146560 390192 146588
rect 358320 146548 358326 146560
rect 390186 146548 390192 146560
rect 390244 146548 390250 146600
rect 359550 146480 359556 146532
rect 359608 146520 359614 146532
rect 392578 146520 392584 146532
rect 359608 146492 392584 146520
rect 359608 146480 359614 146492
rect 392578 146480 392584 146492
rect 392636 146480 392642 146532
rect 355594 146412 355600 146464
rect 355652 146452 355658 146464
rect 362770 146452 362776 146464
rect 355652 146424 362776 146452
rect 355652 146412 355658 146424
rect 362770 146412 362776 146424
rect 362828 146412 362834 146464
rect 362862 146412 362868 146464
rect 362920 146452 362926 146464
rect 391382 146452 391388 146464
rect 362920 146424 391388 146452
rect 362920 146412 362926 146424
rect 391382 146412 391388 146424
rect 391440 146412 391446 146464
rect 359458 146344 359464 146396
rect 359516 146384 359522 146396
rect 397362 146384 397368 146396
rect 359516 146356 397368 146384
rect 359516 146344 359522 146356
rect 397362 146344 397368 146356
rect 397420 146344 397426 146396
rect 355870 146276 355876 146328
rect 355928 146316 355934 146328
rect 362678 146316 362684 146328
rect 355928 146288 362684 146316
rect 355928 146276 355934 146288
rect 362678 146276 362684 146288
rect 362736 146276 362742 146328
rect 362770 146276 362776 146328
rect 362828 146316 362834 146328
rect 398558 146316 398564 146328
rect 362828 146288 398564 146316
rect 362828 146276 362834 146288
rect 398558 146276 398564 146288
rect 398616 146276 398622 146328
rect 358354 144440 358360 144492
rect 358412 144480 358418 144492
rect 386414 144480 386420 144492
rect 358412 144452 386420 144480
rect 358412 144440 358418 144452
rect 386414 144440 386420 144452
rect 386472 144440 386478 144492
rect 358630 144372 358636 144424
rect 358688 144412 358694 144424
rect 385126 144412 385132 144424
rect 358688 144384 385132 144412
rect 358688 144372 358694 144384
rect 385126 144372 385132 144384
rect 385184 144372 385190 144424
rect 359642 144304 359648 144356
rect 359700 144344 359706 144356
rect 407758 144344 407764 144356
rect 359700 144316 407764 144344
rect 359700 144304 359706 144316
rect 407758 144304 407764 144316
rect 407816 144304 407822 144356
rect 358446 144236 358452 144288
rect 358504 144276 358510 144288
rect 387702 144276 387708 144288
rect 358504 144248 387708 144276
rect 358504 144236 358510 144248
rect 387702 144236 387708 144248
rect 387760 144236 387766 144288
rect 238386 122000 238392 122052
rect 238444 122040 238450 122052
rect 239950 122040 239956 122052
rect 238444 122012 239956 122040
rect 238444 122000 238450 122012
rect 239950 122000 239956 122012
rect 240008 122000 240014 122052
rect 235810 120640 235816 120692
rect 235868 120680 235874 120692
rect 283190 120680 283196 120692
rect 235868 120652 283196 120680
rect 235868 120640 235874 120652
rect 283190 120640 283196 120652
rect 283248 120640 283254 120692
rect 235902 120572 235908 120624
rect 235960 120612 235966 120624
rect 355594 120612 355600 120624
rect 235960 120584 355600 120612
rect 235960 120572 235966 120584
rect 355594 120572 355600 120584
rect 355652 120572 355658 120624
rect 279970 120504 279976 120556
rect 280028 120544 280034 120556
rect 290090 120544 290096 120556
rect 280028 120516 290096 120544
rect 280028 120504 280034 120516
rect 290090 120504 290096 120516
rect 290148 120504 290154 120556
rect 50246 120028 50252 120080
rect 50304 120068 50310 120080
rect 63494 120068 63500 120080
rect 50304 120040 63500 120068
rect 50304 120028 50310 120040
rect 63494 120028 63500 120040
rect 63552 120028 63558 120080
rect 126974 120028 126980 120080
rect 127032 120068 127038 120080
rect 128998 120068 129004 120080
rect 127032 120040 129004 120068
rect 127032 120028 127038 120040
rect 128998 120028 129004 120040
rect 129056 120028 129062 120080
rect 129918 120028 129924 120080
rect 129976 120068 129982 120080
rect 358630 120068 358636 120080
rect 129976 120040 358636 120068
rect 129976 120028 129982 120040
rect 358630 120028 358636 120040
rect 358688 120028 358694 120080
rect 50614 119960 50620 120012
rect 50672 120000 50678 120012
rect 61470 120000 61476 120012
rect 50672 119972 61476 120000
rect 50672 119960 50678 119972
rect 61470 119960 61476 119972
rect 61528 119960 61534 120012
rect 127618 119960 127624 120012
rect 127676 120000 127682 120012
rect 350074 120000 350080 120012
rect 127676 119972 350080 120000
rect 127676 119960 127682 119972
rect 350074 119960 350080 119972
rect 350132 119960 350138 120012
rect 127526 119892 127532 119944
rect 127584 119932 127590 119944
rect 289814 119932 289820 119944
rect 127584 119904 289820 119932
rect 127584 119892 127590 119904
rect 289814 119892 289820 119904
rect 289872 119892 289878 119944
rect 127802 119824 127808 119876
rect 127860 119864 127866 119876
rect 284294 119864 284300 119876
rect 127860 119836 284300 119864
rect 127860 119824 127866 119836
rect 284294 119824 284300 119836
rect 284352 119824 284358 119876
rect 128078 119756 128084 119808
rect 128136 119796 128142 119808
rect 283098 119796 283104 119808
rect 128136 119768 283104 119796
rect 128136 119756 128142 119768
rect 283098 119756 283104 119768
rect 283156 119756 283162 119808
rect 127802 119688 127808 119740
rect 127860 119728 127866 119740
rect 129918 119728 129924 119740
rect 127860 119700 129924 119728
rect 127860 119688 127866 119700
rect 129918 119688 129924 119700
rect 129976 119688 129982 119740
rect 238570 119688 238576 119740
rect 238628 119728 238634 119740
rect 358538 119728 358544 119740
rect 238628 119700 358544 119728
rect 238628 119688 238634 119700
rect 358538 119688 358544 119700
rect 358596 119688 358602 119740
rect 238294 119620 238300 119672
rect 238352 119660 238358 119672
rect 318150 119660 318156 119672
rect 238352 119632 318156 119660
rect 238352 119620 238358 119632
rect 318150 119620 318156 119632
rect 318208 119620 318214 119672
rect 235810 119552 235816 119604
rect 235868 119592 235874 119604
rect 284570 119592 284576 119604
rect 235868 119564 284576 119592
rect 235868 119552 235874 119564
rect 284570 119552 284576 119564
rect 284628 119552 284634 119604
rect 235902 119484 235908 119536
rect 235960 119524 235966 119536
rect 284386 119524 284392 119536
rect 235960 119496 284392 119524
rect 235960 119484 235966 119496
rect 284386 119484 284392 119496
rect 284444 119484 284450 119536
rect 238570 119416 238576 119468
rect 238628 119456 238634 119468
rect 284478 119456 284484 119468
rect 238628 119428 284484 119456
rect 238628 119416 238634 119428
rect 284478 119416 284484 119428
rect 284536 119416 284542 119468
rect 49510 118600 49516 118652
rect 49568 118640 49574 118652
rect 72326 118640 72332 118652
rect 49568 118612 72332 118640
rect 49568 118600 49574 118612
rect 72326 118600 72332 118612
rect 72384 118600 72390 118652
rect 109034 118600 109040 118652
rect 109092 118640 109098 118652
rect 125686 118640 125692 118652
rect 109092 118612 125692 118640
rect 109092 118600 109098 118612
rect 125686 118600 125692 118612
rect 125744 118600 125750 118652
rect 234614 118600 234620 118652
rect 234672 118640 234678 118652
rect 245746 118640 245752 118652
rect 234672 118612 245752 118640
rect 234672 118600 234678 118612
rect 245746 118600 245752 118612
rect 245804 118600 245810 118652
rect 247034 118600 247040 118652
rect 247092 118640 247098 118652
rect 250070 118640 250076 118652
rect 247092 118612 250076 118640
rect 247092 118600 247098 118612
rect 250070 118600 250076 118612
rect 250128 118600 250134 118652
rect 50522 118532 50528 118584
rect 50580 118572 50586 118584
rect 84562 118572 84568 118584
rect 50580 118544 84568 118572
rect 50580 118532 50586 118544
rect 84562 118532 84568 118544
rect 84620 118532 84626 118584
rect 114278 118532 114284 118584
rect 114336 118572 114342 118584
rect 125778 118572 125784 118584
rect 114336 118544 125784 118572
rect 114336 118532 114342 118544
rect 125778 118532 125784 118544
rect 125836 118572 125842 118584
rect 126882 118572 126888 118584
rect 125836 118544 126888 118572
rect 125836 118532 125842 118544
rect 126882 118532 126888 118544
rect 126940 118532 126946 118584
rect 237558 118532 237564 118584
rect 237616 118572 237622 118584
rect 246574 118572 246580 118584
rect 237616 118544 246580 118572
rect 237616 118532 237622 118544
rect 246574 118532 246580 118544
rect 246632 118532 246638 118584
rect 48038 118464 48044 118516
rect 48096 118504 48102 118516
rect 81066 118504 81072 118516
rect 48096 118476 81072 118504
rect 48096 118464 48102 118476
rect 81066 118464 81072 118476
rect 81124 118464 81130 118516
rect 116026 118464 116032 118516
rect 116084 118504 116090 118516
rect 129090 118504 129096 118516
rect 116084 118476 129096 118504
rect 116084 118464 116090 118476
rect 129090 118464 129096 118476
rect 129148 118464 129154 118516
rect 132494 118504 132500 118516
rect 132466 118464 132500 118504
rect 132552 118504 132558 118516
rect 359550 118504 359556 118516
rect 132552 118476 359556 118504
rect 132552 118464 132558 118476
rect 359550 118464 359556 118476
rect 359608 118464 359614 118516
rect 49602 118396 49608 118448
rect 49660 118436 49666 118448
rect 79318 118436 79324 118448
rect 49660 118408 79324 118436
rect 49660 118396 49666 118408
rect 79318 118396 79324 118408
rect 79376 118396 79382 118448
rect 102042 118396 102048 118448
rect 102100 118436 102106 118448
rect 117682 118436 117688 118448
rect 102100 118408 117688 118436
rect 102100 118396 102106 118408
rect 117682 118396 117688 118408
rect 117740 118396 117746 118448
rect 117774 118396 117780 118448
rect 117832 118436 117838 118448
rect 124398 118436 124404 118448
rect 117832 118408 124404 118436
rect 117832 118396 117838 118408
rect 124398 118396 124404 118408
rect 124456 118436 124462 118448
rect 125226 118436 125232 118448
rect 124456 118408 125232 118436
rect 124456 118396 124462 118408
rect 125226 118396 125232 118408
rect 125284 118396 125290 118448
rect 47946 118328 47952 118380
rect 48004 118368 48010 118380
rect 77570 118368 77576 118380
rect 48004 118340 77576 118368
rect 48004 118328 48010 118340
rect 77570 118328 77576 118340
rect 77628 118328 77634 118380
rect 103790 118328 103796 118380
rect 103848 118368 103854 118380
rect 128538 118368 128544 118380
rect 103848 118340 128544 118368
rect 103848 118328 103854 118340
rect 128538 118328 128544 118340
rect 128596 118328 128602 118380
rect 48130 118260 48136 118312
rect 48188 118300 48194 118312
rect 75822 118300 75828 118312
rect 48188 118272 75828 118300
rect 48188 118260 48194 118272
rect 75822 118260 75828 118272
rect 75880 118260 75886 118312
rect 107286 118260 107292 118312
rect 107344 118300 107350 118312
rect 132466 118300 132494 118464
rect 239950 118396 239956 118448
rect 240008 118436 240014 118448
rect 349798 118436 349804 118448
rect 240008 118408 349804 118436
rect 240008 118396 240014 118408
rect 349798 118396 349804 118408
rect 349856 118396 349862 118448
rect 238202 118328 238208 118380
rect 238260 118368 238266 118380
rect 359642 118368 359648 118380
rect 238260 118340 359648 118368
rect 238260 118328 238266 118340
rect 359642 118328 359648 118340
rect 359700 118328 359706 118380
rect 107344 118272 132494 118300
rect 107344 118260 107350 118272
rect 238478 118260 238484 118312
rect 238536 118300 238542 118312
rect 349982 118300 349988 118312
rect 238536 118272 349988 118300
rect 238536 118260 238542 118272
rect 349982 118260 349988 118272
rect 350040 118260 350046 118312
rect 105538 118192 105544 118244
rect 105596 118232 105602 118244
rect 129826 118232 129832 118244
rect 105596 118204 129832 118232
rect 105596 118192 105602 118204
rect 129826 118192 129832 118204
rect 129884 118192 129890 118244
rect 238018 118192 238024 118244
rect 238076 118232 238082 118244
rect 349890 118232 349896 118244
rect 238076 118204 349896 118232
rect 238076 118192 238082 118204
rect 349890 118192 349896 118204
rect 349948 118192 349954 118244
rect 110782 118124 110788 118176
rect 110840 118164 110846 118176
rect 132586 118164 132592 118176
rect 110840 118136 132592 118164
rect 110840 118124 110846 118136
rect 132586 118124 132592 118136
rect 132644 118124 132650 118176
rect 237374 118124 237380 118176
rect 237432 118164 237438 118176
rect 248966 118164 248972 118176
rect 237432 118136 248972 118164
rect 237432 118124 237438 118136
rect 248966 118124 248972 118136
rect 249024 118124 249030 118176
rect 264974 118124 264980 118176
rect 265032 118164 265038 118176
rect 294046 118164 294052 118176
rect 265032 118136 294052 118164
rect 265032 118124 265038 118136
rect 294046 118124 294052 118136
rect 294104 118124 294110 118176
rect 112530 118056 112536 118108
rect 112588 118096 112594 118108
rect 131206 118096 131212 118108
rect 112588 118068 131212 118096
rect 112588 118056 112594 118068
rect 131206 118056 131212 118068
rect 131264 118096 131270 118108
rect 131482 118096 131488 118108
rect 131264 118068 131488 118096
rect 131264 118056 131270 118068
rect 131482 118056 131488 118068
rect 131540 118056 131546 118108
rect 237466 118056 237472 118108
rect 237524 118096 237530 118108
rect 247678 118096 247684 118108
rect 237524 118068 247684 118096
rect 237524 118056 237530 118068
rect 247678 118056 247684 118068
rect 247736 118056 247742 118108
rect 271782 118056 271788 118108
rect 271840 118096 271846 118108
rect 292666 118096 292672 118108
rect 271840 118068 292672 118096
rect 271840 118056 271846 118068
rect 292666 118056 292672 118068
rect 292724 118056 292730 118108
rect 117682 117988 117688 118040
rect 117740 118028 117746 118040
rect 124214 118028 124220 118040
rect 117740 118000 124220 118028
rect 117740 117988 117746 118000
rect 124214 117988 124220 118000
rect 124272 118028 124278 118040
rect 125502 118028 125508 118040
rect 124272 118000 125508 118028
rect 124272 117988 124278 118000
rect 125502 117988 125508 118000
rect 125560 117988 125566 118040
rect 126882 117988 126888 118040
rect 126940 118028 126946 118040
rect 359458 118028 359464 118040
rect 126940 118000 359464 118028
rect 126940 117988 126946 118000
rect 359458 117988 359464 118000
rect 359516 117988 359522 118040
rect 61838 117920 61844 117972
rect 61896 117960 61902 117972
rect 360654 117960 360660 117972
rect 61896 117932 360660 117960
rect 61896 117920 61902 117932
rect 360654 117920 360660 117932
rect 360712 117920 360718 117972
rect 89806 117852 89812 117904
rect 89864 117892 89870 117904
rect 124858 117892 124864 117904
rect 89864 117864 124864 117892
rect 89864 117852 89870 117864
rect 124858 117852 124864 117864
rect 124916 117852 124922 117904
rect 91554 117784 91560 117836
rect 91612 117824 91618 117836
rect 125594 117824 125600 117836
rect 91612 117796 125600 117824
rect 91612 117784 91618 117796
rect 125594 117784 125600 117796
rect 125652 117784 125658 117836
rect 121454 117716 121460 117768
rect 121512 117756 121518 117768
rect 244274 117756 244280 117768
rect 121512 117728 244280 117756
rect 121512 117716 121518 117728
rect 244274 117716 244280 117728
rect 244332 117716 244338 117768
rect 45370 117240 45376 117292
rect 45428 117280 45434 117292
rect 67542 117280 67548 117292
rect 45428 117252 67548 117280
rect 45428 117240 45434 117252
rect 67542 117240 67548 117252
rect 67600 117240 67606 117292
rect 128538 117240 128544 117292
rect 128596 117280 128602 117292
rect 358262 117280 358268 117292
rect 128596 117252 358268 117280
rect 128596 117240 128602 117252
rect 358262 117240 358268 117252
rect 358320 117240 358326 117292
rect 46750 117172 46756 117224
rect 46808 117212 46814 117224
rect 65334 117212 65340 117224
rect 46808 117184 65340 117212
rect 46808 117172 46814 117184
rect 65334 117172 65340 117184
rect 65392 117212 65398 117224
rect 66162 117212 66168 117224
rect 65392 117184 66168 117212
rect 65392 117172 65398 117184
rect 66162 117172 66168 117184
rect 66220 117172 66226 117224
rect 107562 117172 107568 117224
rect 107620 117212 107626 117224
rect 129734 117212 129740 117224
rect 107620 117184 129740 117212
rect 107620 117172 107626 117184
rect 129734 117172 129740 117184
rect 129792 117212 129798 117224
rect 358354 117212 358360 117224
rect 129792 117184 358360 117212
rect 129792 117172 129798 117184
rect 358354 117172 358360 117184
rect 358412 117172 358418 117224
rect 106182 117104 106188 117156
rect 106240 117144 106246 117156
rect 131114 117144 131120 117156
rect 106240 117116 131120 117144
rect 106240 117104 106246 117116
rect 131114 117104 131120 117116
rect 131172 117144 131178 117156
rect 358446 117144 358452 117156
rect 131172 117116 358452 117144
rect 131172 117104 131178 117116
rect 358446 117104 358452 117116
rect 358504 117104 358510 117156
rect 191742 117036 191748 117088
rect 191800 117076 191806 117088
rect 355410 117076 355416 117088
rect 191800 117048 355416 117076
rect 191800 117036 191806 117048
rect 355410 117036 355416 117048
rect 355468 117036 355474 117088
rect 212442 116968 212448 117020
rect 212500 117008 212506 117020
rect 358170 117008 358176 117020
rect 212500 116980 358176 117008
rect 212500 116968 212506 116980
rect 358170 116968 358176 116980
rect 358228 116968 358234 117020
rect 241422 116900 241428 116952
rect 241480 116940 241486 116952
rect 352650 116940 352656 116952
rect 241480 116912 352656 116940
rect 241480 116900 241486 116912
rect 352650 116900 352656 116912
rect 352708 116900 352714 116952
rect 66162 115880 66168 115932
rect 66220 115920 66226 115932
rect 295978 115920 295984 115932
rect 66220 115892 295984 115920
rect 66220 115880 66226 115892
rect 295978 115880 295984 115892
rect 296036 115880 296042 115932
rect 67542 115812 67548 115864
rect 67600 115852 67606 115864
rect 297358 115852 297364 115864
rect 67600 115824 297364 115852
rect 67600 115812 67606 115824
rect 297358 115812 297364 115824
rect 297416 115812 297422 115864
rect 234614 115744 234620 115796
rect 234672 115784 234678 115796
rect 355962 115784 355968 115796
rect 234672 115756 355968 115784
rect 234672 115744 234678 115756
rect 355962 115744 355968 115756
rect 356020 115784 356026 115796
rect 358078 115784 358084 115796
rect 356020 115756 358084 115784
rect 356020 115744 356026 115756
rect 358078 115744 358084 115756
rect 358136 115744 358142 115796
rect 252462 114452 252468 114504
rect 252520 114492 252526 114504
rect 289998 114492 290004 114504
rect 252520 114464 290004 114492
rect 252520 114452 252526 114464
rect 289998 114452 290004 114464
rect 290056 114452 290062 114504
rect 360654 88952 360660 89004
rect 360712 88992 360718 89004
rect 537478 88992 537484 89004
rect 360712 88964 537484 88992
rect 360712 88952 360718 88964
rect 537478 88952 537484 88964
rect 537536 88952 537542 89004
rect 73062 87252 73068 87304
rect 73120 87292 73126 87304
rect 91738 87292 91744 87304
rect 73120 87264 91744 87292
rect 73120 87252 73126 87264
rect 91738 87252 91744 87264
rect 91796 87252 91802 87304
rect 74442 87184 74448 87236
rect 74500 87224 74506 87236
rect 86310 87224 86316 87236
rect 74500 87196 86316 87224
rect 74500 87184 74506 87196
rect 86310 87184 86316 87196
rect 86368 87184 86374 87236
rect 76466 87116 76472 87168
rect 76524 87156 76530 87168
rect 90542 87156 90548 87168
rect 76524 87128 90548 87156
rect 76524 87116 76530 87128
rect 90542 87116 90548 87128
rect 90600 87116 90606 87168
rect 84010 87048 84016 87100
rect 84068 87088 84074 87100
rect 98730 87088 98736 87100
rect 84068 87060 98736 87088
rect 84068 87048 84074 87060
rect 98730 87048 98736 87060
rect 98788 87048 98794 87100
rect 358078 86912 358084 86964
rect 358136 86952 358142 86964
rect 580166 86952 580172 86964
rect 358136 86924 580172 86952
rect 358136 86912 358142 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 86310 69640 86316 69692
rect 86368 69680 86374 69692
rect 350442 69680 350448 69692
rect 86368 69652 350448 69680
rect 86368 69640 86374 69652
rect 350442 69640 350448 69652
rect 350500 69640 350506 69692
rect 91738 54476 91744 54528
rect 91796 54516 91802 54528
rect 346946 54516 346952 54528
rect 91796 54488 346952 54516
rect 91796 54476 91802 54488
rect 346946 54476 346952 54488
rect 347004 54476 347010 54528
rect 90542 50328 90548 50380
rect 90600 50368 90606 50380
rect 354030 50368 354036 50380
rect 90600 50340 354036 50368
rect 90600 50328 90606 50340
rect 354030 50328 354036 50340
rect 354088 50328 354094 50380
rect 537478 46860 537484 46912
rect 537536 46900 537542 46912
rect 580166 46900 580172 46912
rect 537536 46872 580172 46900
rect 537536 46860 537542 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 98730 10276 98736 10328
rect 98788 10316 98794 10328
rect 371694 10316 371700 10328
rect 98788 10288 371700 10316
rect 98788 10276 98794 10288
rect 371694 10276 371700 10288
rect 371752 10276 371758 10328
rect 331858 6808 331864 6860
rect 331916 6848 331922 6860
rect 580166 6848 580172 6860
rect 331916 6820 580172 6848
rect 331916 6808 331922 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 271782 4088 271788 4140
rect 271840 4128 271846 4140
rect 292574 4128 292580 4140
rect 271840 4100 292580 4128
rect 271840 4088 271846 4100
rect 292574 4088 292580 4100
rect 292632 4088 292638 4140
rect 446398 3408 446404 3460
rect 446456 3448 446462 3460
rect 583386 3448 583392 3460
rect 446456 3420 583392 3448
rect 446456 3408 446462 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 442902 2796 442908 2848
rect 442960 2836 442966 2848
rect 580994 2836 581000 2848
rect 442960 2808 581000 2836
rect 442960 2796 442966 2808
rect 580994 2796 581000 2808
rect 581052 2796 581058 2848
<< via1 >>
rect 300124 700340 300176 700392
rect 322204 700340 322256 700392
rect 527180 700340 527232 700392
rect 543924 700340 543976 700392
rect 170312 700272 170364 700324
rect 324964 700272 325016 700324
rect 332508 700272 332560 700324
rect 340144 700272 340196 700324
rect 509148 700272 509200 700324
rect 559656 700272 559708 700324
rect 40500 699660 40552 699712
rect 41420 699660 41472 699712
rect 86224 699660 86276 699712
rect 478512 699660 478564 699712
rect 479524 699660 479576 699712
rect 255964 687896 256016 687948
rect 267648 687896 267700 687948
rect 283840 687148 283892 687200
rect 286324 687148 286376 687200
rect 348792 686468 348844 686520
rect 358084 686468 358136 686520
rect 3424 683136 3476 683188
rect 26148 683136 26200 683188
rect 87604 683136 87656 683188
rect 358084 680348 358136 680400
rect 360844 680348 360896 680400
rect 340144 677492 340196 677544
rect 345664 677492 345716 677544
rect 250444 674772 250496 674824
rect 255964 674772 256016 674824
rect 360844 672052 360896 672104
rect 366364 672052 366416 672104
rect 242440 661716 242492 661768
rect 250444 661716 250496 661768
rect 345664 660288 345716 660340
rect 355968 660288 356020 660340
rect 45468 658248 45520 658300
rect 105452 658248 105504 658300
rect 106188 658248 106240 658300
rect 489736 657976 489788 658028
rect 501788 657976 501840 658028
rect 486976 657840 487028 657892
rect 496268 657840 496320 657892
rect 364984 657772 365036 657824
rect 491024 657772 491076 657824
rect 322204 657704 322256 657756
rect 490472 657704 490524 657756
rect 491208 657704 491260 657756
rect 494704 657704 494756 657756
rect 510068 657704 510120 657756
rect 286324 657636 286376 657688
rect 294604 657636 294656 657688
rect 324964 657636 325016 657688
rect 516140 657636 516192 657688
rect 106188 657568 106240 657620
rect 518348 657568 518400 657620
rect 86224 657500 86276 657552
rect 519728 657500 519780 657552
rect 144184 657432 144236 657484
rect 525248 657432 525300 657484
rect 532148 657432 532200 657484
rect 546592 657432 546644 657484
rect 488448 657364 488500 657416
rect 493508 657364 493560 657416
rect 509148 657364 509200 657416
rect 540980 657364 541032 657416
rect 58624 657296 58676 657348
rect 522488 657296 522540 657348
rect 526628 657296 526680 657348
rect 544108 657296 544160 657348
rect 488264 657228 488316 657280
rect 503168 657228 503220 657280
rect 530768 657228 530820 657280
rect 544200 657228 544252 657280
rect 490564 657160 490616 657212
rect 491116 657160 491168 657212
rect 511448 657160 511500 657212
rect 528008 657160 528060 657212
rect 544016 657160 544068 657212
rect 491208 657092 491260 657144
rect 514208 657092 514260 657144
rect 529388 657092 529440 657144
rect 545396 657092 545448 657144
rect 485688 657024 485740 657076
rect 494888 657024 494940 657076
rect 490380 656956 490432 657008
rect 491024 656956 491076 657008
rect 512828 657024 512880 657076
rect 534908 657024 534960 657076
rect 547972 657024 548024 657076
rect 533528 656956 533580 657008
rect 545488 656956 545540 657008
rect 516140 656888 516192 656940
rect 516968 656888 517020 656940
rect 540336 656888 540388 656940
rect 366364 656820 366416 656872
rect 371884 656820 371936 656872
rect 505928 655596 505980 655648
rect 540428 655596 540480 655648
rect 504548 655528 504600 655580
rect 543740 655528 543792 655580
rect 239404 655460 239456 655512
rect 242440 655460 242492 655512
rect 355968 654780 356020 654832
rect 366364 654780 366416 654832
rect 486884 654576 486936 654628
rect 498660 654576 498712 654628
rect 156604 654508 156656 654560
rect 523500 654508 523552 654560
rect 489644 654440 489696 654492
rect 491852 654440 491904 654492
rect 497372 654440 497424 654492
rect 485596 654372 485648 654424
rect 488448 654236 488500 654288
rect 490656 654236 490708 654288
rect 178040 654100 178092 654152
rect 368388 654100 368440 654152
rect 371884 651992 371936 652044
rect 377404 651992 377456 652044
rect 213828 651516 213880 651568
rect 361948 651516 362000 651568
rect 233148 651448 233200 651500
rect 464344 651448 464396 651500
rect 227720 651380 227772 651432
rect 483664 651380 483716 651432
rect 231768 650292 231820 650344
rect 374368 650292 374420 650344
rect 226340 650224 226392 650276
rect 375656 650224 375708 650276
rect 214564 650156 214616 650208
rect 374828 650156 374880 650208
rect 212448 650088 212500 650140
rect 374552 650088 374604 650140
rect 186320 650020 186372 650072
rect 374736 650020 374788 650072
rect 543556 650020 543608 650072
rect 549260 650020 549312 650072
rect 205640 648796 205692 648848
rect 467104 648796 467156 648848
rect 224224 648728 224276 648780
rect 486424 648728 486476 648780
rect 199660 648660 199712 648712
rect 469956 648660 470008 648712
rect 198740 648592 198792 648644
rect 472624 648592 472676 648644
rect 234620 647504 234672 647556
rect 354220 647504 354272 647556
rect 217508 647436 217560 647488
rect 472900 647436 472952 647488
rect 203340 647368 203392 647420
rect 471244 647368 471296 647420
rect 176568 647300 176620 647352
rect 478144 647300 478196 647352
rect 54392 647232 54444 647284
rect 372252 647232 372304 647284
rect 366364 647164 366416 647216
rect 371884 647164 371936 647216
rect 294604 646484 294656 646536
rect 304264 646484 304316 646536
rect 115848 646144 115900 646196
rect 325884 646144 325936 646196
rect 240692 646076 240744 646128
rect 462964 646076 463016 646128
rect 209780 646008 209832 646060
rect 483756 646008 483808 646060
rect 204628 645940 204680 645992
rect 482376 645940 482428 645992
rect 146208 645804 146260 645856
rect 151084 645872 151136 645924
rect 176568 645872 176620 645924
rect 479708 645872 479760 645924
rect 177304 644784 177356 644836
rect 393228 644784 393280 644836
rect 218796 644716 218848 644768
rect 464436 644716 464488 644768
rect 230388 644648 230440 644700
rect 476764 644648 476816 644700
rect 138664 644580 138716 644632
rect 390192 644580 390244 644632
rect 131120 644512 131172 644564
rect 384120 644512 384172 644564
rect 91100 644444 91152 644496
rect 351644 644444 351696 644496
rect 186964 643696 187016 643748
rect 239404 643696 239456 643748
rect 176752 643492 176804 643544
rect 389180 643492 389232 643544
rect 126888 643424 126940 643476
rect 338764 643424 338816 643476
rect 176660 643356 176712 643408
rect 419540 643356 419592 643408
rect 124128 643288 124180 643340
rect 365812 643288 365864 643340
rect 377404 643288 377456 643340
rect 380532 643288 380584 643340
rect 221740 643220 221792 643272
rect 464528 643220 464580 643272
rect 225512 643152 225564 643204
rect 483848 643152 483900 643204
rect 198464 643084 198516 643136
rect 472716 643084 472768 643136
rect 294052 642404 294104 642456
rect 340052 642404 340104 642456
rect 293960 642336 294012 642388
rect 382096 642336 382148 642388
rect 178040 642268 178092 642320
rect 346492 642268 346544 642320
rect 153936 642200 153988 642252
rect 375564 642200 375616 642252
rect 216588 642132 216640 642184
rect 464620 642132 464672 642184
rect 202420 642064 202472 642116
rect 482560 642064 482612 642116
rect 177948 641996 178000 642048
rect 458824 641996 458876 642048
rect 59268 641928 59320 641980
rect 350356 641928 350408 641980
rect 144276 641860 144328 641912
rect 146208 641860 146260 641912
rect 183100 641860 183152 641912
rect 475476 641860 475528 641912
rect 59268 641792 59320 641844
rect 352932 641792 352984 641844
rect 57888 641724 57940 641776
rect 355508 641724 355560 641776
rect 380532 640976 380584 641028
rect 387800 640976 387852 641028
rect 251088 640908 251140 640960
rect 320732 640908 320784 640960
rect 249708 640840 249760 640892
rect 322020 640840 322072 640892
rect 127624 640772 127676 640824
rect 331036 640772 331088 640824
rect 222936 640704 222988 640756
rect 465816 640704 465868 640756
rect 195888 640636 195940 640688
rect 472808 640636 472860 640688
rect 59268 640568 59320 640620
rect 337476 640568 337528 640620
rect 177580 640500 177632 640552
rect 458916 640500 458968 640552
rect 56508 640432 56560 640484
rect 349068 640432 349120 640484
rect 193128 640364 193180 640416
rect 489368 640364 489420 640416
rect 148324 640296 148376 640348
rect 149704 640296 149756 640348
rect 177948 640296 178000 640348
rect 489184 640296 489236 640348
rect 109040 639548 109092 639600
rect 309140 639548 309192 639600
rect 88984 639480 89036 639532
rect 318156 639480 318208 639532
rect 220360 639412 220412 639464
rect 471520 639412 471572 639464
rect 154488 639344 154540 639396
rect 421564 639344 421616 639396
rect 88248 639276 88300 639328
rect 385132 639276 385184 639328
rect 106188 639208 106240 639260
rect 403348 639208 403400 639260
rect 107568 639140 107620 639192
rect 405372 639140 405424 639192
rect 66168 639072 66220 639124
rect 376852 639072 376904 639124
rect 88800 639004 88852 639056
rect 403624 639004 403676 639056
rect 91008 638936 91060 638988
rect 406384 638936 406436 638988
rect 234528 638324 234580 638376
rect 291844 638324 291896 638376
rect 137284 638256 137336 638308
rect 313004 638256 313056 638308
rect 227720 638188 227772 638240
rect 414664 638188 414716 638240
rect 252468 638120 252520 638172
rect 475660 638120 475712 638172
rect 86868 638052 86920 638104
rect 319444 638052 319496 638104
rect 129740 637984 129792 638036
rect 400864 637984 400916 638036
rect 118700 637916 118752 637968
rect 397276 637916 397328 637968
rect 179052 637848 179104 637900
rect 463240 637848 463292 637900
rect 81440 637780 81492 637832
rect 367100 637780 367152 637832
rect 110420 637712 110472 637764
rect 399300 637712 399352 637764
rect 102140 637644 102192 637696
rect 400312 637644 400364 637696
rect 82820 637576 82872 637628
rect 395344 637576 395396 637628
rect 73160 637508 73212 637560
rect 176752 637508 176804 637560
rect 108304 637440 108356 637492
rect 177304 637440 177356 637492
rect 117964 637372 118016 637424
rect 176660 637372 176712 637424
rect 117228 637304 117280 637356
rect 138664 637304 138716 637356
rect 128360 636964 128412 637016
rect 292028 636964 292080 637016
rect 128452 636896 128504 636948
rect 297456 636896 297508 636948
rect 125508 636828 125560 636880
rect 297364 636828 297416 636880
rect 121460 636760 121512 636812
rect 306564 636760 306616 636812
rect 245568 636692 245620 636744
rect 456156 636692 456208 636744
rect 242808 636624 242860 636676
rect 459008 636624 459060 636676
rect 236000 636556 236052 636608
rect 456064 636556 456116 636608
rect 246948 636488 247000 636540
rect 486516 636488 486568 636540
rect 240048 636420 240100 636472
rect 489460 636420 489512 636472
rect 179328 636352 179380 636404
rect 453304 636352 453356 636404
rect 191748 636284 191800 636336
rect 472992 636284 473044 636336
rect 179972 636216 180024 636268
rect 485136 636216 485188 636268
rect 387800 636148 387852 636200
rect 391388 636148 391440 636200
rect 38568 635468 38620 635520
rect 72976 635468 73028 635520
rect 156696 635468 156748 635520
rect 375380 635468 375432 635520
rect 247592 635400 247644 635452
rect 471428 635400 471480 635452
rect 92480 635332 92532 635384
rect 342628 635332 342680 635384
rect 99380 635264 99432 635316
rect 391296 635264 391348 635316
rect 95148 635196 95200 635248
rect 386144 635196 386196 635248
rect 109132 635128 109184 635180
rect 412456 635128 412508 635180
rect 104808 635060 104860 635112
rect 410524 635060 410576 635112
rect 98092 634992 98144 635044
rect 409420 634992 409472 635044
rect 96528 634924 96580 634976
rect 407764 634924 407816 634976
rect 101680 634856 101732 634908
rect 414480 634856 414532 634908
rect 97816 634788 97868 634840
rect 411444 634788 411496 634840
rect 151084 634448 151136 634500
rect 376760 634448 376812 634500
rect 171968 634380 172020 634432
rect 186964 634380 187016 634432
rect 371884 634380 371936 634432
rect 387708 634380 387760 634432
rect 3424 632068 3476 632120
rect 31576 632068 31628 632120
rect 58624 632000 58676 632052
rect 146944 630640 146996 630692
rect 148324 630640 148376 630692
rect 387708 627172 387760 627224
rect 400772 627172 400824 627224
rect 377220 622412 377272 622464
rect 380164 622412 380216 622464
rect 391388 621664 391440 621716
rect 398104 621664 398156 621716
rect 400772 621664 400824 621716
rect 406476 621664 406528 621716
rect 144920 620984 144972 621036
rect 146944 620984 146996 621036
rect 282184 619624 282236 619676
rect 298008 619624 298060 619676
rect 142804 619556 142856 619608
rect 144920 619556 144972 619608
rect 289084 618264 289136 618316
rect 298008 618264 298060 618316
rect 260104 617516 260156 617568
rect 282184 617516 282236 617568
rect 540428 617516 540480 617568
rect 580172 617516 580224 617568
rect 293224 616836 293276 616888
rect 298008 616836 298060 616888
rect 542912 616836 542964 616888
rect 545580 616836 545632 616888
rect 159364 613368 159416 613420
rect 171968 613368 172020 613420
rect 292028 612688 292080 612740
rect 298008 612688 298060 612740
rect 398104 612008 398156 612060
rect 410616 612008 410668 612060
rect 142896 611328 142948 611380
rect 144276 611328 144328 611380
rect 175188 610648 175240 610700
rect 179052 610648 179104 610700
rect 406476 610580 406528 610632
rect 420184 610580 420236 610632
rect 377036 604528 377088 604580
rect 379796 604528 379848 604580
rect 378048 604460 378100 604512
rect 386420 604460 386472 604512
rect 410616 604460 410668 604512
rect 413284 604460 413336 604512
rect 540336 604460 540388 604512
rect 541440 604460 541492 604512
rect 286324 603100 286376 603152
rect 297916 603100 297968 603152
rect 136088 602352 136140 602404
rect 159364 602352 159416 602404
rect 539232 600992 539284 601044
rect 540980 600992 541032 601044
rect 488356 600244 488408 600296
rect 498844 600244 498896 600296
rect 537576 600244 537628 600296
rect 540428 600244 540480 600296
rect 488264 600176 488316 600228
rect 510344 600176 510396 600228
rect 488448 600108 488500 600160
rect 524052 600108 524104 600160
rect 489644 600040 489696 600092
rect 525892 600040 525944 600092
rect 462320 599972 462372 600024
rect 499396 599972 499448 600024
rect 485688 599904 485740 599956
rect 529204 599904 529256 599956
rect 486976 599836 487028 599888
rect 530584 599836 530636 599888
rect 485596 599768 485648 599820
rect 531412 599768 531464 599820
rect 486884 599700 486936 599752
rect 532792 599700 532844 599752
rect 489736 599632 489788 599684
rect 535736 599632 535788 599684
rect 413652 599564 413704 599616
rect 499304 599564 499356 599616
rect 519728 598884 519780 598936
rect 532976 598884 533028 598936
rect 515588 598816 515640 598868
rect 529848 598816 529900 598868
rect 518348 598748 518400 598800
rect 531320 598748 531372 598800
rect 512828 598272 512880 598324
rect 527272 598272 527324 598324
rect 493508 598204 493560 598256
rect 498936 598204 498988 598256
rect 514208 598204 514260 598256
rect 535552 598204 535604 598256
rect 492128 598136 492180 598188
rect 498752 598136 498804 598188
rect 531228 598136 531280 598188
rect 536288 598136 536340 598188
rect 496268 598068 496320 598120
rect 499120 598068 499172 598120
rect 518164 597524 518216 597576
rect 521108 597524 521160 597576
rect 536104 597524 536156 597576
rect 539048 597524 539100 597576
rect 378048 593444 378100 593496
rect 385040 593444 385092 593496
rect 377956 593376 378008 593428
rect 386604 593376 386656 593428
rect 141424 593308 141476 593360
rect 142896 593308 142948 593360
rect 378048 592288 378100 592340
rect 382832 592288 382884 592340
rect 378048 592084 378100 592136
rect 385316 592084 385368 592136
rect 45284 592016 45336 592068
rect 57520 592016 57572 592068
rect 134524 591336 134576 591388
rect 136088 591336 136140 591388
rect 378048 590656 378100 590708
rect 385224 590656 385276 590708
rect 378048 589908 378100 589960
rect 385408 589908 385460 589960
rect 420184 589908 420236 589960
rect 428464 589908 428516 589960
rect 378048 589296 378100 589348
rect 382464 589296 382516 589348
rect 378048 587936 378100 587988
rect 382280 587936 382332 587988
rect 376944 587868 376996 587920
rect 379612 587868 379664 587920
rect 413284 587800 413336 587852
rect 416136 587800 416188 587852
rect 377772 586916 377824 586968
rect 381268 586916 381320 586968
rect 162308 586576 162360 586628
rect 170864 586576 170916 586628
rect 378048 586576 378100 586628
rect 383752 586576 383804 586628
rect 141516 586508 141568 586560
rect 142804 586508 142856 586560
rect 162584 586508 162636 586560
rect 169484 586508 169536 586560
rect 378048 585148 378100 585200
rect 382372 585148 382424 585200
rect 258724 584400 258776 584452
rect 258908 584400 258960 584452
rect 378048 584128 378100 584180
rect 383660 584128 383712 584180
rect 140044 583720 140096 583772
rect 141516 583720 141568 583772
rect 378048 583720 378100 583772
rect 382740 583720 382792 583772
rect 378048 582496 378100 582548
rect 382648 582496 382700 582548
rect 378048 582360 378100 582412
rect 382556 582360 382608 582412
rect 490380 581612 490432 581664
rect 493324 581612 493376 581664
rect 377864 581000 377916 581052
rect 381452 581000 381504 581052
rect 165068 579776 165120 579828
rect 173716 579776 173768 579828
rect 377588 579708 377640 579760
rect 380900 579708 380952 579760
rect 3424 579640 3476 579692
rect 41512 579640 41564 579692
rect 377128 579640 377180 579692
rect 379888 579640 379940 579692
rect 377864 578280 377916 578332
rect 381360 578280 381412 578332
rect 377036 578212 377088 578264
rect 379704 578212 379756 578264
rect 377128 575492 377180 575544
rect 379980 575492 380032 575544
rect 416136 575492 416188 575544
rect 419632 575492 419684 575544
rect 378048 572704 378100 572756
rect 386696 572704 386748 572756
rect 378048 571888 378100 571940
rect 383844 571888 383896 571940
rect 378048 571344 378100 571396
rect 383936 571344 383988 571396
rect 428464 571276 428516 571328
rect 433984 571276 434036 571328
rect 419632 570596 419684 570648
rect 429200 570596 429252 570648
rect 169300 569780 169352 569832
rect 171140 569780 171192 569832
rect 164976 569644 165028 569696
rect 172428 569644 172480 569696
rect 377036 568556 377088 568608
rect 379520 568556 379572 568608
rect 493324 568488 493376 568540
rect 496084 568488 496136 568540
rect 377772 567808 377824 567860
rect 381176 567808 381228 567860
rect 429200 567196 429252 567248
rect 432052 567196 432104 567248
rect 543740 564340 543792 564392
rect 580172 564340 580224 564392
rect 537760 563660 537812 563712
rect 543740 563660 543792 563712
rect 169116 562300 169168 562352
rect 170128 562300 170180 562352
rect 178408 562300 178460 562352
rect 178684 562300 178736 562352
rect 432052 562300 432104 562352
rect 444288 562300 444340 562352
rect 140044 561824 140096 561876
rect 135168 561620 135220 561672
rect 259184 561688 259236 561740
rect 299664 561688 299716 561740
rect 299572 561144 299624 561196
rect 254492 561008 254544 561060
rect 299572 560940 299624 560992
rect 294052 560872 294104 560924
rect 297916 560872 297968 560924
rect 525984 560940 526036 560992
rect 254676 560668 254728 560720
rect 293960 560668 294012 560720
rect 253572 560600 253624 560652
rect 254860 560600 254912 560652
rect 254400 560532 254452 560584
rect 300584 560532 300636 560584
rect 253480 560464 253532 560516
rect 300676 560464 300728 560516
rect 246580 560396 246632 560448
rect 299572 560396 299624 560448
rect 169208 560328 169260 560380
rect 172244 560328 172296 560380
rect 319352 560600 319404 560652
rect 59544 560260 59596 560312
rect 60740 560260 60792 560312
rect 179052 560260 179104 560312
rect 245476 560260 245528 560312
rect 287796 560260 287848 560312
rect 45284 560192 45336 560244
rect 162492 560192 162544 560244
rect 168012 560192 168064 560244
rect 172336 560192 172388 560244
rect 175740 560192 175792 560244
rect 297640 560192 297692 560244
rect 315396 560192 315448 560244
rect 318340 560124 318392 560176
rect 165528 560056 165580 560108
rect 173716 560056 173768 560108
rect 299664 560056 299716 560108
rect 306380 560056 306432 560108
rect 216680 559580 216732 559632
rect 357808 559580 357860 559632
rect 444288 559580 444340 559632
rect 459100 559580 459152 559632
rect 91192 559512 91244 559564
rect 141424 559512 141476 559564
rect 177212 559512 177264 559564
rect 514852 559512 514904 559564
rect 169852 559444 169904 559496
rect 367928 559444 367980 559496
rect 169760 559376 169812 559428
rect 368940 559376 368992 559428
rect 233700 559308 233752 559360
rect 500224 559308 500276 559360
rect 60648 559240 60700 559292
rect 369952 559240 370004 559292
rect 57244 559172 57296 559224
rect 370964 559172 371016 559224
rect 56968 559104 57020 559156
rect 371976 559104 372028 559156
rect 57520 559036 57572 559088
rect 373264 559036 373316 559088
rect 166540 558968 166592 559020
rect 512000 558968 512052 559020
rect 166816 558900 166868 558952
rect 520740 558900 520792 558952
rect 53840 558832 53892 558884
rect 372344 558832 372396 558884
rect 53932 558764 53984 558816
rect 367284 558764 367336 558816
rect 56048 558696 56100 558748
rect 361212 558696 361264 558748
rect 59268 558628 59320 558680
rect 357164 558628 357216 558680
rect 63592 558560 63644 558612
rect 355140 558560 355192 558612
rect 89628 558492 89680 558544
rect 91192 558492 91244 558544
rect 231768 558492 231820 558544
rect 297548 558492 297600 558544
rect 300676 558492 300728 558544
rect 314660 558492 314712 558544
rect 245660 558424 245712 558476
rect 199936 558288 199988 558340
rect 251824 558288 251876 558340
rect 293960 558424 294012 558476
rect 353116 558424 353168 558476
rect 293316 558356 293368 558408
rect 303528 558356 303580 558408
rect 294052 558288 294104 558340
rect 300584 558288 300636 558340
rect 521936 558288 521988 558340
rect 177304 558220 177356 558272
rect 503996 558220 504048 558272
rect 104900 558152 104952 558204
rect 135168 558152 135220 558204
rect 177580 558152 177632 558204
rect 512184 558152 512236 558204
rect 252468 557676 252520 557728
rect 346676 557676 346728 557728
rect 37096 557540 37148 557592
rect 41512 557608 41564 557660
rect 180708 557608 180760 557660
rect 524696 557608 524748 557660
rect 180616 557540 180668 557592
rect 537024 557540 537076 557592
rect 53840 557472 53892 557524
rect 297732 557472 297784 557524
rect 156604 557404 156656 557456
rect 202052 557404 202104 557456
rect 254400 557404 254452 557456
rect 128268 557064 128320 557116
rect 174912 557064 174964 557116
rect 57612 556996 57664 557048
rect 170864 556996 170916 557048
rect 250444 556996 250496 557048
rect 293224 556996 293276 557048
rect 137744 556928 137796 556980
rect 259000 556928 259052 556980
rect 280804 556928 280856 556980
rect 378784 556928 378836 556980
rect 91100 556860 91152 556912
rect 104900 556860 104952 556912
rect 137928 556860 137980 556912
rect 331956 556860 332008 556912
rect 61384 556792 61436 556844
rect 375932 556792 375984 556844
rect 255044 556656 255096 556708
rect 260104 556656 260156 556708
rect 230388 556588 230440 556640
rect 448888 556588 448940 556640
rect 227720 556520 227772 556572
rect 449900 556520 449952 556572
rect 179420 556452 179472 556504
rect 450912 556452 450964 556504
rect 178132 556384 178184 556436
rect 452936 556384 452988 556436
rect 178040 556316 178092 556368
rect 453948 556316 454000 556368
rect 137468 556248 137520 556300
rect 137744 556248 137796 556300
rect 175832 556248 175884 556300
rect 454960 556248 455012 556300
rect 56048 556180 56100 556232
rect 56508 556180 56560 556232
rect 86868 556180 86920 556232
rect 89628 556180 89680 556232
rect 175188 556180 175240 556232
rect 509976 556180 510028 556232
rect 137192 556112 137244 556164
rect 137468 556112 137520 556164
rect 56508 556044 56560 556096
rect 379980 556044 380032 556096
rect 137192 555976 137244 556028
rect 376944 555976 376996 556028
rect 53840 555908 53892 555960
rect 381452 555908 381504 555960
rect 137468 555568 137520 555620
rect 271144 555568 271196 555620
rect 137652 555500 137704 555552
rect 347136 555500 347188 555552
rect 175832 555432 175884 555484
rect 507860 555432 507912 555484
rect 247040 555160 247092 555212
rect 434720 555160 434772 555212
rect 226340 555092 226392 555144
rect 460020 555092 460072 555144
rect 179420 555024 179472 555076
rect 473176 555024 473228 555076
rect 178040 554956 178092 555008
rect 475200 554956 475252 555008
rect 220176 554888 220228 554940
rect 523040 554888 523092 554940
rect 185768 554820 185820 554872
rect 543740 554820 543792 554872
rect 78588 554752 78640 554804
rect 86868 554752 86920 554804
rect 151360 554752 151412 554804
rect 510160 554752 510212 554804
rect 57336 554684 57388 554736
rect 375840 554684 375892 554736
rect 60004 554616 60056 554668
rect 323768 554616 323820 554668
rect 173808 554548 173860 554600
rect 378692 554548 378744 554600
rect 178040 554480 178092 554532
rect 376852 554480 376904 554532
rect 230388 554412 230440 554464
rect 376760 554412 376812 554464
rect 240048 554344 240100 554396
rect 376024 554344 376076 554396
rect 192944 554276 192996 554328
rect 253572 554276 253624 554328
rect 256700 554276 256752 554328
rect 376116 554276 376168 554328
rect 179052 554140 179104 554192
rect 477224 554140 477276 554192
rect 174636 554072 174688 554124
rect 482284 554072 482336 554124
rect 57612 554004 57664 554056
rect 375748 554004 375800 554056
rect 496084 553528 496136 553580
rect 497464 553528 497516 553580
rect 219164 553460 219216 553512
rect 523132 553460 523184 553512
rect 177948 553392 178000 553444
rect 513564 553392 513616 553444
rect 59176 553324 59228 553376
rect 379796 553324 379848 553376
rect 56508 553256 56560 553308
rect 369308 553256 369360 553308
rect 98644 553188 98696 553240
rect 378140 553188 378192 553240
rect 97908 553120 97960 553172
rect 326804 553120 326856 553172
rect 60832 553052 60884 553104
rect 156696 553052 156748 553104
rect 191748 553052 191800 553104
rect 253020 553052 253072 553104
rect 170772 552780 170824 552832
rect 463056 552780 463108 552832
rect 208124 552712 208176 552764
rect 530032 552712 530084 552764
rect 184848 552644 184900 552696
rect 519360 552644 519412 552696
rect 253204 552236 253256 552288
rect 343640 552236 343692 552288
rect 88984 552168 89036 552220
rect 91100 552168 91152 552220
rect 249708 552168 249760 552220
rect 344652 552168 344704 552220
rect 114468 552100 114520 552152
rect 351736 552100 351788 552152
rect 234620 552032 234672 552084
rect 512920 552032 512972 552084
rect 81440 551964 81492 552016
rect 346032 551964 346084 552016
rect 433984 551964 434036 552016
rect 436100 551964 436152 552016
rect 490472 551964 490524 552016
rect 493324 551964 493376 552016
rect 111800 551896 111852 551948
rect 374644 551896 374696 551948
rect 172428 551828 172480 551880
rect 381268 551828 381320 551880
rect 118700 551760 118752 551812
rect 317696 551760 317748 551812
rect 175832 551692 175884 551744
rect 297456 551692 297508 551744
rect 204076 551420 204128 551472
rect 507400 551420 507452 551472
rect 174268 551352 174320 551404
rect 486332 551352 486384 551404
rect 189908 551284 189960 551336
rect 508044 551284 508096 551336
rect 236000 550808 236052 550860
rect 360844 550808 360896 550860
rect 224224 550740 224276 550792
rect 518900 550740 518952 550792
rect 180064 550672 180116 550724
rect 526260 550672 526312 550724
rect 163504 550604 163556 550656
rect 509240 550604 509292 550656
rect 75920 550536 75972 550588
rect 78588 550536 78640 550588
rect 80060 550536 80112 550588
rect 344008 550536 344060 550588
rect 99380 550468 99432 550520
rect 327816 550468 327868 550520
rect 92480 550400 92532 550452
rect 153936 550400 153988 550452
rect 173808 550400 173860 550452
rect 379520 550400 379572 550452
rect 168380 550332 168432 550384
rect 304540 550332 304592 550384
rect 137744 550128 137796 550180
rect 418804 550128 418856 550180
rect 226064 550060 226116 550112
rect 510804 550060 510856 550112
rect 210884 549992 210936 550044
rect 506572 549992 506624 550044
rect 60096 549924 60148 549976
rect 378600 549924 378652 549976
rect 79600 549856 79652 549908
rect 88984 549856 89036 549908
rect 177396 549856 177448 549908
rect 514944 549856 514996 549908
rect 131120 549380 131172 549432
rect 372988 549380 373040 549432
rect 221188 549312 221240 549364
rect 524420 549312 524472 549364
rect 176568 549244 176620 549296
rect 537116 549244 537168 549296
rect 79324 549176 79376 549228
rect 380164 549176 380216 549228
rect 110420 549108 110472 549160
rect 354128 549108 354180 549160
rect 178040 549040 178092 549092
rect 381360 549040 381412 549092
rect 169760 548972 169812 549024
rect 348056 548972 348108 549024
rect 175188 548904 175240 548956
rect 254492 548904 254544 548956
rect 459100 548768 459152 548820
rect 466920 548768 466972 548820
rect 198740 548700 198792 548752
rect 505376 548700 505428 548752
rect 211896 548632 211948 548684
rect 526076 548632 526128 548684
rect 200764 548564 200816 548616
rect 523500 548564 523552 548616
rect 166356 548496 166408 548548
rect 492404 548496 492456 548548
rect 436100 548360 436152 548412
rect 441620 548360 441672 548412
rect 227720 548088 227772 548140
rect 462044 548088 462096 548140
rect 253204 548020 253256 548072
rect 500316 548020 500368 548072
rect 161480 547952 161532 548004
rect 506480 547952 506532 548004
rect 93676 547884 93728 547936
rect 520648 547884 520700 547936
rect 67548 547816 67600 547868
rect 347044 547816 347096 547868
rect 88984 547748 89036 547800
rect 151084 547748 151136 547800
rect 166172 547748 166224 547800
rect 383936 547748 383988 547800
rect 136548 547680 136600 547732
rect 320732 547680 320784 547732
rect 172060 547272 172112 547324
rect 467012 547272 467064 547324
rect 185584 547204 185636 547256
rect 508136 547204 508188 547256
rect 182548 547136 182600 547188
rect 527364 547136 527416 547188
rect 231768 546796 231820 546848
rect 365904 546796 365956 546848
rect 246304 546728 246356 546780
rect 496084 546728 496136 546780
rect 187792 546660 187844 546712
rect 503720 546660 503772 546712
rect 175648 546592 175700 546644
rect 531320 546592 531372 546644
rect 175188 546524 175240 546576
rect 540336 546524 540388 546576
rect 77300 546456 77352 546508
rect 79600 546456 79652 546508
rect 90640 546456 90692 546508
rect 520556 546456 520608 546508
rect 56508 546388 56560 546440
rect 359188 546388 359240 546440
rect 75828 546320 75880 546372
rect 350080 546320 350132 546372
rect 86868 546252 86920 546304
rect 335912 546252 335964 546304
rect 126888 546184 126940 546236
rect 313648 546184 313700 546236
rect 224132 546116 224184 546168
rect 307576 546116 307628 546168
rect 299664 546048 299716 546100
rect 538404 546048 538456 546100
rect 289636 545980 289688 546032
rect 541532 545980 541584 546032
rect 173440 545912 173492 545964
rect 483296 545912 483348 545964
rect 196716 545844 196768 545896
rect 528928 545844 528980 545896
rect 183560 545776 183612 545828
rect 528836 545776 528888 545828
rect 179604 545708 179656 545760
rect 538496 545708 538548 545760
rect 192852 545164 192904 545216
rect 253940 545164 253992 545216
rect 441620 545164 441672 545216
rect 444380 545164 444432 545216
rect 493324 545164 493376 545216
rect 496176 545164 496228 545216
rect 218152 545096 218204 545148
rect 522580 545096 522632 545148
rect 75828 545028 75880 545080
rect 364248 545028 364300 545080
rect 88248 544960 88300 545012
rect 329840 544960 329892 545012
rect 131120 544892 131172 544944
rect 324780 544892 324832 544944
rect 169760 544824 169812 544876
rect 253480 544824 253532 544876
rect 216680 544756 216732 544808
rect 250444 544756 250496 544808
rect 251824 544620 251876 544672
rect 545672 544620 545724 544672
rect 170588 544552 170640 544604
rect 465080 544552 465132 544604
rect 202788 544484 202840 544536
rect 506664 544484 506716 544536
rect 209872 544416 209924 544468
rect 530216 544416 530268 544468
rect 177488 544348 177540 544400
rect 515128 544348 515180 544400
rect 252468 543872 252520 543924
rect 526168 543872 526220 543924
rect 181720 543804 181772 543856
rect 539876 543804 539928 543856
rect 72424 543668 72476 543720
rect 75736 543736 75788 543788
rect 94688 543736 94740 543788
rect 523408 543736 523460 543788
rect 128728 543668 128780 543720
rect 134524 543668 134576 543720
rect 127624 543600 127676 543652
rect 362224 543668 362276 543720
rect 208400 543600 208452 543652
rect 360200 543600 360252 543652
rect 240048 543532 240100 543584
rect 325792 543532 325844 543584
rect 244280 543464 244332 543516
rect 259184 543464 259236 543516
rect 160744 543260 160796 543312
rect 255044 543260 255096 543312
rect 191104 543192 191156 543244
rect 382832 543192 382884 543244
rect 194692 543124 194744 543176
rect 503812 543124 503864 543176
rect 173256 543056 173308 543108
rect 485320 543056 485372 543108
rect 193680 542988 193732 543040
rect 532976 542988 533028 543040
rect 466920 542920 466972 542972
rect 470140 542920 470192 542972
rect 299204 542580 299256 542632
rect 511172 542580 511224 542632
rect 242808 542512 242860 542564
rect 503904 542512 503956 542564
rect 172612 542444 172664 542496
rect 517704 542444 517756 542496
rect 91652 542376 91704 542428
rect 517796 542376 517848 542428
rect 82820 542308 82872 542360
rect 363236 542308 363288 542360
rect 178040 542240 178092 542292
rect 383844 542240 383896 542292
rect 128360 542172 128412 542224
rect 328828 542172 328880 542224
rect 129740 542104 129792 542156
rect 316684 542104 316736 542156
rect 291844 541832 291896 541884
rect 536288 541832 536340 541884
rect 171968 541764 172020 541816
rect 468116 541764 468168 541816
rect 179696 541696 179748 541748
rect 517980 541696 518032 541748
rect 181536 541628 181588 541680
rect 527456 541628 527508 541680
rect 236000 541220 236052 541272
rect 506756 541220 506808 541272
rect 172428 541152 172480 541204
rect 516600 541152 516652 541204
rect 178684 541084 178736 541136
rect 524512 541084 524564 541136
rect 148324 541016 148376 541068
rect 506480 541016 506532 541068
rect 92664 540948 92716 541000
rect 516508 540948 516560 541000
rect 91100 540880 91152 540932
rect 368296 540880 368348 540932
rect 444380 540880 444432 540932
rect 447232 540880 447284 540932
rect 107568 540812 107620 540864
rect 345020 540812 345072 540864
rect 218060 540744 218112 540796
rect 374736 540744 374788 540796
rect 169760 540676 169812 540728
rect 254860 540676 254912 540728
rect 187608 540336 187660 540388
rect 508228 540336 508280 540388
rect 177672 540268 177724 540320
rect 515312 540268 515364 540320
rect 73160 540200 73212 540252
rect 77300 540200 77352 540252
rect 92020 540200 92072 540252
rect 144184 540200 144236 540252
rect 190644 540200 190696 540252
rect 530124 540200 530176 540252
rect 244280 539928 244332 539980
rect 254768 539928 254820 539980
rect 247040 539860 247092 539912
rect 354772 539860 354824 539912
rect 175188 539792 175240 539844
rect 466092 539792 466144 539844
rect 217140 539724 217192 539776
rect 521660 539724 521712 539776
rect 158444 539656 158496 539708
rect 500408 539656 500460 539708
rect 88616 539588 88668 539640
rect 521660 539588 521712 539640
rect 60832 539520 60884 539572
rect 371332 539520 371384 539572
rect 86868 539452 86920 539504
rect 352104 539452 352156 539504
rect 100760 539384 100812 539436
rect 340972 539384 341024 539436
rect 124864 539316 124916 539368
rect 128728 539316 128780 539368
rect 136548 539316 136600 539368
rect 331864 539316 331916 539368
rect 222108 539248 222160 539300
rect 386604 539248 386656 539300
rect 206836 538908 206888 538960
rect 506848 538908 506900 538960
rect 174544 538840 174596 538892
rect 479248 538840 479300 538892
rect 104808 538500 104860 538552
rect 375012 538500 375064 538552
rect 225512 538432 225564 538484
rect 501052 538432 501104 538484
rect 156420 538364 156472 538416
rect 496268 538364 496320 538416
rect 170588 538296 170640 538348
rect 516140 538296 516192 538348
rect 179696 538228 179748 538280
rect 536840 538228 536892 538280
rect 85488 538160 85540 538212
rect 373356 538160 373408 538212
rect 117228 538092 117280 538144
rect 330852 538092 330904 538144
rect 252468 538024 252520 538076
rect 311624 538024 311676 538076
rect 205824 537616 205876 537668
rect 505560 537616 505612 537668
rect 175924 537548 175976 537600
rect 478328 537548 478380 537600
rect 172888 537480 172940 537532
rect 488356 537480 488408 537532
rect 109040 537140 109092 537192
rect 376024 537140 376076 537192
rect 213092 537072 213144 537124
rect 518440 537072 518492 537124
rect 180708 537004 180760 537056
rect 511540 537004 511592 537056
rect 190828 536936 190880 536988
rect 543832 536936 543884 536988
rect 72424 536868 72476 536920
rect 166908 536868 166960 536920
rect 527640 536868 527692 536920
rect 66260 536732 66312 536784
rect 69020 536732 69072 536784
rect 73160 536800 73212 536852
rect 84568 536800 84620 536852
rect 520464 536800 520516 536852
rect 89720 536732 89772 536784
rect 370320 536732 370372 536784
rect 109040 536664 109092 536716
rect 342996 536664 343048 536716
rect 117228 536596 117280 536648
rect 297364 536596 297416 536648
rect 168380 536528 168432 536580
rect 301504 536528 301556 536580
rect 479708 536392 479760 536444
rect 530400 536392 530452 536444
rect 447232 536324 447284 536376
rect 456800 536324 456852 536376
rect 472992 536324 473044 536376
rect 537300 536324 537352 536376
rect 456156 536256 456208 536308
rect 535828 536256 535880 536308
rect 174728 536188 174780 536240
rect 457996 536188 458048 536240
rect 459008 536188 459060 536240
rect 524604 536188 524656 536240
rect 171784 536120 171836 536172
rect 490380 536120 490432 536172
rect 186596 536052 186648 536104
rect 508320 536052 508372 536104
rect 299388 535780 299440 535832
rect 353760 535780 353812 535832
rect 175924 535712 175976 535764
rect 355784 535712 355836 535764
rect 216128 535644 216180 535696
rect 520280 535644 520332 535696
rect 241336 535576 241388 535628
rect 545764 535576 545816 535628
rect 191840 535508 191892 535560
rect 535368 535508 535420 535560
rect 85580 535440 85632 535492
rect 519176 535440 519228 535492
rect 100760 535372 100812 535424
rect 358176 535372 358228 535424
rect 169760 535304 169812 535356
rect 334900 535304 334952 535356
rect 251088 535236 251140 535288
rect 309600 535236 309652 535288
rect 60740 534896 60792 534948
rect 348700 534896 348752 534948
rect 470140 534896 470192 534948
rect 475844 534896 475896 534948
rect 212908 534828 212960 534880
rect 506940 534828 506992 534880
rect 197728 534760 197780 534812
rect 505744 534760 505796 534812
rect 63592 534692 63644 534744
rect 69020 534692 69072 534744
rect 177764 534692 177816 534744
rect 513840 534692 513892 534744
rect 108304 534352 108356 534404
rect 377036 534352 377088 534404
rect 211068 534284 211120 534336
rect 497556 534284 497608 534336
rect 209044 534216 209096 534268
rect 527180 534216 527232 534268
rect 154396 534148 154448 534200
rect 499580 534148 499632 534200
rect 157984 534080 158036 534132
rect 160744 534080 160796 534132
rect 167552 534080 167604 534132
rect 517060 534080 517112 534132
rect 106188 534012 106240 534064
rect 366272 534012 366324 534064
rect 115848 533944 115900 533996
rect 332876 533944 332928 533996
rect 175924 533876 175976 533928
rect 339960 533876 340012 533928
rect 223488 533808 223540 533860
rect 337936 533808 337988 533860
rect 195704 533536 195756 533588
rect 505652 533536 505704 533588
rect 171876 533468 171928 533520
rect 484308 533468 484360 533520
rect 489368 533468 489420 533520
rect 544476 533468 544528 533520
rect 188620 533400 188672 533452
rect 505468 533400 505520 533452
rect 177120 533332 177172 533384
rect 513748 533332 513800 533384
rect 485044 533060 485096 533112
rect 513932 533060 513984 533112
rect 251824 532992 251876 533044
rect 509792 532992 509844 533044
rect 215116 532924 215168 532976
rect 519084 532924 519136 532976
rect 194876 532856 194928 532908
rect 538220 532856 538272 532908
rect 169576 532788 169628 532840
rect 514760 532788 514812 532840
rect 83556 532720 83608 532772
rect 518992 532720 519044 532772
rect 59636 532652 59688 532704
rect 376300 532652 376352 532704
rect 215300 532584 215352 532636
rect 374552 532584 374604 532636
rect 175464 532108 175516 532160
rect 487344 532108 487396 532160
rect 57336 532040 57388 532092
rect 376208 532040 376260 532092
rect 57428 531972 57480 532024
rect 378324 531972 378376 532024
rect 254860 531700 254912 531752
rect 521660 531700 521712 531752
rect 214104 531632 214156 531684
rect 517612 531632 517664 531684
rect 198924 531564 198976 531616
rect 507860 531564 507912 531616
rect 208032 531496 208084 531548
rect 525800 531496 525852 531548
rect 168564 531428 168616 531480
rect 499580 531428 499632 531480
rect 177948 531360 178000 531412
rect 512828 531360 512880 531412
rect 62856 531224 62908 531276
rect 66168 531292 66220 531344
rect 184756 531292 184808 531344
rect 529848 531360 529900 531412
rect 166172 531224 166224 531276
rect 374828 531224 374880 531276
rect 178224 531156 178276 531208
rect 287796 531156 287848 531208
rect 178132 531088 178184 531140
rect 280804 531088 280856 531140
rect 489460 531088 489512 531140
rect 538588 531088 538640 531140
rect 476764 531020 476816 531072
rect 534908 531020 534960 531072
rect 178868 530952 178920 531004
rect 472900 530952 472952 531004
rect 533252 530952 533304 531004
rect 471520 530884 471572 530936
rect 533344 530884 533396 530936
rect 464528 530816 464580 530868
rect 530676 530816 530728 530868
rect 178868 530748 178920 530800
rect 464344 530748 464396 530800
rect 531688 530748 531740 530800
rect 465816 530680 465868 530732
rect 534724 530680 534776 530732
rect 464620 530612 464672 530664
rect 534540 530612 534592 530664
rect 137284 530544 137336 530596
rect 342904 530544 342956 530596
rect 464436 530544 464488 530596
rect 534632 530544 534684 530596
rect 164148 530476 164200 530528
rect 313188 530476 313240 530528
rect 175924 530408 175976 530460
rect 374092 530408 374144 530460
rect 256700 530340 256752 530392
rect 469128 530340 469180 530392
rect 60188 530272 60240 530324
rect 285772 530272 285824 530324
rect 521752 530272 521804 530324
rect 178040 530204 178092 530256
rect 470140 530204 470192 530256
rect 62764 530136 62816 530188
rect 138204 530136 138256 530188
rect 173808 530136 173860 530188
rect 472164 530136 472216 530188
rect 140228 530068 140280 530120
rect 212080 530068 212132 530120
rect 516232 530068 516284 530120
rect 60280 530000 60332 530052
rect 147312 530000 147364 530052
rect 195888 530000 195940 530052
rect 541072 530000 541124 530052
rect 53748 529932 53800 529984
rect 144276 529932 144328 529984
rect 183744 529932 183796 529984
rect 540980 529932 541032 529984
rect 177856 529864 177908 529916
rect 500960 529864 501012 529916
rect 96528 529796 96580 529848
rect 382740 529796 382792 529848
rect 95148 529728 95200 529780
rect 333888 529728 333940 529780
rect 95056 529660 95108 529712
rect 321744 529660 321796 529712
rect 285680 529592 285732 529644
rect 379888 529592 379940 529644
rect 456800 529524 456852 529576
rect 501880 529524 501932 529576
rect 458824 529456 458876 529508
rect 531596 529456 531648 529508
rect 213920 529388 213972 529440
rect 511080 529388 511132 529440
rect 173164 529320 173216 529372
rect 481272 529320 481324 529372
rect 486516 529320 486568 529372
rect 527548 529320 527600 529372
rect 177028 529252 177080 529304
rect 509792 529252 509844 529304
rect 61108 529184 61160 529236
rect 61568 529184 61620 529236
rect 96896 529184 96948 529236
rect 436008 529184 436060 529236
rect 458916 529184 458968 529236
rect 536012 529184 536064 529236
rect 299388 528776 299440 528828
rect 364892 528776 364944 528828
rect 210056 528708 210108 528760
rect 510252 528708 510304 528760
rect 174636 528640 174688 528692
rect 505928 528640 505980 528692
rect 25964 528572 26016 528624
rect 105820 528572 105872 528624
rect 155408 528572 155460 528624
rect 500960 528572 501012 528624
rect 121460 528504 121512 528556
rect 385408 528504 385460 528556
rect 125508 528436 125560 528488
rect 289084 528436 289136 528488
rect 55128 528368 55180 528420
rect 137836 528368 137888 528420
rect 475844 528368 475896 528420
rect 488540 528368 488592 528420
rect 125416 528300 125468 528352
rect 157984 528300 158036 528352
rect 483756 528300 483808 528352
rect 520924 528300 520976 528352
rect 299296 528232 299348 528284
rect 502892 528232 502944 528284
rect 133328 528164 133380 528216
rect 342628 528164 342680 528216
rect 486424 528164 486476 528216
rect 524972 528164 525024 528216
rect 162216 528096 162268 528148
rect 430580 528096 430632 528148
rect 483664 528096 483716 528148
rect 529020 528096 529072 528148
rect 232136 528028 232188 528080
rect 502156 528028 502208 528080
rect 229100 527960 229152 528012
rect 508504 527960 508556 528012
rect 60832 527892 60884 527944
rect 124864 527892 124916 527944
rect 159364 527892 159416 527944
rect 442724 527892 442776 527944
rect 463240 527892 463292 527944
rect 523316 527892 523368 527944
rect 31760 527824 31812 527876
rect 32772 527824 32824 527876
rect 91744 527824 91796 527876
rect 120080 527824 120132 527876
rect 517520 527824 517572 527876
rect 61568 527620 61620 527672
rect 97908 527620 97960 527672
rect 124128 527620 124180 527672
rect 231768 527620 231820 527672
rect 59820 527552 59872 527604
rect 123944 527552 123996 527604
rect 59268 527484 59320 527536
rect 126980 527484 127032 527536
rect 60556 527416 60608 527468
rect 125048 527416 125100 527468
rect 61660 527348 61712 527400
rect 132040 527348 132092 527400
rect 202052 527348 202104 527400
rect 512000 527348 512052 527400
rect 50988 527280 51040 527332
rect 122932 527280 122984 527332
rect 204168 527280 204220 527332
rect 514760 527280 514812 527332
rect 53472 527212 53524 527264
rect 136180 527212 136232 527264
rect 177764 527212 177816 527264
rect 523040 527212 523092 527264
rect 3424 527144 3476 527196
rect 31760 527144 31812 527196
rect 46756 527144 46808 527196
rect 130108 527144 130160 527196
rect 189908 527144 189960 527196
rect 545120 527144 545172 527196
rect 62028 527076 62080 527128
rect 365260 527076 365312 527128
rect 111800 527008 111852 527060
rect 341984 527008 342036 527060
rect 178040 526940 178092 526992
rect 374460 526940 374512 526992
rect 214564 526872 214616 526924
rect 385316 526872 385368 526924
rect 233884 526804 233936 526856
rect 383752 526804 383804 526856
rect 106188 526736 106240 526788
rect 254676 526736 254728 526788
rect 249708 526668 249760 526720
rect 286324 526668 286376 526720
rect 501788 526668 501840 526720
rect 517520 526668 517572 526720
rect 483848 526600 483900 526652
rect 527916 526600 527968 526652
rect 485136 526532 485188 526584
rect 534448 526532 534500 526584
rect 462964 526464 463016 526516
rect 513656 526464 513708 526516
rect 59452 526396 59504 526448
rect 135904 526396 135956 526448
rect 176844 526396 176896 526448
rect 285772 526396 285824 526448
rect 287704 526396 287756 526448
rect 522396 526396 522448 526448
rect 59728 526328 59780 526380
rect 112904 526328 112956 526380
rect 61844 526260 61896 526312
rect 114928 526260 114980 526312
rect 47952 526192 48004 526244
rect 109776 526192 109828 526244
rect 288348 526192 288400 526244
rect 501696 526192 501748 526244
rect 46664 526124 46716 526176
rect 108764 526124 108816 526176
rect 152556 526124 152608 526176
rect 247040 526124 247092 526176
rect 256700 526124 256752 526176
rect 499948 526124 500000 526176
rect 25780 526056 25832 526108
rect 95608 526056 95660 526108
rect 237472 526056 237524 526108
rect 515220 526056 515272 526108
rect 39948 525988 40000 526040
rect 110788 525988 110840 526040
rect 200028 525988 200080 526040
rect 498200 525988 498252 526040
rect 40960 525920 41012 525972
rect 116860 525920 116912 525972
rect 198096 525920 198148 525972
rect 510620 525920 510672 525972
rect 58624 525852 58676 525904
rect 143264 525852 143316 525904
rect 173808 525852 173860 525904
rect 519084 525852 519136 525904
rect 60372 525784 60424 525836
rect 63408 525784 63460 525836
rect 82728 525784 82780 525836
rect 516324 525784 516376 525836
rect 69020 525716 69072 525768
rect 386420 525716 386472 525768
rect 70400 525648 70452 525700
rect 382464 525648 382516 525700
rect 247040 525580 247092 525632
rect 512000 525580 512052 525632
rect 117964 525512 118016 525564
rect 379612 525512 379664 525564
rect 247040 525444 247092 525496
rect 379704 525444 379756 525496
rect 498660 525444 498712 525496
rect 499120 525444 499172 525496
rect 224960 525376 225012 525428
rect 308588 525376 308640 525428
rect 478144 525376 478196 525428
rect 519636 525376 519688 525428
rect 482560 525308 482612 525360
rect 527824 525308 527876 525360
rect 472716 525240 472768 525292
rect 525064 525240 525116 525292
rect 186872 525172 186924 525224
rect 253204 525172 253256 525224
rect 469956 525172 470008 525224
rect 529296 525172 529348 525224
rect 159640 525104 159692 525156
rect 246304 525104 246356 525156
rect 467104 525104 467156 525156
rect 529112 525104 529164 525156
rect 53196 525036 53248 525088
rect 349068 525036 349120 525088
rect 453304 525036 453356 525088
rect 526352 525036 526404 525088
rect 29920 524968 29972 525020
rect 97724 524968 97776 525020
rect 60740 524900 60792 524952
rect 71964 524900 72016 524952
rect 62028 524832 62080 524884
rect 122012 524832 122064 524884
rect 41052 524764 41104 524816
rect 101680 524764 101732 524816
rect 285680 524764 285732 524816
rect 505192 524764 505244 524816
rect 29828 524696 29880 524748
rect 99748 524696 99800 524748
rect 222384 524696 222436 524748
rect 525800 524696 525852 524748
rect 31484 524628 31536 524680
rect 102692 524628 102744 524680
rect 197084 524628 197136 524680
rect 500868 524628 500920 524680
rect 27344 524560 27396 524612
rect 100760 524560 100812 524612
rect 201040 524560 201092 524612
rect 509884 524560 509936 524612
rect 44180 524492 44232 524544
rect 144828 524492 144880 524544
rect 177948 524492 178000 524544
rect 507216 524492 507268 524544
rect 54576 524424 54628 524476
rect 71872 524424 71924 524476
rect 87696 524424 87748 524476
rect 519268 524424 519320 524476
rect 57704 524356 57756 524408
rect 378876 524356 378928 524408
rect 68928 524288 68980 524340
rect 385224 524288 385276 524340
rect 78588 524220 78640 524272
rect 383660 524220 383712 524272
rect 53840 524152 53892 524204
rect 351092 524152 351144 524204
rect 241336 524084 241388 524136
rect 382648 524084 382700 524136
rect 470048 523880 470100 523932
rect 515588 523880 515640 523932
rect 480996 523812 481048 523864
rect 530492 523812 530544 523864
rect 489184 523744 489236 523796
rect 541624 523744 541676 523796
rect 27528 523676 27580 523728
rect 44180 523676 44232 523728
rect 58900 523676 58952 523728
rect 356152 523676 356204 523728
rect 456064 523676 456116 523728
rect 533160 523676 533212 523728
rect 500316 523608 500368 523660
rect 505836 523608 505888 523660
rect 510160 523608 510212 523660
rect 511264 523608 511316 523660
rect 50804 523540 50856 523592
rect 69664 523540 69716 523592
rect 26884 523472 26936 523524
rect 129740 523472 129792 523524
rect 177948 523472 178000 523524
rect 500316 523472 500368 523524
rect 55864 523404 55916 523456
rect 71780 523404 71832 523456
rect 481548 523404 481600 523456
rect 522120 523404 522172 523456
rect 42432 523336 42484 523388
rect 103796 523336 103848 523388
rect 203064 523336 203116 523388
rect 500040 523336 500092 523388
rect 500408 523336 500460 523388
rect 503720 523336 503772 523388
rect 29736 523268 29788 523320
rect 98736 523268 98788 523320
rect 223304 523268 223356 523320
rect 525800 523268 525852 523320
rect 28632 523200 28684 523252
rect 104716 523200 104768 523252
rect 206192 523200 206244 523252
rect 516876 523200 516928 523252
rect 60740 523132 60792 523184
rect 139400 523132 139452 523184
rect 496728 523132 496780 523184
rect 545212 523132 545264 523184
rect 25596 523064 25648 523116
rect 117872 523064 117924 523116
rect 182916 523064 182968 523116
rect 528560 523064 528612 523116
rect 52552 522996 52604 523048
rect 68928 522996 68980 523048
rect 171692 522996 171744 523048
rect 518072 522996 518124 523048
rect 59544 522928 59596 522980
rect 60832 522928 60884 522980
rect 178040 522928 178092 522980
rect 378232 522928 378284 522980
rect 395344 522928 395396 522980
rect 396172 522928 396224 522980
rect 400864 522928 400916 522980
rect 402336 522928 402388 522980
rect 403624 522928 403676 522980
rect 404268 522928 404320 522980
rect 407764 522928 407816 522980
rect 410432 522928 410484 522980
rect 410524 522928 410576 522980
rect 413376 522928 413428 522980
rect 414664 522928 414716 522980
rect 415492 522928 415544 522980
rect 500224 522928 500276 522980
rect 500408 522928 500460 522980
rect 184848 522860 184900 522912
rect 369124 522860 369176 522912
rect 373264 522860 373316 522912
rect 374000 522860 374052 522912
rect 488540 522860 488592 522912
rect 497372 522860 497424 522912
rect 224132 522792 224184 522844
rect 385040 522792 385092 522844
rect 475660 522792 475712 522844
rect 518072 522792 518124 522844
rect 227720 522724 227772 522776
rect 386696 522724 386748 522776
rect 436008 522724 436060 522776
rect 491300 522724 491352 522776
rect 226340 522656 226392 522708
rect 382556 522656 382608 522708
rect 391296 522656 391348 522708
rect 408408 522656 408460 522708
rect 418804 522656 418856 522708
rect 489276 522656 489328 522708
rect 496084 522656 496136 522708
rect 505284 522656 505336 522708
rect 42340 522588 42392 522640
rect 70400 522588 70452 522640
rect 347136 522588 347188 522640
rect 476120 522588 476172 522640
rect 496268 522588 496320 522640
rect 513380 522588 513432 522640
rect 43904 522520 43956 522572
rect 69388 522520 69440 522572
rect 69664 522520 69716 522572
rect 111800 522520 111852 522572
rect 313188 522520 313240 522572
rect 474096 522520 474148 522572
rect 475476 522520 475528 522572
rect 522212 522520 522264 522572
rect 97908 522452 97960 522504
rect 153384 522452 153436 522504
rect 174912 522452 174964 522504
rect 337476 522452 337528 522504
rect 342904 522452 342956 522504
rect 480260 522452 480312 522504
rect 482376 522452 482428 522504
rect 516784 522452 516836 522504
rect 52828 522384 52880 522436
rect 59820 522384 59872 522436
rect 68928 522384 68980 522436
rect 118884 522384 118936 522436
rect 129740 522384 129792 522436
rect 142160 522384 142212 522436
rect 150348 522384 150400 522436
rect 251824 522384 251876 522436
rect 271144 522384 271196 522436
rect 435732 522384 435784 522436
rect 472808 522384 472860 522436
rect 521016 522384 521068 522436
rect 52460 522316 52512 522368
rect 60740 522316 60792 522368
rect 89628 522316 89680 522368
rect 254860 522316 254912 522368
rect 259000 522316 259052 522368
rect 456984 522316 457036 522368
rect 472624 522316 472676 522368
rect 526536 522316 526588 522368
rect 27160 522248 27212 522300
rect 41420 522248 41472 522300
rect 43812 522248 43864 522300
rect 67364 522248 67416 522300
rect 71780 522248 71832 522300
rect 139216 522248 139268 522300
rect 139400 522248 139452 522300
rect 157340 522248 157392 522300
rect 170864 522248 170916 522300
rect 378048 522248 378100 522300
rect 380900 522248 380952 522300
rect 44088 522180 44140 522232
rect 68376 522180 68428 522232
rect 253204 522180 253256 522232
rect 381176 522180 381228 522232
rect 45284 522112 45336 522164
rect 77484 522112 77536 522164
rect 331956 522112 332008 522164
rect 451924 522112 451976 522164
rect 45100 522044 45152 522096
rect 78496 522044 78548 522096
rect 369124 522044 369176 522096
rect 375564 522044 375616 522096
rect 107844 521976 107896 522028
rect 374092 521976 374144 522028
rect 471060 522044 471112 522096
rect 517520 522248 517572 522300
rect 538680 522248 538732 522300
rect 517520 521976 517572 522028
rect 60924 521908 60976 521960
rect 60832 521840 60884 521892
rect 125968 521908 126020 521960
rect 144828 521908 144880 521960
rect 149244 521908 149296 521960
rect 61108 521840 61160 521892
rect 131120 521840 131172 521892
rect 205180 521840 205232 521892
rect 303620 521840 303672 521892
rect 497464 521840 497516 521892
rect 500960 521840 501012 521892
rect 42616 521772 42668 521824
rect 115940 521772 115992 521824
rect 160560 521772 160612 521824
rect 269028 521772 269080 521824
rect 376668 521772 376720 521824
rect 500592 521772 500644 521824
rect 43812 521704 43864 521756
rect 129096 521704 129148 521756
rect 145472 521704 145524 521756
rect 256700 521704 256752 521756
rect 377956 521704 378008 521756
rect 508596 521704 508648 521756
rect 45192 521636 45244 521688
rect 79416 521636 79468 521688
rect 81624 521636 81676 521688
rect 313280 521636 313332 521688
rect 378784 521636 378836 521688
rect 523224 521636 523276 521688
rect 50988 521568 51040 521620
rect 59360 521568 59412 521620
rect 62856 521568 62908 521620
rect 167092 521568 167144 521620
rect 382280 521568 382332 521620
rect 479524 521568 479576 521620
rect 500132 521568 500184 521620
rect 510252 521568 510304 521620
rect 513472 521568 513524 521620
rect 58440 521500 58492 521552
rect 59452 521500 59504 521552
rect 59728 521500 59780 521552
rect 168380 521500 168432 521552
rect 382372 521500 382424 521552
rect 497556 521500 497608 521552
rect 514760 521500 514812 521552
rect 60556 521432 60608 521484
rect 166264 521432 166316 521484
rect 338948 521432 339000 521484
rect 51540 521364 51592 521416
rect 167000 521364 167052 521416
rect 191104 521364 191156 521416
rect 220728 521364 220780 521416
rect 380992 521364 381044 521416
rect 231768 521296 231820 521348
rect 312636 521296 312688 521348
rect 498752 521296 498804 521348
rect 501236 521296 501288 521348
rect 43628 521228 43680 521280
rect 73344 521228 73396 521280
rect 222108 521228 222160 521280
rect 293316 521228 293368 521280
rect 499028 521228 499080 521280
rect 501788 521228 501840 521280
rect 41144 521160 41196 521212
rect 74448 521160 74500 521212
rect 498936 521160 498988 521212
rect 501328 521160 501380 521212
rect 48780 521092 48832 521144
rect 96620 521092 96672 521144
rect 471244 521092 471296 521144
rect 518256 521092 518308 521144
rect 59636 521024 59688 521076
rect 61844 521024 61896 521076
rect 146484 521024 146536 521076
rect 285680 521024 285732 521076
rect 471428 521024 471480 521076
rect 530308 521024 530360 521076
rect 53748 520956 53800 521008
rect 59268 520956 59320 521008
rect 71872 520956 71924 521008
rect 133144 520956 133196 521008
rect 254768 520956 254820 521008
rect 524880 520956 524932 521008
rect 34428 520888 34480 520940
rect 52460 520888 52512 520940
rect 59820 520888 59872 520940
rect 62764 520888 62816 520940
rect 71964 520888 72016 520940
rect 141148 520888 141200 520940
rect 193956 520888 194008 520940
rect 496728 520888 496780 520940
rect 499212 520888 499264 520940
rect 500776 520888 500828 520940
rect 505928 520888 505980 520940
rect 520372 520888 520424 520940
rect 42248 520820 42300 520872
rect 71320 520820 71372 520872
rect 498844 520820 498896 520872
rect 500684 520820 500736 520872
rect 45376 520752 45428 520804
rect 76472 520752 76524 520804
rect 40868 520684 40920 520736
rect 75368 520684 75420 520736
rect 59268 520616 59320 520668
rect 59728 520616 59780 520668
rect 60004 520616 60056 520668
rect 106832 520616 106884 520668
rect 291844 520616 291896 520668
rect 504272 520752 504324 520804
rect 498108 520684 498160 520736
rect 515036 520684 515088 520736
rect 59452 520548 59504 520600
rect 119896 520548 119948 520600
rect 288348 520548 288400 520600
rect 496176 520548 496228 520600
rect 500408 520548 500460 520600
rect 504364 520548 504416 520600
rect 52368 520480 52420 520532
rect 113916 520480 113968 520532
rect 207204 520480 207256 520532
rect 521844 520480 521896 520532
rect 57980 520412 58032 520464
rect 60188 520412 60240 520464
rect 59728 520344 59780 520396
rect 61660 520412 61712 520464
rect 62120 520412 62172 520464
rect 127992 520412 128044 520464
rect 164700 520412 164752 520464
rect 498016 520412 498068 520464
rect 498108 520412 498160 520464
rect 537208 520412 537260 520464
rect 60556 520344 60608 520396
rect 134064 520344 134116 520396
rect 188988 520344 189040 520396
rect 545304 520344 545356 520396
rect 43536 520276 43588 520328
rect 72332 520276 72384 520328
rect 86684 520276 86736 520328
rect 516416 520276 516468 520328
rect 56140 520208 56192 520260
rect 61108 520208 61160 520260
rect 61200 520208 61252 520260
rect 61844 520208 61896 520260
rect 498200 520208 498252 520260
rect 53288 520140 53340 520192
rect 59636 520140 59688 520192
rect 59820 520140 59872 520192
rect 60464 520140 60516 520192
rect 62028 520140 62080 520192
rect 499304 520140 499356 520192
rect 500684 520208 500736 520260
rect 507952 520208 508004 520260
rect 52736 520072 52788 520124
rect 60188 520072 60240 520124
rect 61752 520072 61804 520124
rect 498016 520072 498068 520124
rect 506020 520140 506072 520192
rect 56508 520004 56560 520056
rect 60648 520004 60700 520056
rect 505928 520072 505980 520124
rect 509240 520072 509292 520124
rect 502248 519868 502300 519920
rect 510620 519868 510672 519920
rect 501236 519800 501288 519852
rect 501328 519800 501380 519852
rect 502248 519732 502300 519784
rect 52368 519664 52420 519716
rect 43720 519596 43772 519648
rect 52552 519596 52604 519648
rect 28908 519528 28960 519580
rect 60004 519528 60056 519580
rect 501328 519664 501380 519716
rect 502156 519664 502208 519716
rect 501880 519596 501932 519648
rect 503720 519596 503772 519648
rect 509516 519596 509568 519648
rect 60924 519528 60976 519580
rect 501328 519528 501380 519580
rect 501696 519528 501748 519580
rect 60832 519460 60884 519512
rect 60648 519052 60700 519104
rect 58716 518984 58768 519036
rect 60924 518984 60976 519036
rect 49516 518916 49568 518968
rect 55864 518916 55916 518968
rect 57704 516128 57756 516180
rect 59360 516128 59412 516180
rect 53748 514836 53800 514888
rect 54576 514836 54628 514888
rect 53472 514768 53524 514820
rect 54484 514768 54536 514820
rect 53656 514700 53708 514752
rect 55864 514700 55916 514752
rect 53288 514020 53340 514072
rect 53656 514020 53708 514072
rect 57980 513272 58032 513324
rect 58532 513272 58584 513324
rect 500316 513272 500368 513324
rect 500960 513272 501012 513324
rect 500500 512592 500552 512644
rect 509332 512592 509384 512644
rect 57888 511912 57940 511964
rect 59452 511912 59504 511964
rect 510528 511912 510580 511964
rect 580172 511912 580224 511964
rect 53288 511232 53340 511284
rect 58624 511232 58676 511284
rect 500408 511232 500460 511284
rect 510528 511232 510580 511284
rect 55036 510620 55088 510672
rect 56600 510620 56652 510672
rect 511448 510008 511500 510060
rect 511632 510008 511684 510060
rect 53748 509872 53800 509924
rect 57980 509872 58032 509924
rect 49516 507832 49568 507884
rect 57152 507832 57204 507884
rect 57796 507832 57848 507884
rect 58716 507832 58768 507884
rect 55864 505112 55916 505164
rect 59360 505112 59412 505164
rect 58532 504364 58584 504416
rect 60188 504364 60240 504416
rect 55128 503616 55180 503668
rect 56600 503616 56652 503668
rect 58440 503616 58492 503668
rect 59820 503616 59872 503668
rect 52828 503072 52880 503124
rect 58624 503072 58676 503124
rect 53656 501576 53708 501628
rect 60096 501576 60148 501628
rect 57704 500896 57756 500948
rect 58072 500896 58124 500948
rect 59820 500148 59872 500200
rect 60188 500148 60240 500200
rect 55128 499536 55180 499588
rect 57244 499536 57296 499588
rect 57612 498992 57664 499044
rect 57612 498788 57664 498840
rect 27528 497428 27580 497480
rect 43352 497428 43404 497480
rect 28908 496748 28960 496800
rect 31852 496748 31904 496800
rect 57704 496272 57756 496324
rect 60280 496272 60332 496324
rect 34428 495456 34480 495508
rect 35072 495456 35124 495508
rect 57152 494708 57204 494760
rect 58716 494708 58768 494760
rect 31852 493960 31904 494012
rect 38108 493960 38160 494012
rect 46480 493280 46532 493332
rect 57980 493280 58032 493332
rect 57152 491580 57204 491632
rect 57520 491580 57572 491632
rect 57796 488588 57848 488640
rect 58808 488588 58860 488640
rect 57704 488520 57756 488572
rect 58072 488520 58124 488572
rect 503628 488452 503680 488504
rect 511172 488452 511224 488504
rect 500040 486072 500092 486124
rect 500500 486072 500552 486124
rect 502340 485392 502392 485444
rect 502432 485188 502484 485240
rect 502984 485052 503036 485104
rect 541440 485052 541492 485104
rect 501604 483624 501656 483676
rect 517704 483624 517756 483676
rect 503536 482944 503588 482996
rect 505836 482944 505888 482996
rect 508596 482400 508648 482452
rect 517704 482400 517756 482452
rect 503444 482332 503496 482384
rect 515588 482332 515640 482384
rect 503168 482264 503220 482316
rect 516876 482264 516928 482316
rect 503076 481720 503128 481772
rect 509884 481720 509936 481772
rect 502984 480836 503036 480888
rect 503260 480836 503312 480888
rect 26884 479476 26936 479528
rect 37924 479476 37976 479528
rect 503260 478864 503312 478916
rect 511264 478864 511316 478916
rect 38108 478116 38160 478168
rect 51816 478116 51868 478168
rect 503536 478116 503588 478168
rect 538680 478116 538732 478168
rect 3424 474716 3476 474768
rect 11704 474716 11756 474768
rect 502892 470500 502944 470552
rect 536288 470500 536340 470552
rect 502892 469140 502944 469192
rect 534908 469140 534960 469192
rect 502800 469072 502852 469124
rect 522396 469072 522448 469124
rect 502708 467780 502760 467832
rect 534724 467780 534776 467832
rect 502800 467712 502852 467764
rect 530676 467712 530728 467764
rect 502892 467644 502944 467696
rect 527916 467644 527968 467696
rect 35072 467100 35124 467152
rect 51080 467100 51132 467152
rect 502708 466352 502760 466404
rect 534632 466352 534684 466404
rect 502616 466284 502668 466336
rect 534540 466284 534592 466336
rect 502800 466216 502852 466268
rect 533252 466216 533304 466268
rect 502892 466148 502944 466200
rect 533344 466148 533396 466200
rect 502892 464992 502944 465044
rect 520924 464992 520976 465044
rect 502616 463632 502668 463684
rect 527824 463632 527876 463684
rect 502708 463564 502760 463616
rect 524972 463564 525024 463616
rect 502800 463496 502852 463548
rect 518256 463496 518308 463548
rect 502892 463428 502944 463480
rect 516784 463428 516836 463480
rect 51080 462272 51132 462324
rect 54760 462272 54812 462324
rect 502524 462272 502576 462324
rect 529296 462272 529348 462324
rect 502892 462204 502944 462256
rect 529112 462204 529164 462256
rect 502616 462136 502668 462188
rect 526536 462136 526588 462188
rect 502892 462068 502944 462120
rect 525064 462068 525116 462120
rect 502800 462000 502852 462052
rect 521016 462000 521068 462052
rect 502800 460844 502852 460896
rect 544476 460844 544528 460896
rect 502892 460776 502944 460828
rect 538588 460776 538640 460828
rect 502616 459484 502668 459536
rect 531688 459484 531740 459536
rect 502892 459416 502944 459468
rect 530492 459416 530544 459468
rect 502800 459348 502852 459400
rect 529020 459348 529072 459400
rect 502708 459280 502760 459332
rect 522212 459280 522264 459332
rect 502800 458124 502852 458176
rect 534448 458124 534500 458176
rect 535736 458124 535788 458176
rect 580172 458124 580224 458176
rect 502616 458056 502668 458108
rect 537300 458056 537352 458108
rect 502708 457988 502760 458040
rect 526352 457988 526404 458040
rect 502892 457920 502944 457972
rect 518072 457920 518124 457972
rect 501696 457444 501748 457496
rect 535736 457444 535788 457496
rect 502616 456696 502668 456748
rect 536012 456696 536064 456748
rect 502892 456628 502944 456680
rect 533160 456628 533212 456680
rect 502800 456560 502852 456612
rect 530400 456560 530452 456612
rect 502892 456492 502944 456544
rect 513932 456492 513984 456544
rect 502708 455336 502760 455388
rect 531596 455336 531648 455388
rect 502524 455268 502576 455320
rect 523316 455268 523368 455320
rect 502616 455200 502668 455252
rect 522120 455200 522172 455252
rect 502800 455132 502852 455184
rect 512184 455132 512236 455184
rect 502892 455064 502944 455116
rect 509792 455064 509844 455116
rect 502892 453908 502944 453960
rect 519636 453908 519688 453960
rect 502708 453840 502760 453892
rect 514852 453840 514904 453892
rect 502800 453772 502852 453824
rect 541624 453772 541676 453824
rect 502708 452548 502760 452600
rect 515312 452548 515364 452600
rect 502616 452480 502668 452532
rect 515128 452480 515180 452532
rect 502892 452412 502944 452464
rect 514944 452412 514996 452464
rect 502800 452344 502852 452396
rect 513840 452344 513892 452396
rect 502616 451188 502668 451240
rect 526260 451188 526312 451240
rect 502708 451120 502760 451172
rect 520740 451120 520792 451172
rect 503628 451052 503680 451104
rect 513748 451052 513800 451104
rect 502892 450984 502944 451036
rect 512828 450984 512880 451036
rect 503628 450916 503680 450968
rect 507216 450916 507268 450968
rect 503628 449828 503680 449880
rect 537116 449828 537168 449880
rect 502708 449760 502760 449812
rect 537024 449760 537076 449812
rect 502800 449692 502852 449744
rect 527640 449692 527692 449744
rect 502892 449624 502944 449676
rect 524696 449624 524748 449676
rect 503628 449556 503680 449608
rect 517980 449556 518032 449608
rect 502708 448468 502760 448520
rect 540336 448468 540388 448520
rect 502616 448400 502668 448452
rect 538496 448400 538548 448452
rect 503628 448332 503680 448384
rect 516600 448332 516652 448384
rect 502892 448264 502944 448316
rect 513564 448264 513616 448316
rect 503628 445680 503680 445732
rect 538404 445680 538456 445732
rect 499856 444456 499908 444508
rect 500132 444456 500184 444508
rect 503628 442892 503680 442944
rect 545764 442892 545816 442944
rect 500224 441940 500276 441992
rect 500868 441940 500920 441992
rect 503628 441124 503680 441176
rect 508504 441124 508556 441176
rect 501880 440308 501932 440360
rect 503536 440308 503588 440360
rect 501788 440240 501840 440292
rect 502432 440240 502484 440292
rect 503628 440172 503680 440224
rect 512920 440172 512972 440224
rect 503628 440036 503680 440088
rect 510804 440036 510856 440088
rect 503536 438812 503588 438864
rect 526168 438812 526220 438864
rect 503628 438744 503680 438796
rect 524880 438744 524932 438796
rect 503628 437384 503680 437436
rect 515220 437384 515272 437436
rect 503628 437044 503680 437096
rect 511080 437044 511132 437096
rect 502892 436772 502944 436824
rect 503444 436772 503496 436824
rect 503628 436024 503680 436076
rect 541532 436024 541584 436076
rect 503444 435956 503496 436008
rect 506940 435956 506992 436008
rect 502800 434664 502852 434716
rect 506572 434664 506624 434716
rect 503536 434596 503588 434648
rect 530216 434596 530268 434648
rect 503628 434528 503680 434580
rect 526076 434528 526128 434580
rect 503444 434460 503496 434512
rect 530032 434460 530084 434512
rect 502616 433236 502668 433288
rect 505560 433236 505612 433288
rect 503444 433168 503496 433220
rect 506848 433168 506900 433220
rect 503536 433100 503588 433152
rect 506756 433100 506808 433152
rect 503628 433032 503680 433084
rect 507400 433032 507452 433084
rect 503444 432964 503496 433016
rect 506664 432964 506716 433016
rect 503444 431876 503496 431928
rect 545672 431876 545724 431928
rect 503628 431740 503680 431792
rect 521936 431740 521988 431792
rect 503536 431672 503588 431724
rect 523500 431672 523552 431724
rect 502524 431400 502576 431452
rect 505376 431400 505428 431452
rect 502708 431264 502760 431316
rect 505744 431264 505796 431316
rect 502616 430516 502668 430568
rect 505652 430516 505704 430568
rect 503628 430448 503680 430500
rect 528928 430448 528980 430500
rect 503444 430380 503496 430432
rect 525984 430380 526036 430432
rect 503536 430312 503588 430364
rect 532976 430312 533028 430364
rect 57704 429156 57756 429208
rect 58532 429156 58584 429208
rect 502524 429088 502576 429140
rect 505468 429088 505520 429140
rect 503628 429020 503680 429072
rect 529940 429020 529992 429072
rect 503628 428816 503680 428868
rect 530124 428816 530176 428868
rect 503628 428612 503680 428664
rect 508044 428612 508096 428664
rect 503628 428340 503680 428392
rect 508228 428340 508280 428392
rect 503444 427728 503496 427780
rect 528836 427728 528888 427780
rect 503536 427660 503588 427712
rect 527364 427660 527416 427712
rect 503628 427592 503680 427644
rect 519360 427592 519412 427644
rect 502800 427524 502852 427576
rect 508136 427524 508188 427576
rect 502708 427456 502760 427508
rect 508320 427456 508372 427508
rect 503444 426368 503496 426420
rect 530308 426368 530360 426420
rect 503628 426300 503680 426352
rect 527456 426300 527508 426352
rect 503536 426232 503588 426284
rect 515036 426232 515088 426284
rect 503628 425008 503680 425060
rect 537208 425008 537260 425060
rect 503444 424940 503496 424992
rect 535828 424940 535880 424992
rect 503536 424872 503588 424924
rect 527548 424872 527600 424924
rect 503628 424804 503680 424856
rect 513656 424804 513708 424856
rect 503628 423580 503680 423632
rect 524604 423580 524656 423632
rect 3424 422288 3476 422340
rect 14464 422288 14516 422340
rect 43352 420180 43404 420232
rect 46204 420180 46256 420232
rect 54760 400868 54812 400920
rect 57520 400868 57572 400920
rect 37924 392572 37976 392624
rect 51080 392572 51132 392624
rect 60372 391620 60424 391672
rect 62028 391620 62080 391672
rect 498200 390600 498252 390652
rect 500316 390600 500368 390652
rect 325516 390260 325568 390312
rect 503352 390260 503404 390312
rect 14464 390192 14516 390244
rect 96528 390192 96580 390244
rect 306288 390192 306340 390244
rect 501696 390192 501748 390244
rect 58532 390124 58584 390176
rect 144184 390124 144236 390176
rect 343088 390124 343140 390176
rect 544200 390124 544252 390176
rect 57520 390056 57572 390108
rect 220728 390056 220780 390108
rect 346216 390056 346268 390108
rect 545488 390056 545540 390108
rect 62028 389988 62080 390040
rect 273904 389988 273956 390040
rect 308128 389988 308180 390040
rect 500408 389988 500460 390040
rect 51816 389920 51868 389972
rect 274732 389920 274784 389972
rect 485780 389920 485832 389972
rect 501880 389920 501932 389972
rect 46204 389852 46256 389904
rect 294604 389852 294656 389904
rect 398104 389852 398156 389904
rect 498200 389852 498252 389904
rect 51080 389784 51132 389836
rect 326344 389784 326396 389836
rect 360476 389784 360528 389836
rect 525892 389784 525944 389836
rect 309784 389104 309836 389156
rect 537760 389104 537812 389156
rect 311164 389036 311216 389088
rect 537576 389036 537628 389088
rect 346308 388968 346360 389020
rect 543924 388968 543976 389020
rect 349804 388900 349856 388952
rect 505836 388900 505888 388952
rect 319720 388832 319772 388884
rect 398104 388832 398156 388884
rect 400312 388832 400364 388884
rect 545580 388832 545632 388884
rect 398840 388492 398892 388544
rect 499948 388492 500000 388544
rect 11704 388424 11756 388476
rect 95148 388424 95200 388476
rect 359648 388424 359700 388476
rect 509516 388424 509568 388476
rect 96528 387744 96580 387796
rect 339316 387744 339368 387796
rect 343640 387744 343692 387796
rect 344560 387744 344612 387796
rect 546592 387744 546644 387796
rect 95148 387676 95200 387728
rect 337568 387676 337620 387728
rect 544108 387676 544160 387728
rect 314844 387608 314896 387660
rect 315304 387608 315356 387660
rect 539232 387608 539284 387660
rect 37096 387540 37148 387592
rect 89720 387540 89772 387592
rect 292120 387540 292172 387592
rect 359648 387540 359700 387592
rect 32772 387472 32824 387524
rect 91192 387472 91244 387524
rect 221832 387472 221884 387524
rect 343640 387472 343692 387524
rect 348424 387472 348476 387524
rect 547972 387472 548024 387524
rect 45468 387404 45520 387456
rect 106188 387404 106240 387456
rect 327080 387404 327132 387456
rect 85580 387336 85632 387388
rect 86868 387336 86920 387388
rect 328828 387336 328880 387388
rect 86960 387268 87012 387320
rect 88248 387268 88300 387320
rect 330576 387268 330628 387320
rect 31576 387200 31628 387252
rect 89628 387200 89680 387252
rect 332324 387200 332376 387252
rect 341524 387200 341576 387252
rect 360200 387200 360252 387252
rect 27160 387132 27212 387184
rect 85580 387132 85632 387184
rect 89720 387132 89772 387184
rect 91008 387132 91060 387184
rect 334072 387132 334124 387184
rect 359740 387132 359792 387184
rect 403992 387132 404044 387184
rect 26148 387064 26200 387116
rect 86960 387064 87012 387116
rect 91192 387064 91244 387116
rect 92388 387064 92440 387116
rect 335820 387064 335872 387116
rect 339316 387064 339368 387116
rect 360108 387064 360160 387116
rect 360384 387064 360436 387116
rect 419724 387064 419776 387116
rect 293868 386996 293920 387048
rect 355968 386996 356020 387048
rect 360476 386996 360528 387048
rect 360108 386520 360160 386572
rect 394608 386520 394660 386572
rect 360200 386452 360252 386504
rect 395988 386452 396040 386504
rect 302884 386384 302936 386436
rect 498200 386384 498252 386436
rect 220728 386316 220780 386368
rect 227720 386316 227772 386368
rect 394608 386316 394660 386368
rect 544016 386316 544068 386368
rect 395988 386248 396040 386300
rect 545396 386248 545448 386300
rect 466368 385636 466420 385688
rect 485780 385636 485832 385688
rect 282092 384956 282144 385008
rect 491392 384956 491444 385008
rect 355968 384888 356020 384940
rect 542728 384888 542780 384940
rect 357348 384820 357400 384872
rect 542820 384820 542872 384872
rect 274732 384344 274784 384396
rect 287704 384344 287756 384396
rect 498200 384344 498252 384396
rect 529940 384344 529992 384396
rect 239956 384276 240008 384328
rect 580356 384276 580408 384328
rect 234620 383664 234672 383716
rect 313924 383664 313976 383716
rect 498844 383664 498896 383716
rect 501788 383664 501840 383716
rect 294604 382916 294656 382968
rect 308496 382916 308548 382968
rect 445668 382916 445720 382968
rect 466368 382916 466420 382968
rect 273904 382236 273956 382288
rect 276664 382236 276716 382288
rect 529940 382236 529992 382288
rect 531228 382236 531280 382288
rect 532792 382236 532844 382288
rect 240048 382168 240100 382220
rect 535552 382168 535604 382220
rect 266360 382100 266412 382152
rect 527272 382100 527324 382152
rect 227720 380128 227772 380180
rect 236000 380128 236052 380180
rect 282552 378836 282604 378888
rect 541256 378836 541308 378888
rect 144184 378768 144236 378820
rect 146944 378768 146996 378820
rect 282276 378768 282328 378820
rect 541348 378768 541400 378820
rect 239312 378156 239364 378208
rect 580172 378156 580224 378208
rect 436744 377408 436796 377460
rect 445668 377408 445720 377460
rect 234620 376660 234672 376712
rect 530768 376660 530820 376712
rect 485964 376592 486016 376644
rect 549260 376592 549312 376644
rect 282460 376048 282512 376100
rect 539968 376048 540020 376100
rect 231216 375980 231268 376032
rect 537668 375980 537720 376032
rect 236000 375368 236052 375420
rect 238852 375368 238904 375420
rect 287704 375300 287756 375352
rect 294604 375300 294656 375352
rect 276020 373940 276072 373992
rect 511448 373940 511500 373992
rect 238852 373260 238904 373312
rect 264980 373260 265032 373312
rect 97908 371832 97960 371884
rect 341524 371832 341576 371884
rect 3424 371220 3476 371272
rect 97908 371220 97960 371272
rect 264980 369112 265032 369164
rect 276020 369112 276072 369164
rect 359372 369112 359424 369164
rect 435456 369112 435508 369164
rect 495440 368772 495492 368824
rect 498844 368772 498896 368824
rect 358360 367752 358412 367804
rect 479156 367752 479208 367804
rect 276020 366664 276072 366716
rect 293592 366664 293644 366716
rect 294604 366664 294656 366716
rect 306012 366664 306064 366716
rect 57428 366596 57480 366648
rect 341524 366596 341576 366648
rect 29736 366528 29788 366580
rect 333244 366528 333296 366580
rect 356704 366528 356756 366580
rect 452936 366528 452988 366580
rect 29828 366460 29880 366512
rect 358084 366460 358136 366512
rect 487804 366460 487856 366512
rect 495440 366460 495492 366512
rect 43536 366392 43588 366444
rect 502340 366392 502392 366444
rect 42248 366324 42300 366376
rect 501144 366324 501196 366376
rect 420920 365032 420972 365084
rect 436744 365032 436796 365084
rect 43628 364964 43680 365016
rect 502432 364964 502484 365016
rect 146944 364352 146996 364404
rect 153844 364352 153896 364404
rect 60280 364216 60332 364268
rect 341708 364216 341760 364268
rect 46664 364148 46716 364200
rect 333428 364148 333480 364200
rect 42432 364080 42484 364132
rect 336004 364080 336056 364132
rect 40960 364012 41012 364064
rect 338764 364012 338816 364064
rect 47400 363944 47452 363996
rect 347044 363944 347096 363996
rect 29920 363876 29972 363928
rect 333336 363876 333388 363928
rect 39948 363808 40000 363860
rect 347136 363808 347188 363860
rect 43720 363740 43772 363792
rect 359464 363740 359516 363792
rect 477500 363740 477552 363792
rect 487804 363740 487856 363792
rect 42340 363672 42392 363724
rect 499672 363672 499724 363724
rect 45100 363604 45152 363656
rect 505100 363604 505152 363656
rect 45192 362176 45244 362228
rect 503904 362176 503956 362228
rect 60464 361360 60516 361412
rect 336372 361360 336424 361412
rect 59268 361292 59320 361344
rect 336188 361292 336240 361344
rect 58624 361224 58676 361276
rect 336280 361224 336332 361276
rect 57888 361156 57940 361208
rect 338856 361156 338908 361208
rect 41052 361088 41104 361140
rect 336096 361088 336148 361140
rect 25780 361020 25832 361072
rect 347228 361020 347280 361072
rect 25964 360952 26016 361004
rect 355324 360952 355376 361004
rect 25596 360884 25648 360936
rect 359556 360884 359608 360936
rect 408500 360884 408552 360936
rect 420920 360884 420972 360936
rect 45284 360816 45336 360868
rect 503812 360816 503864 360868
rect 253204 359524 253256 359576
rect 430212 359524 430264 359576
rect 40868 359456 40920 359508
rect 502524 359456 502576 359508
rect 252468 358844 252520 358896
rect 289084 358844 289136 358896
rect 252376 358776 252428 358828
rect 294604 358776 294656 358828
rect 271788 358640 271840 358692
rect 282920 358640 282972 358692
rect 272432 358572 272484 358624
rect 472164 358572 472216 358624
rect 273352 358504 273404 358556
rect 473912 358504 473964 358556
rect 274272 358436 274324 358488
rect 475660 358436 475712 358488
rect 275192 358368 275244 358420
rect 477408 358368 477460 358420
rect 60188 358300 60240 358352
rect 302240 358300 302292 358352
rect 57336 358232 57388 358284
rect 338948 358232 339000 358284
rect 56232 358164 56284 358216
rect 347320 358164 347372 358216
rect 54576 358096 54628 358148
rect 349896 358096 349948 358148
rect 53288 358028 53340 358080
rect 349804 358028 349856 358080
rect 402244 358028 402296 358080
rect 408500 358028 408552 358080
rect 474648 357620 474700 357672
rect 477500 357620 477552 357672
rect 271788 357416 271840 357468
rect 303620 357416 303672 357468
rect 260472 356804 260524 356856
rect 449440 356804 449492 356856
rect 261392 356736 261444 356788
rect 451188 356736 451240 356788
rect 45376 356668 45428 356720
rect 502708 356668 502760 356720
rect 238392 355920 238444 355972
rect 284300 355920 284352 355972
rect 276020 355852 276072 355904
rect 532700 355852 532752 355904
rect 269028 355784 269080 355836
rect 534080 355784 534132 355836
rect 60096 355716 60148 355768
rect 341892 355716 341944 355768
rect 58716 355648 58768 355700
rect 341800 355648 341852 355700
rect 57244 355580 57296 355632
rect 344376 355580 344428 355632
rect 238208 355512 238260 355564
rect 529940 355512 529992 355564
rect 53104 355444 53156 355496
rect 344284 355444 344336 355496
rect 58808 355376 58860 355428
rect 355416 355376 355468 355428
rect 452660 355376 452712 355428
rect 474648 355376 474700 355428
rect 237748 355308 237800 355360
rect 536104 355308 536156 355360
rect 240048 354628 240100 354680
rect 580448 354628 580500 354680
rect 237840 353948 237892 354000
rect 452660 353948 452712 354000
rect 239404 353404 239456 353456
rect 296812 353404 296864 353456
rect 237104 353336 237156 353388
rect 295340 353336 295392 353388
rect 237012 353268 237064 353320
rect 296720 353268 296772 353320
rect 240048 353200 240100 353252
rect 402244 353200 402296 353252
rect 531228 353200 531280 353252
rect 580172 353200 580224 353252
rect 282092 353132 282144 353184
rect 539600 353132 539652 353184
rect 60556 353064 60608 353116
rect 350080 353064 350132 353116
rect 52736 352996 52788 353048
rect 347504 352996 347556 353048
rect 52368 352928 52420 352980
rect 347412 352928 347464 352980
rect 56140 352860 56192 352912
rect 352656 352860 352708 352912
rect 54484 352792 54536 352844
rect 352748 352792 352800 352844
rect 46480 352724 46532 352776
rect 349988 352724 350040 352776
rect 46756 352656 46808 352708
rect 352564 352656 352616 352708
rect 28632 352588 28684 352640
rect 355508 352588 355560 352640
rect 27344 352520 27396 352572
rect 355600 352520 355652 352572
rect 235356 351908 235408 351960
rect 288440 351908 288492 351960
rect 234988 351772 235040 351824
rect 235356 351772 235408 351824
rect 359924 351432 359976 351484
rect 503260 351432 503312 351484
rect 282000 351364 282052 351416
rect 541164 351364 541216 351416
rect 239588 351296 239640 351348
rect 510068 351296 510120 351348
rect 239864 351228 239916 351280
rect 580264 351228 580316 351280
rect 43260 351160 43312 351212
rect 503720 351160 503772 351212
rect 229928 351092 229980 351144
rect 280252 351092 280304 351144
rect 230296 351024 230348 351076
rect 283012 351024 283064 351076
rect 224684 350956 224736 351008
rect 280344 350956 280396 351008
rect 221464 350888 221516 350940
rect 277952 350888 278004 350940
rect 224224 350820 224276 350872
rect 290556 350820 290608 350872
rect 217416 350752 217468 350804
rect 288716 350752 288768 350804
rect 217324 350684 217376 350736
rect 291568 350684 291620 350736
rect 237932 350616 237984 350668
rect 318064 350616 318116 350668
rect 222108 350548 222160 350600
rect 311256 350548 311308 350600
rect 232504 350480 232556 350532
rect 240048 350480 240100 350532
rect 226340 350344 226392 350396
rect 298100 350344 298152 350396
rect 282736 350276 282788 350328
rect 539784 350276 539836 350328
rect 50804 350208 50856 350260
rect 336464 350208 336516 350260
rect 55864 350140 55916 350192
rect 344468 350140 344520 350192
rect 42616 350072 42668 350124
rect 339040 350072 339092 350124
rect 43812 350004 43864 350056
rect 352840 350004 352892 350056
rect 48780 349936 48832 349988
rect 359648 349936 359700 349988
rect 43904 349868 43956 349920
rect 501236 349868 501288 349920
rect 41144 349800 41196 349852
rect 502616 349800 502668 349852
rect 153844 349732 153896 349784
rect 158720 349732 158772 349784
rect 254584 349324 254636 349376
rect 292580 349324 292632 349376
rect 234988 349256 235040 349308
rect 580264 349256 580316 349308
rect 220176 349188 220228 349240
rect 283380 349188 283432 349240
rect 221648 349120 221700 349172
rect 302332 349120 302384 349172
rect 259368 348576 259420 348628
rect 302516 348576 302568 348628
rect 233976 348508 234028 348560
rect 282920 348508 282972 348560
rect 226524 348440 226576 348492
rect 278044 348440 278096 348492
rect 212264 348372 212316 348424
rect 312544 348372 312596 348424
rect 249708 348304 249760 348356
rect 301044 348304 301096 348356
rect 232688 348236 232740 348288
rect 284300 348236 284352 348288
rect 226432 348168 226484 348220
rect 290648 348168 290700 348220
rect 226340 348100 226392 348152
rect 299572 348100 299624 348152
rect 222108 348032 222160 348084
rect 296076 348032 296128 348084
rect 212448 347964 212500 348016
rect 287796 347964 287848 348016
rect 220728 347896 220780 347948
rect 298836 347896 298888 347948
rect 211988 347828 212040 347880
rect 292856 347828 292908 347880
rect 224224 347760 224276 347812
rect 322296 347760 322348 347812
rect 60648 347216 60700 347268
rect 350264 347216 350316 347268
rect 50620 347148 50672 347200
rect 344560 347148 344612 347200
rect 47952 347080 48004 347132
rect 350172 347080 350224 347132
rect 31484 347012 31536 347064
rect 358176 347012 358228 347064
rect 266360 346944 266412 346996
rect 285772 346944 285824 346996
rect 273260 346876 273312 346928
rect 298284 346876 298336 346928
rect 243544 346808 243596 346860
rect 283196 346808 283248 346860
rect 226064 346740 226116 346792
rect 280528 346740 280580 346792
rect 224224 346672 224276 346724
rect 291200 346672 291252 346724
rect 220728 346604 220780 346656
rect 289268 346604 289320 346656
rect 223304 346536 223356 346588
rect 303068 346536 303120 346588
rect 225052 346468 225104 346520
rect 314108 346468 314160 346520
rect 224960 346400 225012 346452
rect 325056 346400 325108 346452
rect 260748 346332 260800 346384
rect 360384 346332 360436 346384
rect 503628 346332 503680 346384
rect 523408 346332 523460 346384
rect 253112 346264 253164 346316
rect 273260 346264 273312 346316
rect 229744 345856 229796 345908
rect 280160 345856 280212 345908
rect 227720 345788 227772 345840
rect 278964 345788 279016 345840
rect 225880 345720 225932 345772
rect 284300 345720 284352 345772
rect 216680 345652 216732 345704
rect 304356 345652 304408 345704
rect 274640 345584 274692 345636
rect 295524 345584 295576 345636
rect 244280 345516 244332 345568
rect 298192 345516 298244 345568
rect 223212 345448 223264 345500
rect 289360 345448 289412 345500
rect 228364 345380 228416 345432
rect 299480 345380 299532 345432
rect 158720 345312 158772 345364
rect 161572 345312 161624 345364
rect 226340 345312 226392 345364
rect 307300 345312 307352 345364
rect 223304 345244 223356 345296
rect 305828 345244 305880 345296
rect 209136 345176 209188 345228
rect 296904 345176 296956 345228
rect 223120 345108 223172 345160
rect 327724 345108 327776 345160
rect 220728 345040 220780 345092
rect 334624 345040 334676 345092
rect 243544 344972 243596 345024
rect 360292 344972 360344 345024
rect 228456 344360 228508 344412
rect 254584 344360 254636 344412
rect 271788 344360 271840 344412
rect 287244 344360 287296 344412
rect 251088 344292 251140 344344
rect 279332 344292 279384 344344
rect 293592 344292 293644 344344
rect 304540 344292 304592 344344
rect 255320 344224 255372 344276
rect 292764 344224 292816 344276
rect 236000 344156 236052 344208
rect 285036 344156 285088 344208
rect 218060 344088 218112 344140
rect 293316 344088 293368 344140
rect 231124 344020 231176 344072
rect 316684 344020 316736 344072
rect 216680 343952 216732 344004
rect 307116 343952 307168 344004
rect 228272 343884 228324 343936
rect 319444 343884 319496 343936
rect 224224 343816 224276 343868
rect 319536 343816 319588 343868
rect 214564 343748 214616 343800
rect 314016 343748 314068 343800
rect 125508 343680 125560 343732
rect 322204 343680 322256 343732
rect 61936 343612 61988 343664
rect 302884 343612 302936 343664
rect 231124 343204 231176 343256
rect 280712 343204 280764 343256
rect 276112 343136 276164 343188
rect 358360 343136 358412 343188
rect 262312 343068 262364 343120
rect 356704 343068 356756 343120
rect 250352 343000 250404 343052
rect 253204 343000 253256 343052
rect 253480 343000 253532 343052
rect 359372 343000 359424 343052
rect 161572 342932 161624 342984
rect 176660 342932 176712 342984
rect 239220 342932 239272 342984
rect 358544 342932 358596 342984
rect 60004 342864 60056 342916
rect 350356 342864 350408 342916
rect 221740 342796 221792 342848
rect 276020 342796 276072 342848
rect 224224 342728 224276 342780
rect 282920 342728 282972 342780
rect 209228 342660 209280 342712
rect 279424 342660 279476 342712
rect 214564 342592 214616 342644
rect 286600 342592 286652 342644
rect 214472 342524 214524 342576
rect 287980 342524 288032 342576
rect 220360 342456 220412 342508
rect 305644 342456 305696 342508
rect 306104 342456 306156 342508
rect 244280 342388 244332 342440
rect 339224 342388 339276 342440
rect 214656 342320 214708 342372
rect 311348 342320 311400 342372
rect 214380 342252 214432 342304
rect 320824 342252 320876 342304
rect 240048 342184 240100 342236
rect 356796 342184 356848 342236
rect 270408 341708 270460 341760
rect 295708 341708 295760 341760
rect 256700 341640 256752 341692
rect 285864 341640 285916 341692
rect 231124 341572 231176 341624
rect 280620 341572 280672 341624
rect 216680 341504 216732 341556
rect 285680 341504 285732 341556
rect 224960 341436 225012 341488
rect 300400 341436 300452 341488
rect 228548 341368 228600 341420
rect 323584 341368 323636 341420
rect 223304 341300 223356 341352
rect 321008 341300 321060 341352
rect 236000 341232 236052 341284
rect 342904 341232 342956 341284
rect 220728 341164 220780 341216
rect 336556 341164 336608 341216
rect 68928 341096 68980 341148
rect 311164 341096 311216 341148
rect 66076 341028 66128 341080
rect 307852 341028 307904 341080
rect 308404 341028 308456 341080
rect 66168 340960 66220 341012
rect 309784 340960 309836 341012
rect 71596 340892 71648 340944
rect 315304 340892 315356 340944
rect 216680 340824 216732 340876
rect 348424 340824 348476 340876
rect 503628 340824 503680 340876
rect 520648 340824 520700 340876
rect 216864 340756 216916 340808
rect 342812 340756 342864 340808
rect 278044 340416 278096 340468
rect 303712 340416 303764 340468
rect 276020 340348 276072 340400
rect 302424 340348 302476 340400
rect 236920 340280 236972 340332
rect 355048 340280 355100 340332
rect 238392 340212 238444 340264
rect 359740 340212 359792 340264
rect 103428 340144 103480 340196
rect 346308 340144 346360 340196
rect 279056 340076 279108 340128
rect 281356 340076 281408 340128
rect 242440 340008 242492 340060
rect 275744 340008 275796 340060
rect 280068 340008 280120 340060
rect 281172 340008 281224 340060
rect 241428 339940 241480 339992
rect 250996 339940 251048 339992
rect 279792 339940 279844 339992
rect 281264 339940 281316 339992
rect 250904 339872 250956 339924
rect 300952 339872 301004 339924
rect 229928 339804 229980 339856
rect 289544 339804 289596 339856
rect 221924 339736 221976 339788
rect 283564 339736 283616 339788
rect 222016 339668 222068 339720
rect 284300 339668 284352 339720
rect 216772 339600 216824 339652
rect 294788 339600 294840 339652
rect 220728 339532 220780 339584
rect 309968 339532 310020 339584
rect 274640 339464 274692 339516
rect 298100 339464 298152 339516
rect 176660 339396 176712 339448
rect 181444 339396 181496 339448
rect 279332 339396 279384 339448
rect 279424 339396 279476 339448
rect 279516 339396 279568 339448
rect 279608 339396 279660 339448
rect 279976 339396 280028 339448
rect 283748 339396 283800 339448
rect 358360 339396 358412 339448
rect 284852 339192 284904 339244
rect 280160 338920 280212 338972
rect 294328 338920 294380 338972
rect 298376 338852 298428 338904
rect 301228 338784 301280 338836
rect 280068 338716 280120 338768
rect 324964 338716 325016 338768
rect 239128 338580 239180 338632
rect 239772 338580 239824 338632
rect 228640 338444 228692 338496
rect 231124 338444 231176 338496
rect 217508 338308 217560 338360
rect 292948 338308 293000 338360
rect 280160 338240 280212 338292
rect 289912 338240 289964 338292
rect 280068 338172 280120 338224
rect 291476 338172 291528 338224
rect 280160 336132 280212 336184
rect 281080 336132 281132 336184
rect 503628 333888 503680 333940
rect 516508 333888 516560 333940
rect 326344 330488 326396 330540
rect 329196 330488 329248 330540
rect 503628 328380 503680 328432
rect 517796 328380 517848 328432
rect 304540 322872 304592 322924
rect 308680 322872 308732 322924
rect 503628 322872 503680 322924
rect 520556 322872 520608 322924
rect 90364 320832 90416 320884
rect 125600 320832 125652 320884
rect 3424 319404 3476 319456
rect 98644 319404 98696 319456
rect 88984 317432 89036 317484
rect 124864 317364 124916 317416
rect 228272 317364 228324 317416
rect 281816 307708 281868 307760
rect 284300 307708 284352 307760
rect 329196 307708 329248 307760
rect 331956 307708 332008 307760
rect 503628 304920 503680 304972
rect 519268 304920 519320 304972
rect 106188 303628 106240 303680
rect 129924 303628 129976 303680
rect 181444 303628 181496 303680
rect 186964 303628 187016 303680
rect 306012 303560 306064 303612
rect 309048 303560 309100 303612
rect 79416 303084 79468 303136
rect 90364 303084 90416 303136
rect 83924 303016 83976 303068
rect 106188 303016 106240 303068
rect 77852 302948 77904 303000
rect 88984 302948 89036 303000
rect 126796 302948 126848 303000
rect 221832 302948 221884 303000
rect 63500 302880 63552 302932
rect 64328 302880 64380 302932
rect 220360 302880 220412 302932
rect 66168 302812 66220 302864
rect 67180 302812 67232 302864
rect 71596 302812 71648 302864
rect 72148 302812 72200 302864
rect 94320 302744 94372 302796
rect 95148 302744 95200 302796
rect 132500 302608 132552 302660
rect 102600 302540 102652 302592
rect 103428 302540 103480 302592
rect 111800 302540 111852 302592
rect 104808 302472 104860 302524
rect 124220 302472 124272 302524
rect 89628 302404 89680 302456
rect 124312 302404 124364 302456
rect 46848 302336 46900 302388
rect 57152 302336 57204 302388
rect 92388 302336 92440 302388
rect 129832 302336 129884 302388
rect 45376 302268 45428 302320
rect 55588 302268 55640 302320
rect 82728 302268 82780 302320
rect 95148 302268 95200 302320
rect 88248 302200 88300 302252
rect 131120 302200 131172 302252
rect 95148 301452 95200 301504
rect 128452 301452 128504 301504
rect 100484 301044 100536 301096
rect 125784 301044 125836 301096
rect 126796 301044 126848 301096
rect 98644 300976 98696 301028
rect 131304 300976 131356 301028
rect 46756 300908 46808 300960
rect 53932 300908 53984 300960
rect 91008 300908 91060 300960
rect 128360 300908 128412 300960
rect 47860 300840 47912 300892
rect 58900 300840 58952 300892
rect 86132 300840 86184 300892
rect 86868 300840 86920 300892
rect 129740 300840 129792 300892
rect 128452 300772 128504 300824
rect 129004 300772 129056 300824
rect 228640 300772 228692 300824
rect 47584 299548 47636 299600
rect 50252 299480 50304 299532
rect 52460 299480 52512 299532
rect 100300 299480 100352 299532
rect 357348 299480 357400 299532
rect 531964 299412 532016 299464
rect 580172 299412 580224 299464
rect 357348 299276 357400 299328
rect 281908 298120 281960 298172
rect 292672 298120 292724 298172
rect 309048 298052 309100 298104
rect 315580 298052 315632 298104
rect 503628 298052 503680 298104
rect 516416 298052 516468 298104
rect 331956 295332 332008 295384
rect 337384 295332 337436 295384
rect 281816 292544 281868 292596
rect 284300 292544 284352 292596
rect 503628 292476 503680 292528
rect 519176 292476 519228 292528
rect 281908 291184 281960 291236
rect 284484 291184 284536 291236
rect 281908 289824 281960 289876
rect 284576 289824 284628 289876
rect 281908 288396 281960 288448
rect 294052 288396 294104 288448
rect 339224 288328 339276 288380
rect 357532 288328 357584 288380
rect 503628 286968 503680 287020
rect 520464 286968 520516 287020
rect 337384 285676 337436 285728
rect 342260 285676 342312 285728
rect 342904 282820 342956 282872
rect 357532 282820 357584 282872
rect 342260 279420 342312 279472
rect 351184 279420 351236 279472
rect 285036 277312 285088 277364
rect 357532 277312 357584 277364
rect 315580 275272 315632 275324
rect 318248 275272 318300 275324
rect 503628 274592 503680 274644
rect 516324 274592 516376 274644
rect 289544 273164 289596 273216
rect 357532 273164 357584 273216
rect 307300 271804 307352 271856
rect 357532 271804 357584 271856
rect 290648 270444 290700 270496
rect 357532 270444 357584 270496
rect 282092 269016 282144 269068
rect 284852 269016 284904 269068
rect 282828 268948 282880 269000
rect 287244 268948 287296 269000
rect 3424 267656 3476 267708
rect 47584 267656 47636 267708
rect 282828 266296 282880 266348
rect 295708 266296 295760 266348
rect 282828 264868 282880 264920
rect 294328 264868 294380 264920
rect 282736 263508 282788 263560
rect 292948 263508 293000 263560
rect 282828 263440 282880 263492
rect 291568 263440 291620 263492
rect 282828 262148 282880 262200
rect 288716 262148 288768 262200
rect 325056 262148 325108 262200
rect 357532 262148 357584 262200
rect 282828 260788 282880 260840
rect 301044 260788 301096 260840
rect 318248 260788 318300 260840
rect 323768 260788 323820 260840
rect 186964 259360 187016 259412
rect 189724 259360 189776 259412
rect 282828 259360 282880 259412
rect 302516 259360 302568 259412
rect 282644 259292 282696 259344
rect 299572 259292 299624 259344
rect 282736 259224 282788 259276
rect 292856 259224 292908 259276
rect 282736 258000 282788 258052
rect 299664 258000 299716 258052
rect 282828 257932 282880 257984
rect 298284 257932 298336 257984
rect 282644 256640 282696 256692
rect 299480 256640 299532 256692
rect 300400 256640 300452 256692
rect 357532 256640 357584 256692
rect 282828 256572 282880 256624
rect 298192 256572 298244 256624
rect 282736 256504 282788 256556
rect 296904 256504 296956 256556
rect 286600 255212 286652 255264
rect 357532 255212 357584 255264
rect 282828 255144 282880 255196
rect 301228 255144 301280 255196
rect 282644 253852 282696 253904
rect 302332 253852 302384 253904
rect 282736 253784 282788 253836
rect 298376 253784 298428 253836
rect 282828 253716 282880 253768
rect 292580 253716 292632 253768
rect 282736 252492 282788 252544
rect 303712 252492 303764 252544
rect 282828 252424 282880 252476
rect 300952 252424 301004 252476
rect 282828 251132 282880 251184
rect 302424 251132 302476 251184
rect 309968 251132 310020 251184
rect 357532 251132 357584 251184
rect 502800 251132 502852 251184
rect 505100 251132 505152 251184
rect 282736 251064 282788 251116
rect 298100 251064 298152 251116
rect 282552 250996 282604 251048
rect 285680 250996 285732 251048
rect 308680 250452 308732 250504
rect 319720 250452 319772 250504
rect 282828 249704 282880 249756
rect 295524 249704 295576 249756
rect 282736 249636 282788 249688
rect 292764 249636 292816 249688
rect 282644 248072 282696 248124
rect 285864 248072 285916 248124
rect 282828 246984 282880 247036
rect 289912 246984 289964 247036
rect 322296 246984 322348 247036
rect 357532 246984 357584 247036
rect 321008 245556 321060 245608
rect 357532 245556 357584 245608
rect 299112 244876 299164 244928
rect 355692 244876 355744 244928
rect 530584 244876 530636 244928
rect 580172 244876 580224 244928
rect 50344 244196 50396 244248
rect 50712 244196 50764 244248
rect 323768 244196 323820 244248
rect 326344 244196 326396 244248
rect 319536 244128 319588 244180
rect 357532 244196 357584 244248
rect 305828 240048 305880 240100
rect 357532 240048 357584 240100
rect 81440 238688 81492 238740
rect 221740 238688 221792 238740
rect 282828 238688 282880 238740
rect 291476 238688 291528 238740
rect 88984 238620 89036 238672
rect 221648 238620 221700 238672
rect 97908 238552 97960 238604
rect 228456 238552 228508 238604
rect 86868 238484 86920 238536
rect 209228 238484 209280 238536
rect 88248 238416 88300 238468
rect 209320 238416 209372 238468
rect 102140 238348 102192 238400
rect 220176 238348 220228 238400
rect 104808 238280 104860 238332
rect 217508 238280 217560 238332
rect 99380 238212 99432 238264
rect 211988 238212 212040 238264
rect 106188 238144 106240 238196
rect 217416 238144 217468 238196
rect 98644 238076 98696 238128
rect 209136 238076 209188 238128
rect 108304 238008 108356 238060
rect 217324 238008 217376 238060
rect 281540 235900 281592 235952
rect 283748 235900 283800 235952
rect 293316 235900 293368 235952
rect 357532 235900 357584 235952
rect 189724 234540 189776 234592
rect 192484 234540 192536 234592
rect 314108 231752 314160 231804
rect 357532 231752 357584 231804
rect 294788 226244 294840 226296
rect 357716 226244 357768 226296
rect 311348 226176 311400 226228
rect 357532 226176 357584 226228
rect 296076 224884 296128 224936
rect 357532 224884 357584 224936
rect 290556 223524 290608 223576
rect 357532 223524 357584 223576
rect 307116 222096 307168 222148
rect 357716 222096 357768 222148
rect 336556 222028 336608 222080
rect 357532 222028 357584 222080
rect 308496 218016 308548 218068
rect 314660 218016 314712 218068
rect 287980 217948 288032 218000
rect 357532 217948 357584 218000
rect 327724 216588 327776 216640
rect 357532 216588 357584 216640
rect 303068 215228 303120 215280
rect 357532 215228 357584 215280
rect 3424 213936 3476 213988
rect 102784 213936 102836 213988
rect 298836 212440 298888 212492
rect 357532 212440 357584 212492
rect 319720 212372 319772 212424
rect 321928 212372 321980 212424
rect 314660 211760 314712 211812
rect 322388 211760 322440 211812
rect 320824 211080 320876 211132
rect 357532 211080 357584 211132
rect 314016 209720 314068 209772
rect 357532 209720 357584 209772
rect 102784 209040 102836 209092
rect 111708 209040 111760 209092
rect 289360 208292 289412 208344
rect 357532 208292 357584 208344
rect 192484 207000 192536 207052
rect 197360 207000 197412 207052
rect 289268 206932 289320 206984
rect 357532 206932 357584 206984
rect 334624 206864 334676 206916
rect 357532 206660 357584 206712
rect 529204 206252 529256 206304
rect 580172 206252 580224 206304
rect 289084 205572 289136 205624
rect 357532 205572 357584 205624
rect 313924 204212 313976 204264
rect 357532 204212 357584 204264
rect 321928 204144 321980 204196
rect 326436 204144 326488 204196
rect 326344 202784 326396 202836
rect 330484 202784 330536 202836
rect 197360 202104 197412 202156
rect 226064 202104 226116 202156
rect 322388 202104 322440 202156
rect 332508 202104 332560 202156
rect 294604 201424 294656 201476
rect 357532 201424 357584 201476
rect 311256 201356 311308 201408
rect 357532 201220 357584 201272
rect 326436 198704 326488 198756
rect 329104 198704 329156 198756
rect 332508 197956 332560 198008
rect 352932 197956 352984 198008
rect 287796 195916 287848 195968
rect 357532 195916 357584 195968
rect 226064 194488 226116 194540
rect 229928 194488 229980 194540
rect 282828 191836 282880 191888
rect 292580 191836 292632 191888
rect 351184 189728 351236 189780
rect 358268 189728 358320 189780
rect 329104 189048 329156 189100
rect 338028 189048 338080 189100
rect 38568 186940 38620 186992
rect 238392 186940 238444 186992
rect 111708 185580 111760 185632
rect 129096 185580 129148 185632
rect 54484 184900 54536 184952
rect 124220 184900 124272 184952
rect 124404 184900 124456 184952
rect 330484 184152 330536 184204
rect 351184 184152 351236 184204
rect 352932 184152 352984 184204
rect 359740 184152 359792 184204
rect 338028 181432 338080 181484
rect 358636 181432 358688 181484
rect 350172 180616 350224 180668
rect 379612 180616 379664 180668
rect 488448 180616 488500 180668
rect 522580 180616 522632 180668
rect 347136 180548 347188 180600
rect 380808 180548 380860 180600
rect 492496 180548 492548 180600
rect 525800 180548 525852 180600
rect 350356 180480 350408 180532
rect 384580 180480 384632 180532
rect 489552 180480 489604 180532
rect 523132 180480 523184 180532
rect 344560 180412 344612 180464
rect 382556 180412 382608 180464
rect 477408 180412 477460 180464
rect 521844 180412 521896 180464
rect 344468 180344 344520 180396
rect 383752 180344 383804 180396
rect 479432 180344 479484 180396
rect 527180 180344 527232 180396
rect 336464 180276 336516 180328
rect 381636 180276 381688 180328
rect 475384 180276 475436 180328
rect 523224 180276 523276 180328
rect 339040 180208 339092 180260
rect 385684 180208 385736 180260
rect 449072 180208 449124 180260
rect 524512 180208 524564 180260
rect 338764 180140 338816 180192
rect 386604 180140 386656 180192
rect 449808 180140 449860 180192
rect 536840 180140 536892 180192
rect 350264 180072 350316 180124
rect 377588 180072 377640 180124
rect 476120 180072 476172 180124
rect 480168 180072 480220 180124
rect 513472 180072 513524 180124
rect 355324 180004 355376 180056
rect 375564 180004 375616 180056
rect 358084 179936 358136 179988
rect 369492 179936 369544 179988
rect 491116 180004 491168 180056
rect 524420 180004 524472 180056
rect 503168 179936 503220 179988
rect 351184 179868 351236 179920
rect 367008 179868 367060 179920
rect 355416 179324 355468 179376
rect 423404 179324 423456 179376
rect 451740 179324 451792 179376
rect 539876 179324 539928 179376
rect 341800 179256 341852 179308
rect 409236 179256 409288 179308
rect 455788 179256 455840 179308
rect 543740 179256 543792 179308
rect 347504 179188 347556 179240
rect 408224 179188 408276 179240
rect 458824 179188 458876 179240
rect 545304 179188 545356 179240
rect 341524 179120 341576 179172
rect 402152 179120 402204 179172
rect 459836 179120 459888 179172
rect 545120 179120 545172 179172
rect 347412 179052 347464 179104
rect 407212 179052 407264 179104
rect 460848 179052 460900 179104
rect 543832 179052 543884 179104
rect 341708 178984 341760 179036
rect 396080 178984 396132 179036
rect 463884 178984 463936 179036
rect 545212 178984 545264 179036
rect 344376 178916 344428 178968
rect 398104 178916 398156 178968
rect 444656 178916 444708 178968
rect 520372 178916 520424 178968
rect 352748 178848 352800 178900
rect 406200 178848 406252 178900
rect 443644 178848 443696 178900
rect 519084 178848 519136 178900
rect 338856 178780 338908 178832
rect 390008 178780 390060 178832
rect 465908 178780 465960 178832
rect 541072 178780 541124 178832
rect 344284 178712 344336 178764
rect 395068 178712 395120 178764
rect 446680 178712 446732 178764
rect 521752 178712 521804 178764
rect 358268 178644 358320 178696
rect 369124 178644 369176 178696
rect 464896 178644 464948 178696
rect 538220 178644 538272 178696
rect 359740 178576 359792 178628
rect 369860 178576 369912 178628
rect 442632 178576 442684 178628
rect 501604 178576 501656 178628
rect 336004 178440 336056 178492
rect 373816 178440 373868 178492
rect 358636 178032 358688 178084
rect 347228 177964 347280 178016
rect 359648 177964 359700 178016
rect 366364 177964 366416 178016
rect 427452 177964 427504 178016
rect 472992 177964 473044 178016
rect 499580 177964 499632 178016
rect 355600 177896 355652 177948
rect 370780 177896 370832 177948
rect 467932 177896 467984 177948
rect 510620 177896 510672 177948
rect 365720 177828 365772 177880
rect 367008 177828 367060 177880
rect 376852 177828 376904 177880
rect 466920 177828 466972 177880
rect 509332 177828 509384 177880
rect 350080 177760 350132 177812
rect 404176 177760 404228 177812
rect 468944 177760 468996 177812
rect 507860 177760 507912 177812
rect 349988 177692 350040 177744
rect 403164 177692 403216 177744
rect 483112 177692 483164 177744
rect 518440 177692 518492 177744
rect 333244 177624 333296 177676
rect 368756 177624 368808 177676
rect 369860 177624 369912 177676
rect 419356 177624 419408 177676
rect 486148 177624 486200 177676
rect 520280 177624 520332 177676
rect 352656 177556 352708 177608
rect 401140 177556 401192 177608
rect 482100 177556 482152 177608
rect 516232 177556 516284 177608
rect 352564 177488 352616 177540
rect 400128 177488 400180 177540
rect 485136 177488 485188 177540
rect 518992 177488 519044 177540
rect 352840 177420 352892 177472
rect 399116 177420 399168 177472
rect 484124 177420 484176 177472
rect 517612 177420 517664 177472
rect 333336 177352 333388 177404
rect 367744 177352 367796 177404
rect 369124 177352 369176 177404
rect 412272 177352 412324 177404
rect 469956 177352 470008 177404
rect 502984 177352 503036 177404
rect 359464 177284 359516 177336
rect 388996 177284 389048 177336
rect 470968 177284 471020 177336
rect 503076 177284 503128 177336
rect 333428 177216 333480 177268
rect 378876 177216 378928 177268
rect 453764 177216 453816 177268
rect 540980 177216 541032 177268
rect 336280 177148 336332 177200
rect 394056 177148 394108 177200
rect 494244 177148 494296 177200
rect 518900 177148 518952 177200
rect 336188 177080 336240 177132
rect 397092 177080 397144 177132
rect 347320 176604 347372 176656
rect 417332 176604 417384 176656
rect 426440 176604 426492 176656
rect 513380 176604 513432 176656
rect 347044 176536 347096 176588
rect 393044 176536 393096 176588
rect 445668 176536 445720 176588
rect 531320 176536 531372 176588
rect 452752 176468 452804 176520
rect 528560 176468 528612 176520
rect 429476 176400 429528 176452
rect 505284 176400 505336 176452
rect 440608 176332 440660 176384
rect 516140 176332 516192 176384
rect 434536 176264 434588 176316
rect 509240 176264 509292 176316
rect 305644 175924 305696 175976
rect 371056 175924 371108 175976
rect 416320 175176 416372 175228
rect 505192 175176 505244 175228
rect 430488 175108 430540 175160
rect 517704 175108 517756 175160
rect 447692 175040 447744 175092
rect 523960 175040 524012 175092
rect 436560 174972 436612 175024
rect 511356 174972 511408 175024
rect 450728 174904 450780 174956
rect 512644 174904 512696 174956
rect 308404 170348 308456 170400
rect 372252 170348 372304 170400
rect 282828 169736 282880 169788
rect 290004 169736 290056 169788
rect 360108 169260 360160 169312
rect 393780 169260 393832 169312
rect 315304 169192 315356 169244
rect 377036 169192 377088 169244
rect 349988 169124 350040 169176
rect 580264 169124 580316 169176
rect 349804 169056 349856 169108
rect 580356 169056 580408 169108
rect 349896 168988 349948 169040
rect 580540 168988 580592 169040
rect 282828 168376 282880 168428
rect 290096 168376 290148 168428
rect 282460 168308 282512 168360
rect 291200 168308 291252 168360
rect 282644 167016 282696 167068
rect 289820 167016 289872 167068
rect 282828 166948 282880 167000
rect 303620 166948 303672 167000
rect 524328 166948 524380 167000
rect 580172 166948 580224 167000
rect 282828 165520 282880 165572
rect 296812 165520 296864 165572
rect 302884 164840 302936 164892
rect 368664 164840 368716 164892
rect 3424 164160 3476 164212
rect 54484 164160 54536 164212
rect 282828 164160 282880 164212
rect 296720 164160 296772 164212
rect 282644 164092 282696 164144
rect 295340 164092 295392 164144
rect 282644 162800 282696 162852
rect 302240 162800 302292 162852
rect 282828 162732 282880 162784
rect 288440 162732 288492 162784
rect 324964 162120 325016 162172
rect 384212 162120 384264 162172
rect 282828 161372 282880 161424
rect 290188 161372 290240 161424
rect 309784 160692 309836 160744
rect 373448 160692 373500 160744
rect 229836 155864 229888 155916
rect 237380 155864 237432 155916
rect 229928 154504 229980 154556
rect 237380 154504 237432 154556
rect 318156 151784 318208 151836
rect 580172 151784 580224 151836
rect 311164 149676 311216 149728
rect 374644 149676 374696 149728
rect 322204 148384 322256 148436
rect 381820 148384 381872 148436
rect 319444 148316 319496 148368
rect 380624 148316 380676 148368
rect 358728 146956 358780 147008
rect 363604 146956 363656 147008
rect 355968 146888 356020 146940
rect 364984 146888 365036 146940
rect 355416 146752 355468 146804
rect 362868 146752 362920 146804
rect 352656 146684 352708 146736
rect 365904 146684 365956 146736
rect 358176 146616 358228 146668
rect 388996 146616 389048 146668
rect 358268 146548 358320 146600
rect 390192 146548 390244 146600
rect 359556 146480 359608 146532
rect 392584 146480 392636 146532
rect 355600 146412 355652 146464
rect 362776 146412 362828 146464
rect 362868 146412 362920 146464
rect 391388 146412 391440 146464
rect 359464 146344 359516 146396
rect 397368 146344 397420 146396
rect 355876 146276 355928 146328
rect 362684 146276 362736 146328
rect 362776 146276 362828 146328
rect 398564 146276 398616 146328
rect 358360 144440 358412 144492
rect 386420 144440 386472 144492
rect 358636 144372 358688 144424
rect 385132 144372 385184 144424
rect 359648 144304 359700 144356
rect 407764 144304 407816 144356
rect 358452 144236 358504 144288
rect 387708 144236 387760 144288
rect 238392 122000 238444 122052
rect 239956 122000 240008 122052
rect 235816 120640 235868 120692
rect 283196 120640 283248 120692
rect 235908 120572 235960 120624
rect 355600 120572 355652 120624
rect 279976 120504 280028 120556
rect 290096 120504 290148 120556
rect 50252 120028 50304 120080
rect 63500 120028 63552 120080
rect 126980 120028 127032 120080
rect 129004 120028 129056 120080
rect 129924 120028 129976 120080
rect 358636 120028 358688 120080
rect 50620 119960 50672 120012
rect 61476 119960 61528 120012
rect 127624 119960 127676 120012
rect 350080 119960 350132 120012
rect 127532 119892 127584 119944
rect 289820 119892 289872 119944
rect 127808 119824 127860 119876
rect 284300 119824 284352 119876
rect 128084 119756 128136 119808
rect 283104 119756 283156 119808
rect 127808 119688 127860 119740
rect 129924 119688 129976 119740
rect 238576 119688 238628 119740
rect 358544 119688 358596 119740
rect 238300 119620 238352 119672
rect 318156 119620 318208 119672
rect 235816 119552 235868 119604
rect 284576 119552 284628 119604
rect 235908 119484 235960 119536
rect 284392 119484 284444 119536
rect 238576 119416 238628 119468
rect 284484 119416 284536 119468
rect 49516 118600 49568 118652
rect 72332 118600 72384 118652
rect 109040 118600 109092 118652
rect 125692 118600 125744 118652
rect 234620 118600 234672 118652
rect 245752 118600 245804 118652
rect 247040 118600 247092 118652
rect 250076 118600 250128 118652
rect 50528 118532 50580 118584
rect 84568 118532 84620 118584
rect 114284 118532 114336 118584
rect 125784 118532 125836 118584
rect 126888 118532 126940 118584
rect 237564 118532 237616 118584
rect 246580 118532 246632 118584
rect 48044 118464 48096 118516
rect 81072 118464 81124 118516
rect 116032 118464 116084 118516
rect 129096 118464 129148 118516
rect 132500 118464 132552 118516
rect 359556 118464 359608 118516
rect 49608 118396 49660 118448
rect 79324 118396 79376 118448
rect 102048 118396 102100 118448
rect 117688 118396 117740 118448
rect 117780 118396 117832 118448
rect 124404 118396 124456 118448
rect 125232 118396 125284 118448
rect 47952 118328 48004 118380
rect 77576 118328 77628 118380
rect 103796 118328 103848 118380
rect 128544 118328 128596 118380
rect 48136 118260 48188 118312
rect 75828 118260 75880 118312
rect 107292 118260 107344 118312
rect 239956 118396 240008 118448
rect 349804 118396 349856 118448
rect 238208 118328 238260 118380
rect 359648 118328 359700 118380
rect 238484 118260 238536 118312
rect 349988 118260 350040 118312
rect 105544 118192 105596 118244
rect 129832 118192 129884 118244
rect 238024 118192 238076 118244
rect 349896 118192 349948 118244
rect 110788 118124 110840 118176
rect 132592 118124 132644 118176
rect 237380 118124 237432 118176
rect 248972 118124 249024 118176
rect 264980 118124 265032 118176
rect 294052 118124 294104 118176
rect 112536 118056 112588 118108
rect 131212 118056 131264 118108
rect 131488 118056 131540 118108
rect 237472 118056 237524 118108
rect 247684 118056 247736 118108
rect 271788 118056 271840 118108
rect 292672 118056 292724 118108
rect 117688 117988 117740 118040
rect 124220 117988 124272 118040
rect 125508 117988 125560 118040
rect 126888 117988 126940 118040
rect 359464 117988 359516 118040
rect 61844 117920 61896 117972
rect 360660 117920 360712 117972
rect 89812 117852 89864 117904
rect 124864 117852 124916 117904
rect 91560 117784 91612 117836
rect 125600 117784 125652 117836
rect 121460 117716 121512 117768
rect 244280 117716 244332 117768
rect 45376 117240 45428 117292
rect 67548 117240 67600 117292
rect 128544 117240 128596 117292
rect 358268 117240 358320 117292
rect 46756 117172 46808 117224
rect 65340 117172 65392 117224
rect 66168 117172 66220 117224
rect 107568 117172 107620 117224
rect 129740 117172 129792 117224
rect 358360 117172 358412 117224
rect 106188 117104 106240 117156
rect 131120 117104 131172 117156
rect 358452 117104 358504 117156
rect 191748 117036 191800 117088
rect 355416 117036 355468 117088
rect 212448 116968 212500 117020
rect 358176 116968 358228 117020
rect 241428 116900 241480 116952
rect 352656 116900 352708 116952
rect 66168 115880 66220 115932
rect 295984 115880 296036 115932
rect 67548 115812 67600 115864
rect 297364 115812 297416 115864
rect 234620 115744 234672 115796
rect 355968 115744 356020 115796
rect 358084 115744 358136 115796
rect 252468 114452 252520 114504
rect 290004 114452 290056 114504
rect 360660 88952 360712 89004
rect 537484 88952 537536 89004
rect 73068 87252 73120 87304
rect 91744 87252 91796 87304
rect 74448 87184 74500 87236
rect 86316 87184 86368 87236
rect 76472 87116 76524 87168
rect 90548 87116 90600 87168
rect 84016 87048 84068 87100
rect 98736 87048 98788 87100
rect 358084 86912 358136 86964
rect 580172 86912 580224 86964
rect 86316 69640 86368 69692
rect 350448 69640 350500 69692
rect 91744 54476 91796 54528
rect 346952 54476 347004 54528
rect 90548 50328 90600 50380
rect 354036 50328 354088 50380
rect 537484 46860 537536 46912
rect 580172 46860 580224 46912
rect 98736 10276 98788 10328
rect 371700 10276 371752 10328
rect 331864 6808 331916 6860
rect 580172 6808 580224 6860
rect 271788 4088 271840 4140
rect 292580 4088 292632 4140
rect 446404 3408 446456 3460
rect 583392 3408 583444 3460
rect 442908 2796 442960 2848
rect 581000 2796 581052 2848
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 579698 3464 579935
rect 3424 579692 3476 579698
rect 3424 579634 3476 579640
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 4066 398168 4122 398177
rect 4066 398103 4122 398112
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 4080 358737 4108 398103
rect 4066 358728 4122 358737
rect 4066 358663 4122 358672
rect 3424 319456 3476 319462
rect 3424 319398 3476 319404
rect 3436 319297 3464 319398
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 8128 312497 8156 703520
rect 24320 700369 24348 703520
rect 24306 700360 24362 700369
rect 24306 700295 24362 700304
rect 31022 700360 31078 700369
rect 31022 700295 31078 700304
rect 26148 683188 26200 683194
rect 26148 683130 26200 683136
rect 25686 645144 25742 645153
rect 25686 645079 25742 645088
rect 25502 542872 25558 542881
rect 25502 542807 25558 542816
rect 11704 474768 11756 474774
rect 11704 474710 11756 474716
rect 11716 388482 11744 474710
rect 25516 432313 25544 542807
rect 25596 523116 25648 523122
rect 25596 523058 25648 523064
rect 25502 432304 25558 432313
rect 25502 432239 25558 432248
rect 14464 422340 14516 422346
rect 14464 422282 14516 422288
rect 14476 390250 14504 422282
rect 14464 390244 14516 390250
rect 14464 390186 14516 390192
rect 11704 388476 11756 388482
rect 11704 388418 11756 388424
rect 25608 360942 25636 523058
rect 25700 481273 25728 645079
rect 25870 644192 25926 644201
rect 25870 644127 25926 644136
rect 25780 526108 25832 526114
rect 25780 526050 25832 526056
rect 25686 481264 25742 481273
rect 25686 481199 25742 481208
rect 25792 361078 25820 526050
rect 25884 475833 25912 644127
rect 26054 643240 26110 643249
rect 26054 643175 26110 643184
rect 25964 528624 26016 528630
rect 25964 528566 26016 528572
rect 25870 475824 25926 475833
rect 25870 475759 25926 475768
rect 25780 361072 25832 361078
rect 25780 361014 25832 361020
rect 25976 361010 26004 528566
rect 26068 471481 26096 643175
rect 26054 471472 26110 471481
rect 26054 471407 26110 471416
rect 26160 387122 26188 683130
rect 27434 655072 27490 655081
rect 27434 655007 27490 655016
rect 26790 654256 26846 654265
rect 26790 654191 26846 654200
rect 26804 393689 26832 654191
rect 27250 549672 27306 549681
rect 27250 549607 27306 549616
rect 26974 538520 27030 538529
rect 26974 538455 27030 538464
rect 26884 523524 26936 523530
rect 26884 523466 26936 523472
rect 26896 479534 26924 523466
rect 26884 479528 26936 479534
rect 26884 479470 26936 479476
rect 26988 420889 27016 538455
rect 27066 534168 27122 534177
rect 27066 534103 27122 534112
rect 26974 420880 27030 420889
rect 26974 420815 27030 420824
rect 27080 400761 27108 534103
rect 27160 522300 27212 522306
rect 27160 522242 27212 522248
rect 27066 400752 27122 400761
rect 27066 400687 27122 400696
rect 26790 393680 26846 393689
rect 26790 393615 26846 393624
rect 27172 387190 27200 522242
rect 27264 410553 27292 549607
rect 27344 524612 27396 524618
rect 27344 524554 27396 524560
rect 27250 410544 27306 410553
rect 27250 410479 27306 410488
rect 27160 387184 27212 387190
rect 27160 387126 27212 387132
rect 26148 387116 26200 387122
rect 26148 387058 26200 387064
rect 25964 361004 26016 361010
rect 25964 360946 26016 360952
rect 25596 360936 25648 360942
rect 25596 360878 25648 360884
rect 27356 352578 27384 524554
rect 27448 395865 27476 655007
rect 30194 654528 30250 654537
rect 30194 654463 30250 654472
rect 28262 652896 28318 652905
rect 28262 652831 28318 652840
rect 27528 523728 27580 523734
rect 27528 523670 27580 523676
rect 27540 497486 27568 523670
rect 27528 497480 27580 497486
rect 27528 497422 27580 497428
rect 27434 395856 27490 395865
rect 27434 395791 27490 395800
rect 28276 394233 28304 652831
rect 30010 641336 30066 641345
rect 30010 641271 30066 641280
rect 28538 638616 28594 638625
rect 28538 638551 28594 638560
rect 28446 553072 28502 553081
rect 28446 553007 28502 553016
rect 28354 544096 28410 544105
rect 28354 544031 28410 544040
rect 28368 408921 28396 544031
rect 28460 410009 28488 553007
rect 28552 467673 28580 638551
rect 28722 633992 28778 634001
rect 28722 633927 28778 633936
rect 28632 523252 28684 523258
rect 28632 523194 28684 523200
rect 28538 467664 28594 467673
rect 28538 467599 28594 467608
rect 28446 410000 28502 410009
rect 28446 409935 28502 409944
rect 28354 408912 28410 408921
rect 28354 408847 28410 408856
rect 28262 394224 28318 394233
rect 28262 394159 28318 394168
rect 28644 352646 28672 523194
rect 28736 461145 28764 633927
rect 28814 633856 28870 633865
rect 28814 633791 28870 633800
rect 28722 461136 28778 461145
rect 28722 461071 28778 461080
rect 28828 460601 28856 633791
rect 29920 525020 29972 525026
rect 29920 524962 29972 524968
rect 29828 524748 29880 524754
rect 29828 524690 29880 524696
rect 29736 523320 29788 523326
rect 29736 523262 29788 523268
rect 28908 519580 28960 519586
rect 28908 519522 28960 519528
rect 28920 496806 28948 519522
rect 28908 496800 28960 496806
rect 28908 496742 28960 496748
rect 28814 460592 28870 460601
rect 28814 460527 28870 460536
rect 29748 366586 29776 523262
rect 29736 366580 29788 366586
rect 29736 366522 29788 366528
rect 29840 366518 29868 524690
rect 29828 366512 29880 366518
rect 29828 366454 29880 366460
rect 29932 363934 29960 524962
rect 30024 468217 30052 641271
rect 30102 542328 30158 542337
rect 30102 542263 30158 542272
rect 30010 468208 30066 468217
rect 30010 468143 30066 468152
rect 29920 363928 29972 363934
rect 29920 363870 29972 363876
rect 28632 352640 28684 352646
rect 28632 352582 28684 352588
rect 27344 352572 27396 352578
rect 27344 352514 27396 352520
rect 30116 350441 30144 542263
rect 30208 390969 30236 654463
rect 30286 654392 30342 654401
rect 30286 654327 30342 654336
rect 30300 391513 30328 654327
rect 30286 391504 30342 391513
rect 30286 391439 30342 391448
rect 30194 390960 30250 390969
rect 30194 390895 30250 390904
rect 31036 354385 31064 700295
rect 40512 699718 40540 703520
rect 43074 700360 43130 700369
rect 43074 700295 43130 700304
rect 40500 699712 40552 699718
rect 40500 699654 40552 699660
rect 41420 699712 41472 699718
rect 41420 699654 41472 699660
rect 33046 654664 33102 654673
rect 33046 654599 33102 654608
rect 31666 651672 31722 651681
rect 31666 651607 31722 651616
rect 31298 642424 31354 642433
rect 31298 642359 31354 642368
rect 31206 532944 31262 532953
rect 31206 532879 31262 532888
rect 31114 525192 31170 525201
rect 31114 525127 31170 525136
rect 31128 503713 31156 525127
rect 31114 503704 31170 503713
rect 31114 503639 31170 503648
rect 31220 420345 31248 532879
rect 31312 480729 31340 642359
rect 31576 632120 31628 632126
rect 31576 632062 31628 632068
rect 31484 524680 31536 524686
rect 31484 524622 31536 524628
rect 31390 514856 31446 514865
rect 31390 514791 31446 514800
rect 31298 480720 31354 480729
rect 31298 480655 31354 480664
rect 31206 420336 31262 420345
rect 31206 420271 31262 420280
rect 31404 354521 31432 514791
rect 31390 354512 31446 354521
rect 31390 354447 31446 354456
rect 31022 354376 31078 354385
rect 31022 354311 31078 354320
rect 30102 350432 30158 350441
rect 30102 350367 30158 350376
rect 31496 347070 31524 524622
rect 31588 387258 31616 632062
rect 31680 393145 31708 651607
rect 32862 642016 32918 642025
rect 32862 641951 32918 641960
rect 32678 539880 32734 539889
rect 32678 539815 32734 539824
rect 32586 535664 32642 535673
rect 32586 535599 32642 535608
rect 31760 527876 31812 527882
rect 31760 527818 31812 527824
rect 31772 527202 31800 527818
rect 31760 527196 31812 527202
rect 31760 527138 31812 527144
rect 32494 526960 32550 526969
rect 32494 526895 32550 526904
rect 32402 523424 32458 523433
rect 32402 523359 32458 523368
rect 32416 498681 32444 523359
rect 32402 498672 32458 498681
rect 32402 498607 32458 498616
rect 31852 496800 31904 496806
rect 31852 496742 31904 496748
rect 31864 494018 31892 496742
rect 31852 494012 31904 494018
rect 31852 493954 31904 493960
rect 32508 427417 32536 526895
rect 32494 427408 32550 427417
rect 32494 427343 32550 427352
rect 32600 421977 32628 535599
rect 32692 423065 32720 539815
rect 32772 527876 32824 527882
rect 32772 527818 32824 527824
rect 32678 423056 32734 423065
rect 32678 422991 32734 423000
rect 32586 421968 32642 421977
rect 32586 421903 32642 421912
rect 31666 393136 31722 393145
rect 31666 393071 31722 393080
rect 32784 387530 32812 527818
rect 32876 469305 32904 641951
rect 32954 638072 33010 638081
rect 32954 638007 33010 638016
rect 32862 469296 32918 469305
rect 32862 469231 32918 469240
rect 32968 464953 32996 638007
rect 32954 464944 33010 464953
rect 32954 464879 33010 464888
rect 33060 392057 33088 654599
rect 41326 653712 41382 653721
rect 41326 653647 41382 653656
rect 33782 653032 33838 653041
rect 33782 652967 33838 652976
rect 33796 392601 33824 652967
rect 39670 651128 39726 651137
rect 39670 651063 39726 651072
rect 35714 640520 35770 640529
rect 35714 640455 35770 640464
rect 34334 640112 34390 640121
rect 34334 640047 34390 640056
rect 34242 553752 34298 553761
rect 34242 553687 34298 553696
rect 33874 546816 33930 546825
rect 33874 546751 33930 546760
rect 33888 504665 33916 546751
rect 34150 542464 34206 542473
rect 34150 542399 34206 542408
rect 34058 533760 34114 533769
rect 34058 533695 34114 533704
rect 33966 530768 34022 530777
rect 33966 530703 34022 530712
rect 33874 504656 33930 504665
rect 33874 504591 33930 504600
rect 33980 401305 34008 530703
rect 33966 401296 34022 401305
rect 33966 401231 34022 401240
rect 34072 398585 34100 533695
rect 34164 399129 34192 542399
rect 34256 408377 34284 553687
rect 34348 467129 34376 640047
rect 35622 549536 35678 549545
rect 35622 549471 35678 549480
rect 35530 546000 35586 546009
rect 35530 545935 35586 545944
rect 35254 538656 35310 538665
rect 35254 538591 35310 538600
rect 35162 526552 35218 526561
rect 35162 526487 35218 526496
rect 34428 520940 34480 520946
rect 34428 520882 34480 520888
rect 34440 495514 34468 520882
rect 34428 495508 34480 495514
rect 34428 495450 34480 495456
rect 35072 495508 35124 495514
rect 35072 495450 35124 495456
rect 35084 467158 35112 495450
rect 35072 467152 35124 467158
rect 34334 467120 34390 467129
rect 35072 467094 35124 467100
rect 34334 467055 34390 467064
rect 35176 421433 35204 526487
rect 35268 426873 35296 538591
rect 35346 537024 35402 537033
rect 35346 536959 35402 536968
rect 35254 426864 35310 426873
rect 35254 426799 35310 426808
rect 35162 421424 35218 421433
rect 35162 421359 35218 421368
rect 35360 412185 35388 536959
rect 35438 524648 35494 524657
rect 35438 524583 35494 524592
rect 35346 412176 35402 412185
rect 35346 412111 35402 412120
rect 34242 408368 34298 408377
rect 34242 408303 34298 408312
rect 35452 400217 35480 524583
rect 35438 400208 35494 400217
rect 35438 400143 35494 400152
rect 35544 399673 35572 545935
rect 35530 399664 35586 399673
rect 35530 399599 35586 399608
rect 34150 399120 34206 399129
rect 34150 399055 34206 399064
rect 34058 398576 34114 398585
rect 34058 398511 34114 398520
rect 35636 398041 35664 549471
rect 35728 480185 35756 640455
rect 37186 639296 37242 639305
rect 37186 639231 37242 639240
rect 35806 638208 35862 638217
rect 35806 638143 35862 638152
rect 35714 480176 35770 480185
rect 35714 480111 35770 480120
rect 35622 398032 35678 398041
rect 35622 397967 35678 397976
rect 35820 395321 35848 638143
rect 36634 557832 36690 557841
rect 36634 557767 36690 557776
rect 36542 533080 36598 533089
rect 36542 533015 36598 533024
rect 36556 413273 36584 533015
rect 36648 429593 36676 557767
rect 37096 557592 37148 557598
rect 37096 557534 37148 557540
rect 37002 551032 37058 551041
rect 37002 550967 37058 550976
rect 36910 545320 36966 545329
rect 36910 545255 36966 545264
rect 36818 543960 36874 543969
rect 36818 543895 36874 543904
rect 36726 539744 36782 539753
rect 36726 539679 36782 539688
rect 36634 429584 36690 429593
rect 36634 429519 36690 429528
rect 36542 413264 36598 413273
rect 36542 413199 36598 413208
rect 36740 404025 36768 539679
rect 36726 404016 36782 404025
rect 36726 403951 36782 403960
rect 36832 403481 36860 543895
rect 36818 403472 36874 403481
rect 36818 403407 36874 403416
rect 36924 402937 36952 545255
rect 37016 405113 37044 550967
rect 37002 405104 37058 405113
rect 37002 405039 37058 405048
rect 36910 402928 36966 402937
rect 36910 402863 36966 402872
rect 35806 395312 35862 395321
rect 35806 395247 35862 395256
rect 33782 392592 33838 392601
rect 33782 392527 33838 392536
rect 33046 392048 33102 392057
rect 33046 391983 33102 391992
rect 37108 387598 37136 557534
rect 37200 462777 37228 639231
rect 38568 635520 38620 635526
rect 38568 635462 38620 635468
rect 38474 635080 38530 635089
rect 38474 635015 38530 635024
rect 38106 552392 38162 552401
rect 38106 552327 38162 552336
rect 37922 531992 37978 532001
rect 37922 531927 37978 531936
rect 37936 504121 37964 531927
rect 38014 523696 38070 523705
rect 38014 523631 38070 523640
rect 37922 504112 37978 504121
rect 37922 504047 37978 504056
rect 37922 503704 37978 503713
rect 37922 503639 37978 503648
rect 37936 491881 37964 503639
rect 37922 491872 37978 491881
rect 37922 491807 37978 491816
rect 38028 488889 38056 523631
rect 38120 506297 38148 552327
rect 38382 547904 38438 547913
rect 38382 547839 38438 547848
rect 38198 541240 38254 541249
rect 38198 541175 38254 541184
rect 38106 506288 38162 506297
rect 38106 506223 38162 506232
rect 38108 494012 38160 494018
rect 38108 493954 38160 493960
rect 38014 488880 38070 488889
rect 38014 488815 38070 488824
rect 37924 479528 37976 479534
rect 37924 479470 37976 479476
rect 37186 462768 37242 462777
rect 37186 462703 37242 462712
rect 37936 392630 37964 479470
rect 38120 478174 38148 493954
rect 38108 478168 38160 478174
rect 38108 478110 38160 478116
rect 38212 404569 38240 541175
rect 38290 534984 38346 534993
rect 38290 534919 38346 534928
rect 38198 404560 38254 404569
rect 38198 404495 38254 404504
rect 38304 396953 38332 534919
rect 38396 406201 38424 547839
rect 38488 477465 38516 635015
rect 38474 477456 38530 477465
rect 38474 477391 38530 477400
rect 38382 406192 38438 406201
rect 38382 406127 38438 406136
rect 38290 396944 38346 396953
rect 38290 396879 38346 396888
rect 37924 392624 37976 392630
rect 37924 392566 37976 392572
rect 37096 387592 37148 387598
rect 37096 387534 37148 387540
rect 32772 387524 32824 387530
rect 32772 387466 32824 387472
rect 31576 387252 31628 387258
rect 31576 387194 31628 387200
rect 31484 347064 31536 347070
rect 31484 347006 31536 347012
rect 8114 312488 8170 312497
rect 8114 312423 8170 312432
rect 3424 267708 3476 267714
rect 3424 267650 3476 267656
rect 3436 267209 3464 267650
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3436 213994 3464 214911
rect 35162 214160 35218 214169
rect 35162 214095 35218 214104
rect 3424 213988 3476 213994
rect 3424 213930 3476 213936
rect 5262 213072 5318 213081
rect 5262 213007 5318 213016
rect 3424 164212 3476 164218
rect 3424 164154 3476 164160
rect 3436 162897 3464 164154
rect 3422 162888 3478 162897
rect 3422 162823 3478 162832
rect 570 46200 626 46209
rect 570 46135 626 46144
rect 584 480 612 46135
rect 4066 17232 4122 17241
rect 4066 17167 4122 17176
rect 2870 8936 2926 8945
rect 2870 8871 2926 8880
rect 1674 5264 1730 5273
rect 1674 5199 1730 5208
rect 1688 480 1716 5199
rect 2884 480 2912 8871
rect 4080 480 4108 17167
rect 5276 480 5304 213007
rect 31022 211984 31078 211993
rect 31022 211919 31078 211928
rect 6458 210896 6514 210905
rect 6458 210831 6514 210840
rect 6472 480 6500 210831
rect 21822 118144 21878 118153
rect 21822 118079 21878 118088
rect 7562 115968 7618 115977
rect 7562 115903 7618 115912
rect 7576 71641 7604 115903
rect 13542 112704 13598 112713
rect 13542 112639 13598 112648
rect 9954 104136 10010 104145
rect 9954 104071 10010 104080
rect 7562 71632 7618 71641
rect 7562 71567 7618 71576
rect 8758 20224 8814 20233
rect 8758 20159 8814 20168
rect 7654 3496 7710 3505
rect 7654 3431 7710 3440
rect 7668 480 7696 3431
rect 8772 480 8800 20159
rect 9968 480 9996 104071
rect 11702 100056 11758 100065
rect 11702 99991 11758 100000
rect 11716 3505 11744 99991
rect 12346 6216 12402 6225
rect 12346 6151 12402 6160
rect 11702 3496 11758 3505
rect 11702 3431 11758 3440
rect 12360 480 12388 6151
rect 13556 480 13584 112639
rect 18234 109848 18290 109857
rect 18234 109783 18290 109792
rect 14738 98832 14794 98841
rect 14738 98767 14794 98776
rect 14752 480 14780 98767
rect 17038 3496 17094 3505
rect 17038 3431 17094 3440
rect 17052 480 17080 3431
rect 18248 480 18276 109783
rect 18602 106992 18658 107001
rect 18602 106927 18658 106936
rect 18616 3505 18644 106927
rect 18602 3496 18658 3505
rect 18602 3431 18658 3440
rect 19430 2816 19486 2825
rect 19430 2751 19486 2760
rect 19444 480 19472 2751
rect 21836 480 21864 118079
rect 30102 117464 30158 117473
rect 30102 117399 30158 117408
rect 26514 117328 26570 117337
rect 26514 117263 26570 117272
rect 24214 94480 24270 94489
rect 24214 94415 24270 94424
rect 23018 93392 23074 93401
rect 23018 93327 23074 93336
rect 23032 480 23060 93327
rect 24228 480 24256 94415
rect 26528 480 26556 117263
rect 28906 89040 28962 89049
rect 28906 88975 28962 88984
rect 27710 16144 27766 16153
rect 27710 16079 27766 16088
rect 27724 480 27752 16079
rect 28920 480 28948 88975
rect 30116 480 30144 117399
rect 31036 17241 31064 211919
rect 33598 117736 33654 117745
rect 33598 117671 33654 117680
rect 32402 109712 32458 109721
rect 32402 109647 32458 109656
rect 31022 17232 31078 17241
rect 31022 17167 31078 17176
rect 31298 6352 31354 6361
rect 31298 6287 31354 6296
rect 31312 480 31340 6287
rect 32416 480 32444 109647
rect 33612 480 33640 117671
rect 34794 97200 34850 97209
rect 34794 97135 34850 97144
rect 34808 480 34836 97135
rect 35176 8945 35204 214095
rect 38580 186998 38608 635462
rect 39486 558240 39542 558249
rect 39486 558175 39542 558184
rect 39210 552664 39266 552673
rect 39210 552599 39266 552608
rect 39224 507929 39252 552599
rect 39394 527368 39450 527377
rect 39394 527303 39450 527312
rect 39302 521248 39358 521257
rect 39302 521183 39358 521192
rect 39210 507920 39266 507929
rect 39210 507855 39266 507864
rect 39316 397497 39344 521183
rect 39408 402393 39436 527303
rect 39500 431769 39528 558175
rect 39578 535528 39634 535537
rect 39578 535463 39634 535472
rect 39486 431760 39542 431769
rect 39486 431695 39542 431704
rect 39394 402384 39450 402393
rect 39394 402319 39450 402328
rect 39302 397488 39358 397497
rect 39302 397423 39358 397432
rect 39592 396409 39620 535463
rect 39684 502353 39712 651063
rect 39762 650992 39818 651001
rect 39762 650927 39818 650936
rect 39670 502344 39726 502353
rect 39670 502279 39726 502288
rect 39776 494737 39804 650927
rect 39854 650720 39910 650729
rect 39854 650655 39910 650664
rect 39762 494728 39818 494737
rect 39762 494663 39818 494672
rect 39868 491201 39896 650655
rect 40774 650448 40830 650457
rect 40774 650383 40830 650392
rect 40682 536888 40738 536897
rect 40682 536823 40738 536832
rect 40498 532808 40554 532817
rect 40498 532743 40554 532752
rect 39948 526040 40000 526046
rect 39948 525982 40000 525988
rect 39854 491192 39910 491201
rect 39854 491127 39910 491136
rect 39578 396400 39634 396409
rect 39578 396335 39634 396344
rect 39960 363866 39988 525982
rect 40512 419257 40540 532743
rect 40590 530088 40646 530097
rect 40590 530023 40646 530032
rect 40498 419248 40554 419257
rect 40498 419183 40554 419192
rect 40604 405657 40632 530023
rect 40590 405648 40646 405657
rect 40590 405583 40646 405592
rect 40696 401849 40724 536823
rect 40788 506569 40816 650383
rect 41234 648952 41290 648961
rect 41234 648887 41290 648896
rect 40960 525972 41012 525978
rect 40960 525914 41012 525920
rect 40868 520736 40920 520742
rect 40868 520678 40920 520684
rect 40774 506560 40830 506569
rect 40774 506495 40830 506504
rect 40682 401840 40738 401849
rect 40682 401775 40738 401784
rect 39948 363860 40000 363866
rect 39948 363802 40000 363808
rect 40880 359514 40908 520678
rect 40972 364070 41000 525914
rect 41052 524816 41104 524822
rect 41052 524758 41104 524764
rect 40960 364064 41012 364070
rect 40960 364006 41012 364012
rect 41064 361146 41092 524758
rect 41144 521212 41196 521218
rect 41144 521154 41196 521160
rect 41052 361140 41104 361146
rect 41052 361082 41104 361088
rect 40868 359508 40920 359514
rect 40868 359450 40920 359456
rect 41156 349858 41184 521154
rect 41248 473113 41276 648887
rect 41234 473104 41290 473113
rect 41234 473039 41290 473048
rect 41340 461689 41368 653647
rect 41432 522306 41460 699654
rect 42154 650584 42210 650593
rect 42154 650519 42210 650528
rect 41512 579692 41564 579698
rect 41512 579634 41564 579640
rect 41524 557666 41552 579634
rect 42062 557968 42118 557977
rect 42062 557903 42118 557912
rect 41512 557660 41564 557666
rect 41512 557602 41564 557608
rect 41878 530632 41934 530641
rect 41878 530567 41934 530576
rect 41420 522300 41472 522306
rect 41420 522242 41472 522248
rect 41892 509017 41920 530567
rect 41970 520704 42026 520713
rect 41970 520639 42026 520648
rect 41878 509008 41934 509017
rect 41878 508943 41934 508952
rect 41326 461680 41382 461689
rect 41326 461615 41382 461624
rect 41984 419801 42012 520639
rect 42076 435033 42104 557903
rect 42168 498137 42196 650519
rect 42706 650312 42762 650321
rect 42706 650247 42762 650256
rect 42522 642152 42578 642161
rect 42522 642087 42578 642096
rect 42432 523388 42484 523394
rect 42432 523330 42484 523336
rect 42340 522640 42392 522646
rect 42340 522582 42392 522588
rect 42248 520872 42300 520878
rect 42248 520814 42300 520820
rect 42154 498128 42210 498137
rect 42154 498063 42210 498072
rect 42062 435024 42118 435033
rect 42062 434959 42118 434968
rect 41970 419792 42026 419801
rect 41970 419727 42026 419736
rect 42260 366382 42288 520814
rect 42248 366376 42300 366382
rect 42248 366318 42300 366324
rect 42352 363730 42380 522582
rect 42444 364138 42472 523330
rect 42536 479097 42564 642087
rect 42616 521824 42668 521830
rect 42616 521766 42668 521772
rect 42522 479088 42578 479097
rect 42522 479023 42578 479032
rect 42432 364132 42484 364138
rect 42432 364074 42484 364080
rect 42340 363724 42392 363730
rect 42340 363666 42392 363672
rect 42628 350130 42656 521766
rect 42720 469849 42748 650247
rect 42706 469840 42762 469849
rect 42706 469775 42762 469784
rect 43088 353297 43116 700295
rect 45468 658300 45520 658306
rect 45468 658242 45520 658248
rect 43994 647592 44050 647601
rect 43994 647527 44050 647536
rect 43902 582176 43958 582185
rect 43902 582111 43958 582120
rect 43442 558104 43498 558113
rect 43442 558039 43498 558048
rect 43166 548040 43222 548049
rect 43166 547975 43222 547984
rect 43180 496097 43208 547975
rect 43258 527640 43314 527649
rect 43258 527575 43314 527584
rect 43272 498817 43300 527575
rect 43258 498808 43314 498817
rect 43258 498743 43314 498752
rect 43352 497480 43404 497486
rect 43352 497422 43404 497428
rect 43258 496768 43314 496777
rect 43258 496703 43314 496712
rect 43166 496088 43222 496097
rect 43166 496023 43222 496032
rect 43074 353288 43130 353297
rect 43074 353223 43130 353232
rect 43272 351218 43300 496703
rect 43364 420238 43392 497422
rect 43456 493377 43484 558039
rect 43916 552537 43944 582111
rect 43902 552528 43958 552537
rect 43902 552463 43958 552472
rect 43904 522572 43956 522578
rect 43904 522514 43956 522520
rect 43812 522300 43864 522306
rect 43812 522242 43864 522248
rect 43824 521937 43852 522242
rect 43810 521928 43866 521937
rect 43810 521863 43866 521872
rect 43812 521756 43864 521762
rect 43812 521698 43864 521704
rect 43628 521280 43680 521286
rect 43628 521222 43680 521228
rect 43536 520328 43588 520334
rect 43536 520270 43588 520276
rect 43442 493368 43498 493377
rect 43442 493303 43498 493312
rect 43352 420232 43404 420238
rect 43352 420174 43404 420180
rect 43548 366450 43576 520270
rect 43536 366444 43588 366450
rect 43536 366386 43588 366392
rect 43640 365022 43668 521222
rect 43720 519648 43772 519654
rect 43720 519590 43772 519596
rect 43628 365016 43680 365022
rect 43628 364958 43680 364964
rect 43732 363798 43760 519590
rect 43720 363792 43772 363798
rect 43720 363734 43772 363740
rect 43260 351212 43312 351218
rect 43260 351154 43312 351160
rect 42616 350124 42668 350130
rect 42616 350066 42668 350072
rect 43824 350062 43852 521698
rect 43812 350056 43864 350062
rect 43812 349998 43864 350004
rect 43916 349926 43944 522514
rect 44008 472025 44036 647527
rect 45006 639024 45062 639033
rect 45006 638959 45062 638968
rect 44914 578912 44970 578921
rect 44914 578847 44970 578856
rect 44822 576736 44878 576745
rect 44822 576671 44878 576680
rect 44836 555801 44864 576671
rect 44822 555792 44878 555801
rect 44822 555727 44878 555736
rect 44928 555529 44956 578847
rect 44914 555520 44970 555529
rect 44914 555455 44970 555464
rect 44638 549808 44694 549817
rect 44638 549743 44694 549752
rect 44178 527504 44234 527513
rect 44178 527439 44234 527448
rect 44192 525201 44220 527439
rect 44178 525192 44234 525201
rect 44178 525127 44234 525136
rect 44180 524544 44232 524550
rect 44180 524486 44232 524492
rect 44192 523734 44220 524486
rect 44180 523728 44232 523734
rect 44180 523670 44232 523676
rect 44088 522232 44140 522238
rect 44088 522174 44140 522180
rect 44100 521801 44128 522174
rect 44086 521792 44142 521801
rect 44086 521727 44142 521736
rect 44652 510105 44680 549743
rect 44730 538248 44786 538257
rect 44730 538183 44786 538192
rect 44638 510096 44694 510105
rect 44638 510031 44694 510040
rect 44744 500857 44772 538183
rect 44914 533624 44970 533633
rect 44914 533559 44970 533568
rect 44822 528728 44878 528737
rect 44822 528663 44878 528672
rect 44730 500848 44786 500857
rect 44730 500783 44786 500792
rect 44836 475561 44864 528663
rect 44822 475552 44878 475561
rect 44822 475487 44878 475496
rect 44928 472705 44956 533559
rect 45020 494057 45048 638959
rect 45284 592068 45336 592074
rect 45284 592010 45336 592016
rect 45098 591968 45154 591977
rect 45098 591903 45154 591912
rect 45112 560153 45140 591903
rect 45190 589792 45246 589801
rect 45190 589727 45246 589736
rect 45098 560144 45154 560153
rect 45098 560079 45154 560088
rect 45204 557433 45232 589727
rect 45296 560250 45324 592010
rect 45374 590880 45430 590889
rect 45374 590815 45430 590824
rect 45284 560244 45336 560250
rect 45284 560186 45336 560192
rect 45388 558657 45416 590815
rect 45374 558648 45430 558657
rect 45374 558583 45430 558592
rect 45190 557424 45246 557433
rect 45190 557359 45246 557368
rect 45284 522164 45336 522170
rect 45284 522106 45336 522112
rect 45100 522096 45152 522102
rect 45100 522038 45152 522044
rect 45006 494048 45062 494057
rect 45006 493983 45062 493992
rect 44914 472696 44970 472705
rect 44914 472631 44970 472640
rect 43994 472016 44050 472025
rect 43994 471951 44050 471960
rect 45112 363662 45140 522038
rect 45192 521688 45244 521694
rect 45192 521630 45244 521636
rect 45100 363656 45152 363662
rect 45100 363598 45152 363604
rect 45204 362234 45232 521630
rect 45192 362228 45244 362234
rect 45192 362170 45244 362176
rect 45296 360874 45324 522106
rect 45376 520804 45428 520810
rect 45376 520746 45428 520752
rect 45284 360868 45336 360874
rect 45284 360810 45336 360816
rect 45388 356726 45416 520746
rect 45480 387462 45508 658242
rect 58624 657348 58676 657354
rect 58624 657290 58676 657296
rect 53562 649632 53618 649641
rect 53562 649567 53618 649576
rect 51446 649360 51502 649369
rect 51446 649295 51502 649304
rect 46846 644056 46902 644065
rect 46846 643991 46902 644000
rect 46754 594144 46810 594153
rect 46754 594079 46810 594088
rect 46662 580000 46718 580009
rect 46662 579935 46718 579944
rect 46570 577824 46626 577833
rect 46570 577759 46626 577768
rect 46584 557025 46612 577759
rect 46570 557016 46626 557025
rect 46570 556951 46626 556960
rect 46676 555257 46704 579935
rect 46768 559881 46796 594079
rect 46754 559872 46810 559881
rect 46754 559807 46810 559816
rect 46662 555248 46718 555257
rect 46662 555183 46718 555192
rect 46570 551304 46626 551313
rect 46570 551239 46626 551248
rect 46386 545456 46442 545465
rect 46386 545391 46442 545400
rect 46294 534304 46350 534313
rect 46294 534239 46350 534248
rect 46110 522608 46166 522617
rect 46110 522543 46166 522552
rect 46018 519480 46074 519489
rect 46018 519415 46074 519424
rect 45468 387456 45520 387462
rect 45468 387398 45520 387404
rect 46032 363633 46060 519415
rect 46124 508473 46152 522543
rect 46202 520840 46258 520849
rect 46202 520775 46258 520784
rect 46110 508464 46166 508473
rect 46110 508399 46166 508408
rect 46216 498953 46244 520775
rect 46202 498944 46258 498953
rect 46202 498879 46258 498888
rect 46204 420232 46256 420238
rect 46204 420174 46256 420180
rect 46216 389910 46244 420174
rect 46308 418169 46336 534239
rect 46400 418713 46428 545391
rect 46478 520432 46534 520441
rect 46478 520367 46534 520376
rect 46492 496233 46520 520367
rect 46584 516633 46612 551239
rect 46756 527196 46808 527202
rect 46756 527138 46808 527144
rect 46664 526176 46716 526182
rect 46664 526118 46716 526124
rect 46570 516624 46626 516633
rect 46570 516559 46626 516568
rect 46478 496224 46534 496233
rect 46478 496159 46534 496168
rect 46480 493332 46532 493338
rect 46480 493274 46532 493280
rect 46386 418704 46442 418713
rect 46386 418639 46442 418648
rect 46294 418160 46350 418169
rect 46294 418095 46350 418104
rect 46204 389904 46256 389910
rect 46204 389846 46256 389852
rect 46018 363624 46074 363633
rect 46018 363559 46074 363568
rect 45376 356720 45428 356726
rect 45376 356662 45428 356668
rect 46492 352782 46520 493274
rect 46676 364206 46704 526118
rect 46664 364200 46716 364206
rect 46664 364142 46716 364148
rect 46480 352776 46532 352782
rect 46480 352718 46532 352724
rect 46768 352714 46796 527138
rect 46860 394777 46888 643991
rect 49606 643784 49662 643793
rect 49606 643719 49662 643728
rect 48042 643512 48098 643521
rect 48042 643447 48098 643456
rect 47950 581088 48006 581097
rect 47950 581023 48006 581032
rect 47858 575648 47914 575657
rect 47858 575583 47914 575592
rect 47872 556073 47900 575583
rect 47964 556753 47992 581023
rect 47950 556744 48006 556753
rect 47950 556679 48006 556688
rect 47858 556064 47914 556073
rect 47858 555999 47914 556008
rect 47766 548176 47822 548185
rect 47766 548111 47822 548120
rect 47674 545592 47730 545601
rect 47674 545527 47730 545536
rect 47582 522064 47638 522073
rect 47582 521999 47638 522008
rect 47490 521112 47546 521121
rect 47490 521047 47546 521056
rect 47398 519208 47454 519217
rect 47398 519143 47454 519152
rect 47412 508609 47440 519143
rect 47398 508600 47454 508609
rect 47398 508535 47454 508544
rect 47398 506560 47454 506569
rect 47398 506495 47454 506504
rect 46846 394768 46902 394777
rect 46846 394703 46902 394712
rect 47412 364002 47440 506495
rect 47504 499769 47532 521047
rect 47490 499760 47546 499769
rect 47490 499695 47546 499704
rect 47596 496369 47624 521999
rect 47582 496360 47638 496369
rect 47582 496295 47638 496304
rect 47688 425785 47716 545527
rect 47674 425776 47730 425785
rect 47674 425711 47730 425720
rect 47780 424697 47808 548111
rect 47952 526244 48004 526250
rect 47952 526186 48004 526192
rect 47858 521928 47914 521937
rect 47858 521863 47914 521872
rect 47872 505889 47900 521863
rect 47858 505880 47914 505889
rect 47858 505815 47914 505824
rect 47766 424688 47822 424697
rect 47766 424623 47822 424632
rect 47400 363996 47452 364002
rect 47400 363938 47452 363944
rect 46756 352708 46808 352714
rect 46756 352650 46808 352656
rect 43904 349920 43956 349926
rect 43904 349862 43956 349868
rect 41144 349852 41196 349858
rect 41144 349794 41196 349800
rect 47964 347138 47992 526186
rect 48056 458969 48084 643447
rect 48226 642696 48282 642705
rect 48226 642631 48282 642640
rect 48134 640928 48190 640937
rect 48134 640863 48190 640872
rect 48042 458960 48098 458969
rect 48042 458895 48098 458904
rect 48148 456793 48176 640863
rect 48240 457337 48268 642631
rect 49514 595232 49570 595241
rect 49514 595167 49570 595176
rect 49422 587616 49478 587625
rect 49422 587551 49478 587560
rect 49330 586392 49386 586401
rect 49330 586327 49386 586336
rect 49238 585440 49294 585449
rect 49238 585375 49294 585384
rect 49252 557297 49280 585375
rect 49238 557288 49294 557297
rect 49238 557223 49294 557232
rect 49344 557161 49372 586327
rect 49330 557152 49386 557161
rect 49330 557087 49386 557096
rect 49436 555665 49464 587551
rect 49528 560561 49556 595167
rect 49514 560552 49570 560561
rect 49514 560487 49570 560496
rect 49422 555656 49478 555665
rect 49422 555591 49478 555600
rect 49422 552120 49478 552129
rect 49422 552055 49478 552064
rect 49330 544640 49386 544649
rect 49330 544575 49386 544584
rect 49238 541512 49294 541521
rect 49238 541447 49294 541456
rect 49146 538792 49202 538801
rect 49146 538727 49202 538736
rect 49054 537160 49110 537169
rect 49054 537095 49110 537104
rect 48962 535936 49018 535945
rect 48962 535871 49018 535880
rect 48870 521792 48926 521801
rect 48870 521727 48926 521736
rect 48780 521144 48832 521150
rect 48780 521086 48832 521092
rect 48226 457328 48282 457337
rect 48226 457263 48282 457272
rect 48134 456784 48190 456793
rect 48134 456719 48190 456728
rect 48792 349994 48820 521086
rect 48884 506841 48912 521727
rect 48870 506832 48926 506841
rect 48870 506767 48926 506776
rect 48976 436665 49004 535871
rect 49068 438297 49096 537095
rect 49054 438288 49110 438297
rect 49054 438223 49110 438232
rect 49160 437209 49188 538727
rect 49146 437200 49202 437209
rect 49146 437135 49202 437144
rect 48962 436656 49018 436665
rect 48962 436591 49018 436600
rect 49252 432857 49280 541447
rect 49344 433401 49372 544575
rect 49436 436121 49464 552055
rect 49516 518968 49568 518974
rect 49516 518910 49568 518916
rect 49528 507890 49556 518910
rect 49516 507884 49568 507890
rect 49516 507826 49568 507832
rect 49620 459513 49648 643719
rect 50618 641880 50674 641889
rect 50618 641815 50674 641824
rect 50066 639976 50122 639985
rect 50066 639911 50122 639920
rect 50080 463321 50108 639911
rect 50526 550080 50582 550089
rect 50526 550015 50582 550024
rect 50434 546952 50490 546961
rect 50434 546887 50490 546896
rect 50342 545184 50398 545193
rect 50342 545119 50398 545128
rect 50250 540016 50306 540025
rect 50250 539951 50306 539960
rect 50158 523152 50214 523161
rect 50158 523087 50214 523096
rect 50066 463312 50122 463321
rect 50066 463247 50122 463256
rect 49606 459504 49662 459513
rect 49606 459439 49662 459448
rect 49422 436112 49478 436121
rect 49422 436047 49478 436056
rect 49330 433392 49386 433401
rect 49330 433327 49386 433336
rect 49238 432848 49294 432857
rect 49238 432783 49294 432792
rect 50172 426329 50200 523087
rect 50264 435577 50292 539951
rect 50250 435568 50306 435577
rect 50250 435503 50306 435512
rect 50356 430681 50384 545119
rect 50342 430672 50398 430681
rect 50342 430607 50398 430616
rect 50158 426320 50214 426329
rect 50158 426255 50214 426264
rect 50448 424153 50476 546887
rect 50434 424144 50490 424153
rect 50434 424079 50490 424088
rect 50540 422521 50568 550015
rect 50632 483041 50660 641815
rect 50710 637800 50766 637809
rect 50710 637735 50766 637744
rect 50618 483032 50674 483041
rect 50618 482967 50674 482976
rect 50618 482896 50674 482905
rect 50618 482831 50674 482840
rect 50526 422512 50582 422521
rect 50526 422447 50582 422456
rect 48780 349988 48832 349994
rect 48780 349930 48832 349936
rect 50632 347206 50660 482831
rect 50724 464409 50752 637735
rect 50894 637528 50950 637537
rect 50894 637463 50950 637472
rect 50804 523592 50856 523598
rect 50804 523534 50856 523540
rect 50710 464400 50766 464409
rect 50710 464335 50766 464344
rect 50816 350266 50844 523534
rect 50908 462233 50936 637463
rect 51460 528554 51488 649295
rect 52274 649224 52330 649233
rect 52274 649159 52330 649168
rect 51814 648136 51870 648145
rect 51814 648071 51870 648080
rect 51630 533352 51686 533361
rect 51630 533287 51686 533296
rect 51276 528526 51488 528554
rect 50988 527332 51040 527338
rect 50988 527274 51040 527280
rect 51000 527241 51028 527274
rect 50986 527232 51042 527241
rect 50986 527167 51042 527176
rect 50988 521620 51040 521626
rect 50988 521562 51040 521568
rect 51000 520305 51028 521562
rect 50986 520296 51042 520305
rect 50986 520231 51042 520240
rect 51276 520010 51304 528526
rect 51538 526688 51594 526697
rect 51460 526646 51538 526674
rect 51460 520146 51488 526646
rect 51538 526623 51594 526632
rect 51540 521416 51592 521422
rect 51540 521358 51592 521364
rect 51552 520305 51580 521358
rect 51538 520296 51594 520305
rect 51538 520231 51594 520240
rect 51460 520118 51580 520146
rect 51276 519982 51488 520010
rect 51080 467152 51132 467158
rect 51080 467094 51132 467100
rect 51092 462330 51120 467094
rect 51460 465497 51488 519982
rect 51446 465488 51502 465497
rect 51446 465423 51502 465432
rect 51080 462324 51132 462330
rect 51080 462266 51132 462272
rect 50894 462224 50950 462233
rect 50894 462159 50950 462168
rect 51552 433945 51580 520118
rect 51644 434489 51672 533287
rect 51722 529000 51778 529009
rect 51722 528935 51778 528944
rect 51630 434480 51686 434489
rect 51630 434415 51686 434424
rect 51538 433936 51594 433945
rect 51538 433871 51594 433880
rect 51736 417625 51764 528935
rect 51828 482361 51856 648071
rect 52182 647728 52238 647737
rect 52182 647663 52238 647672
rect 52090 647456 52146 647465
rect 52090 647391 52146 647400
rect 51906 642968 51962 642977
rect 51906 642903 51962 642912
rect 51814 482352 51870 482361
rect 51814 482287 51870 482296
rect 51816 478168 51868 478174
rect 51816 478110 51868 478116
rect 51722 417616 51778 417625
rect 51722 417551 51778 417560
rect 51080 392624 51132 392630
rect 51080 392566 51132 392572
rect 51092 389842 51120 392566
rect 51828 389978 51856 478110
rect 51920 476377 51948 642903
rect 51998 641472 52054 641481
rect 51998 641407 52054 641416
rect 51906 476368 51962 476377
rect 51906 476303 51962 476312
rect 51906 475552 51962 475561
rect 51906 475487 51962 475496
rect 51920 407289 51948 475487
rect 52012 472569 52040 641407
rect 52104 476921 52132 647391
rect 52090 476912 52146 476921
rect 52090 476847 52146 476856
rect 52196 474745 52224 647663
rect 52182 474736 52238 474745
rect 52182 474671 52238 474680
rect 52288 474201 52316 649159
rect 53010 646776 53066 646785
rect 53010 646711 53066 646720
rect 52918 639568 52974 639577
rect 52918 639503 52974 639512
rect 52552 523048 52604 523054
rect 52552 522990 52604 522996
rect 52460 522368 52512 522374
rect 52460 522310 52512 522316
rect 52472 520946 52500 522310
rect 52460 520940 52512 520946
rect 52460 520882 52512 520888
rect 52368 520532 52420 520538
rect 52368 520474 52420 520480
rect 52380 520305 52408 520474
rect 52366 520296 52422 520305
rect 52366 520231 52422 520240
rect 52368 519716 52420 519722
rect 52368 519658 52420 519664
rect 52380 519353 52408 519658
rect 52564 519654 52592 522990
rect 52828 522436 52880 522442
rect 52828 522378 52880 522384
rect 52736 520124 52788 520130
rect 52736 520066 52788 520072
rect 52552 519648 52604 519654
rect 52552 519590 52604 519596
rect 52366 519344 52422 519353
rect 52366 519279 52422 519288
rect 52366 476232 52422 476241
rect 52366 476167 52422 476176
rect 52274 474192 52330 474201
rect 52274 474127 52330 474136
rect 52182 472696 52238 472705
rect 52182 472631 52238 472640
rect 51998 472560 52054 472569
rect 51998 472495 52054 472504
rect 52196 407833 52224 472631
rect 52182 407824 52238 407833
rect 52182 407759 52238 407768
rect 51906 407280 51962 407289
rect 51906 407215 51962 407224
rect 51816 389972 51868 389978
rect 51816 389914 51868 389920
rect 51080 389836 51132 389842
rect 51080 389778 51132 389784
rect 52380 352986 52408 476167
rect 52748 353054 52776 520066
rect 52840 503130 52868 522378
rect 52828 503124 52880 503130
rect 52828 503066 52880 503072
rect 52932 463865 52960 639503
rect 53024 470393 53052 646711
rect 53378 640384 53434 640393
rect 53378 640319 53434 640328
rect 53196 525088 53248 525094
rect 53196 525030 53248 525036
rect 53102 503704 53158 503713
rect 53102 503639 53158 503648
rect 53010 470384 53066 470393
rect 53010 470319 53066 470328
rect 52918 463856 52974 463865
rect 52918 463791 52974 463800
rect 53116 355502 53144 503639
rect 53208 425241 53236 525030
rect 53288 520192 53340 520198
rect 53288 520134 53340 520140
rect 53300 514078 53328 520134
rect 53288 514072 53340 514078
rect 53288 514014 53340 514020
rect 53288 511284 53340 511290
rect 53288 511226 53340 511232
rect 53194 425232 53250 425241
rect 53194 425167 53250 425176
rect 53300 358086 53328 511226
rect 53392 475289 53420 640319
rect 53470 574560 53526 574569
rect 53470 574495 53526 574504
rect 53484 556889 53512 574495
rect 53470 556880 53526 556889
rect 53470 556815 53526 556824
rect 53472 527264 53524 527270
rect 53472 527206 53524 527212
rect 53484 514826 53512 527206
rect 53472 514820 53524 514826
rect 53472 514762 53524 514768
rect 53576 478553 53604 649567
rect 54850 649088 54906 649097
rect 54850 649023 54906 649032
rect 54114 648000 54170 648009
rect 54114 647935 54170 647944
rect 53840 558884 53892 558890
rect 53840 558826 53892 558832
rect 53852 558113 53880 558826
rect 53932 558816 53984 558822
rect 53932 558758 53984 558764
rect 53838 558104 53894 558113
rect 53838 558039 53894 558048
rect 53944 557977 53972 558758
rect 53930 557968 53986 557977
rect 53930 557903 53986 557912
rect 53840 557524 53892 557530
rect 53840 557466 53892 557472
rect 53852 556209 53880 557466
rect 53838 556200 53894 556209
rect 53838 556135 53894 556144
rect 53840 555960 53892 555966
rect 53840 555902 53892 555908
rect 53852 554985 53880 555902
rect 53838 554976 53894 554985
rect 53838 554911 53894 554920
rect 53748 529984 53800 529990
rect 53748 529926 53800 529932
rect 53760 529825 53788 529926
rect 53746 529816 53802 529825
rect 53746 529751 53802 529760
rect 53840 524204 53892 524210
rect 53840 524146 53892 524152
rect 53852 523161 53880 524146
rect 53838 523152 53894 523161
rect 53838 523087 53894 523096
rect 53748 521008 53800 521014
rect 53748 520950 53800 520956
rect 53760 518894 53788 520950
rect 53668 518866 53788 518894
rect 53668 514758 53696 518866
rect 53748 514888 53800 514894
rect 53748 514830 53800 514836
rect 53656 514752 53708 514758
rect 53656 514694 53708 514700
rect 53656 514072 53708 514078
rect 53656 514014 53708 514020
rect 53668 501634 53696 514014
rect 53760 509930 53788 514830
rect 53748 509924 53800 509930
rect 53748 509866 53800 509872
rect 53656 501628 53708 501634
rect 53656 501570 53708 501576
rect 53562 478544 53618 478553
rect 53562 478479 53618 478488
rect 53378 475280 53434 475289
rect 53378 475215 53434 475224
rect 54128 470937 54156 647935
rect 54392 647284 54444 647290
rect 54392 647226 54444 647232
rect 54404 644474 54432 647226
rect 54312 644446 54432 644474
rect 54114 470928 54170 470937
rect 54114 470863 54170 470872
rect 54312 460057 54340 644446
rect 54758 641744 54814 641753
rect 54758 641679 54814 641688
rect 54666 635488 54722 635497
rect 54666 635423 54722 635432
rect 54574 634672 54630 634681
rect 54574 634607 54630 634616
rect 54588 599593 54616 634607
rect 54574 599584 54630 599593
rect 54574 599519 54630 599528
rect 54680 597417 54708 635423
rect 54666 597408 54722 597417
rect 54666 597343 54722 597352
rect 54666 588704 54722 588713
rect 54666 588639 54722 588648
rect 54574 584352 54630 584361
rect 54574 584287 54630 584296
rect 54482 572384 54538 572393
rect 54482 572319 54538 572328
rect 54496 558793 54524 572319
rect 54482 558784 54538 558793
rect 54482 558719 54538 558728
rect 54588 558521 54616 584287
rect 54574 558512 54630 558521
rect 54574 558447 54630 558456
rect 54680 556617 54708 588639
rect 54666 556608 54722 556617
rect 54666 556543 54722 556552
rect 54666 544232 54722 544241
rect 54666 544167 54722 544176
rect 54390 538384 54446 538393
rect 54390 538319 54446 538328
rect 54298 460048 54354 460057
rect 54298 459983 54354 459992
rect 54404 412729 54432 538319
rect 54576 524476 54628 524482
rect 54576 524418 54628 524424
rect 54588 514894 54616 524418
rect 54576 514888 54628 514894
rect 54576 514830 54628 514836
rect 54484 514820 54536 514826
rect 54484 514762 54536 514768
rect 54390 412720 54446 412729
rect 54390 412655 54446 412664
rect 53288 358080 53340 358086
rect 53288 358022 53340 358028
rect 53104 355496 53156 355502
rect 53104 355438 53156 355444
rect 52736 353048 52788 353054
rect 52736 352990 52788 352996
rect 52368 352980 52420 352986
rect 52368 352922 52420 352928
rect 54496 352850 54524 514762
rect 54574 513360 54630 513369
rect 54574 513295 54630 513304
rect 54588 358154 54616 513295
rect 54680 411641 54708 544167
rect 54772 481817 54800 641679
rect 54758 481808 54814 481817
rect 54758 481743 54814 481752
rect 54864 478009 54892 649023
rect 56230 648816 56286 648825
rect 56230 648751 56286 648760
rect 55586 640792 55642 640801
rect 55586 640727 55642 640736
rect 54942 640656 54998 640665
rect 54942 640591 54998 640600
rect 54850 478000 54906 478009
rect 54850 477935 54906 477944
rect 54956 466041 54984 640591
rect 55126 583264 55182 583273
rect 55126 583199 55182 583208
rect 55034 573472 55090 573481
rect 55034 573407 55090 573416
rect 55048 555393 55076 573407
rect 55140 559337 55168 583199
rect 55126 559328 55182 559337
rect 55126 559263 55182 559272
rect 55034 555384 55090 555393
rect 55034 555319 55090 555328
rect 55128 528420 55180 528426
rect 55128 528362 55180 528368
rect 55140 527241 55168 528362
rect 55126 527232 55182 527241
rect 55126 527167 55182 527176
rect 55034 520160 55090 520169
rect 55034 520095 55090 520104
rect 55048 510678 55076 520095
rect 55036 510672 55088 510678
rect 55036 510614 55088 510620
rect 55128 503668 55180 503674
rect 55128 503610 55180 503616
rect 55140 499594 55168 503610
rect 55128 499588 55180 499594
rect 55128 499530 55180 499536
rect 55600 466585 55628 640727
rect 56046 635624 56102 635633
rect 56046 635559 56102 635568
rect 56060 596329 56088 635559
rect 56138 612640 56194 612649
rect 56138 612575 56194 612584
rect 56046 596320 56102 596329
rect 56046 596255 56102 596264
rect 55954 570208 56010 570217
rect 55954 570143 56010 570152
rect 55770 566808 55826 566817
rect 55770 566743 55826 566752
rect 55784 552945 55812 566743
rect 55968 557954 55996 570143
rect 56048 558748 56100 558754
rect 56048 558690 56100 558696
rect 56060 558249 56088 558690
rect 56046 558240 56102 558249
rect 56046 558175 56102 558184
rect 56046 557968 56102 557977
rect 55968 557926 56046 557954
rect 56046 557903 56102 557912
rect 56048 556232 56100 556238
rect 56048 556174 56100 556180
rect 55770 552936 55826 552945
rect 55770 552871 55826 552880
rect 56060 552809 56088 556174
rect 56046 552800 56102 552809
rect 56046 552735 56102 552744
rect 56046 546680 56102 546689
rect 56046 546615 56102 546624
rect 55678 542736 55734 542745
rect 55678 542671 55734 542680
rect 55586 466576 55642 466585
rect 55586 466511 55642 466520
rect 54942 466032 54998 466041
rect 54942 465967 54998 465976
rect 54760 462324 54812 462330
rect 54760 462266 54812 462272
rect 54666 411632 54722 411641
rect 54666 411567 54722 411576
rect 54772 400926 54800 462266
rect 55692 431225 55720 542671
rect 55954 542600 56010 542609
rect 55954 542535 56010 542544
rect 55770 541376 55826 541385
rect 55770 541311 55826 541320
rect 55678 431216 55734 431225
rect 55678 431151 55734 431160
rect 55784 411097 55812 541311
rect 55864 523456 55916 523462
rect 55864 523398 55916 523404
rect 55876 518974 55904 523398
rect 55864 518968 55916 518974
rect 55864 518910 55916 518916
rect 55864 514752 55916 514758
rect 55864 514694 55916 514700
rect 55876 505170 55904 514694
rect 55864 505164 55916 505170
rect 55864 505106 55916 505112
rect 55862 499896 55918 499905
rect 55862 499831 55918 499840
rect 55770 411088 55826 411097
rect 55770 411023 55826 411032
rect 54760 400920 54812 400926
rect 54760 400862 54812 400868
rect 54576 358148 54628 358154
rect 54576 358090 54628 358096
rect 54484 352844 54536 352850
rect 54484 352786 54536 352792
rect 50804 350260 50856 350266
rect 50804 350202 50856 350208
rect 55876 350198 55904 499831
rect 55968 409465 55996 542535
rect 55954 409456 56010 409465
rect 55954 409391 56010 409400
rect 56060 406745 56088 546615
rect 56152 545873 56180 612575
rect 56138 545864 56194 545873
rect 56138 545799 56194 545808
rect 56140 520260 56192 520266
rect 56140 520202 56192 520208
rect 56046 406736 56102 406745
rect 56046 406671 56102 406680
rect 56152 352918 56180 520202
rect 56244 479641 56272 648751
rect 56414 647864 56470 647873
rect 56414 647799 56470 647808
rect 56322 641064 56378 641073
rect 56322 640999 56378 641008
rect 56230 479632 56286 479641
rect 56230 479567 56286 479576
rect 56230 478952 56286 478961
rect 56230 478887 56286 478896
rect 56244 358222 56272 478887
rect 56336 468761 56364 640999
rect 56428 473657 56456 647799
rect 57886 642832 57942 642841
rect 57808 642790 57886 642818
rect 56506 640520 56562 640529
rect 56506 640455 56508 640464
rect 56560 640455 56562 640464
rect 56508 640426 56560 640432
rect 57702 635760 57758 635769
rect 57702 635695 57758 635704
rect 57610 624608 57666 624617
rect 57610 624543 57666 624552
rect 56966 622432 57022 622441
rect 56966 622367 57022 622376
rect 56506 568032 56562 568041
rect 56506 567967 56562 567976
rect 56520 556238 56548 567967
rect 56980 559162 57008 622367
rect 57242 621344 57298 621353
rect 57242 621279 57298 621288
rect 57058 605024 57114 605033
rect 57058 604959 57114 604968
rect 56968 559156 57020 559162
rect 56968 559098 57020 559104
rect 56508 556232 56560 556238
rect 56508 556174 56560 556180
rect 56508 556096 56560 556102
rect 56508 556038 56560 556044
rect 56520 554849 56548 556038
rect 56506 554840 56562 554849
rect 56506 554775 56562 554784
rect 56508 553308 56560 553314
rect 56508 553250 56560 553256
rect 56520 552129 56548 553250
rect 56506 552120 56562 552129
rect 56506 552055 56562 552064
rect 56508 546440 56560 546446
rect 56508 546382 56560 546388
rect 56520 545193 56548 546382
rect 56506 545184 56562 545193
rect 56506 545119 56562 545128
rect 57072 536217 57100 604959
rect 57150 562456 57206 562465
rect 57150 562391 57206 562400
rect 57164 543017 57192 562391
rect 57256 559230 57284 621279
rect 57334 611552 57390 611561
rect 57334 611487 57390 611496
rect 57244 559224 57296 559230
rect 57244 559166 57296 559172
rect 57348 557534 57376 611487
rect 57426 609376 57482 609385
rect 57426 609311 57482 609320
rect 57256 557506 57376 557534
rect 57256 549953 57284 557506
rect 57336 554736 57388 554742
rect 57336 554678 57388 554684
rect 57242 549944 57298 549953
rect 57242 549879 57298 549888
rect 57348 547874 57376 554678
rect 57256 547846 57376 547874
rect 57150 543008 57206 543017
rect 57150 542943 57206 542952
rect 57058 536208 57114 536217
rect 57058 536143 57114 536152
rect 56966 532400 57022 532409
rect 56966 532335 57022 532344
rect 56508 520056 56560 520062
rect 56508 519998 56560 520004
rect 56520 514049 56548 519998
rect 56506 514040 56562 514049
rect 56506 513975 56562 513984
rect 56980 511737 57008 532335
rect 57150 532264 57206 532273
rect 57150 532199 57206 532208
rect 57058 526416 57114 526425
rect 57058 526351 57114 526360
rect 57072 512825 57100 526351
rect 57058 512816 57114 512825
rect 57058 512751 57114 512760
rect 56966 511728 57022 511737
rect 56966 511663 57022 511672
rect 57164 511193 57192 532199
rect 57256 513369 57284 547846
rect 57440 547097 57468 609311
rect 57518 593056 57574 593065
rect 57518 592991 57574 593000
rect 57532 592074 57560 592991
rect 57520 592068 57572 592074
rect 57520 592010 57572 592016
rect 57624 567194 57652 624543
rect 57716 600681 57744 635695
rect 57808 631145 57836 642790
rect 57886 642767 57942 642776
rect 57886 641880 57942 641889
rect 57886 641815 57942 641824
rect 57900 641782 57928 641815
rect 57888 641776 57940 641782
rect 57888 641718 57940 641724
rect 58530 637392 58586 637401
rect 58530 637327 58586 637336
rect 58346 634808 58402 634817
rect 58346 634743 58402 634752
rect 57794 631136 57850 631145
rect 57794 631071 57850 631080
rect 57886 625696 57942 625705
rect 57886 625631 57942 625640
rect 57794 623520 57850 623529
rect 57794 623455 57850 623464
rect 57702 600672 57758 600681
rect 57702 600607 57758 600616
rect 57532 567166 57652 567194
rect 57532 559094 57560 567166
rect 57702 563544 57758 563553
rect 57702 563479 57758 563488
rect 57610 560280 57666 560289
rect 57610 560215 57666 560224
rect 57520 559088 57572 559094
rect 57520 559030 57572 559036
rect 57624 557054 57652 560215
rect 57612 557048 57664 557054
rect 57612 556990 57664 556996
rect 57612 554056 57664 554062
rect 57612 553998 57664 554004
rect 57426 547088 57482 547097
rect 57426 547023 57482 547032
rect 57518 532128 57574 532137
rect 57336 532092 57388 532098
rect 57518 532063 57574 532072
rect 57336 532034 57388 532040
rect 57348 517177 57376 532034
rect 57428 532024 57480 532030
rect 57428 531966 57480 531972
rect 57334 517168 57390 517177
rect 57334 517103 57390 517112
rect 57440 515545 57468 531966
rect 57426 515536 57482 515545
rect 57426 515471 57482 515480
rect 57242 513360 57298 513369
rect 57242 513295 57298 513304
rect 57532 512281 57560 532063
rect 57624 516089 57652 553998
rect 57716 544513 57744 563479
rect 57808 550633 57836 623455
rect 57794 550624 57850 550633
rect 57794 550559 57850 550568
rect 57702 544504 57758 544513
rect 57702 544439 57758 544448
rect 57900 539481 57928 625631
rect 58254 615904 58310 615913
rect 58254 615839 58310 615848
rect 58070 603936 58126 603945
rect 58070 603871 58126 603880
rect 58084 540433 58112 603871
rect 58268 547369 58296 615839
rect 58360 598505 58388 634743
rect 58438 614816 58494 614825
rect 58438 614751 58494 614760
rect 58346 598496 58402 598505
rect 58346 598431 58402 598440
rect 58346 564632 58402 564641
rect 58346 564567 58402 564576
rect 58360 553353 58388 564567
rect 58346 553344 58402 553353
rect 58346 553279 58402 553288
rect 58254 547360 58310 547369
rect 58254 547295 58310 547304
rect 58070 540424 58126 540433
rect 58070 540359 58126 540368
rect 57886 539472 57942 539481
rect 57886 539407 57942 539416
rect 57794 531584 57850 531593
rect 57794 531519 57850 531528
rect 57704 524408 57756 524414
rect 57704 524350 57756 524356
rect 57716 523161 57744 524350
rect 57702 523152 57758 523161
rect 57702 523087 57758 523096
rect 57704 516180 57756 516186
rect 57704 516122 57756 516128
rect 57610 516080 57666 516089
rect 57610 516015 57666 516024
rect 57518 512272 57574 512281
rect 57518 512207 57574 512216
rect 57150 511184 57206 511193
rect 57150 511119 57206 511128
rect 56600 510672 56652 510678
rect 56600 510614 56652 510620
rect 57518 510640 57574 510649
rect 56612 503674 56640 510614
rect 57518 510575 57574 510584
rect 57152 507884 57204 507890
rect 57152 507826 57204 507832
rect 56600 503668 56652 503674
rect 56600 503610 56652 503616
rect 57058 496088 57114 496097
rect 57058 496023 57114 496032
rect 57072 489977 57100 496023
rect 57164 494766 57192 507826
rect 57426 503704 57482 503713
rect 57426 503639 57482 503648
rect 57334 500712 57390 500721
rect 57334 500647 57390 500656
rect 57244 499588 57296 499594
rect 57244 499530 57296 499536
rect 57152 494760 57204 494766
rect 57152 494702 57204 494708
rect 57150 493368 57206 493377
rect 57150 493303 57206 493312
rect 57164 491638 57192 493303
rect 57152 491632 57204 491638
rect 57152 491574 57204 491580
rect 57150 491192 57206 491201
rect 57150 491127 57206 491136
rect 57058 489968 57114 489977
rect 57058 489903 57114 489912
rect 56414 473648 56470 473657
rect 56414 473583 56470 473592
rect 56322 468752 56378 468761
rect 56322 468687 56378 468696
rect 57164 428505 57192 491127
rect 57150 428496 57206 428505
rect 57150 428431 57206 428440
rect 56232 358216 56284 358222
rect 56232 358158 56284 358164
rect 57256 355638 57284 499530
rect 57348 358290 57376 500647
rect 57440 366654 57468 503639
rect 57532 498930 57560 510575
rect 57610 505880 57666 505889
rect 57610 505815 57666 505824
rect 57624 499050 57652 505815
rect 57716 500954 57744 516122
rect 57808 515001 57836 531519
rect 57886 531448 57942 531457
rect 57886 531383 57942 531392
rect 57794 514992 57850 515001
rect 57794 514927 57850 514936
rect 57900 513913 57928 531383
rect 58452 529825 58480 614751
rect 58544 601769 58572 637327
rect 58636 632058 58664 657290
rect 66534 646912 66590 646921
rect 66534 646847 66590 646856
rect 62670 645280 62726 645289
rect 62670 645215 62726 645224
rect 59266 642424 59322 642433
rect 59266 642359 59322 642368
rect 59082 642288 59138 642297
rect 59082 642223 59138 642232
rect 59096 633321 59124 642223
rect 59280 641986 59308 642359
rect 59268 641980 59320 641986
rect 59268 641922 59320 641928
rect 59174 641880 59230 641889
rect 59174 641815 59230 641824
rect 59268 641844 59320 641850
rect 59188 640778 59216 641815
rect 59268 641786 59320 641792
rect 59280 641753 59308 641786
rect 59266 641744 59322 641753
rect 59266 641679 59322 641688
rect 59188 640750 59400 640778
rect 59268 640620 59320 640626
rect 59268 640562 59320 640568
rect 59174 640520 59230 640529
rect 59174 640455 59230 640464
rect 59082 633312 59138 633321
rect 59082 633247 59138 633256
rect 58624 632052 58676 632058
rect 58624 631994 58676 632000
rect 59188 630057 59216 640455
rect 59280 640393 59308 640562
rect 59266 640384 59322 640393
rect 59266 640319 59322 640328
rect 59372 640234 59400 640750
rect 59280 640206 59400 640234
rect 59280 632233 59308 640206
rect 62684 634916 62712 645215
rect 66074 639840 66130 639849
rect 66074 639775 66130 639784
rect 66088 636313 66116 639775
rect 66168 639124 66220 639130
rect 66168 639066 66220 639072
rect 66180 639033 66208 639066
rect 66166 639024 66222 639033
rect 66166 638959 66222 638968
rect 63958 636304 64014 636313
rect 63958 636239 64014 636248
rect 66074 636304 66130 636313
rect 66074 636239 66130 636248
rect 63972 634916 64000 636239
rect 65246 635216 65302 635225
rect 65246 635151 65302 635160
rect 65260 634916 65288 635151
rect 66548 634916 66576 646847
rect 71686 646232 71742 646241
rect 71686 646167 71742 646176
rect 67822 646096 67878 646105
rect 67822 646031 67878 646040
rect 67836 634916 67864 646031
rect 70398 636984 70454 636993
rect 70398 636919 70454 636928
rect 69110 636304 69166 636313
rect 69110 636239 69166 636248
rect 69124 634916 69152 636239
rect 70412 634916 70440 636919
rect 71700 634916 71728 646167
rect 72988 635526 73016 703520
rect 89180 700369 89208 703520
rect 89166 700360 89222 700369
rect 89166 700295 89222 700304
rect 86224 699712 86276 699718
rect 86224 699654 86276 699660
rect 86236 657558 86264 699654
rect 87604 683188 87656 683194
rect 87604 683130 87656 683136
rect 86224 657552 86276 657558
rect 87616 657529 87644 683130
rect 105464 658306 105492 703520
rect 135902 700360 135958 700369
rect 135902 700295 135958 700304
rect 105452 658300 105504 658306
rect 105452 658242 105504 658248
rect 106188 658300 106240 658306
rect 106188 658242 106240 658248
rect 106200 657626 106228 658242
rect 106188 657620 106240 657626
rect 106188 657562 106240 657568
rect 86224 657494 86276 657500
rect 87602 657520 87658 657529
rect 87602 657455 87658 657464
rect 115846 646776 115902 646785
rect 115846 646711 115902 646720
rect 115478 646640 115534 646649
rect 115478 646575 115534 646584
rect 112902 646504 112958 646513
rect 112902 646439 112958 646448
rect 73066 646368 73122 646377
rect 73066 646303 73122 646312
rect 72976 635520 73028 635526
rect 72976 635462 73028 635468
rect 73080 634930 73108 646303
rect 91098 645144 91154 645153
rect 91098 645079 91154 645088
rect 92294 645144 92350 645153
rect 92294 645079 92350 645088
rect 84566 645008 84622 645017
rect 84566 644943 84622 644952
rect 80702 644872 80758 644881
rect 80702 644807 80758 644816
rect 76838 644736 76894 644745
rect 76838 644671 76894 644680
rect 75550 644600 75606 644609
rect 75550 644535 75606 644544
rect 73160 637560 73212 637566
rect 73160 637502 73212 637508
rect 73172 636313 73200 637502
rect 74262 637120 74318 637129
rect 74262 637055 74318 637064
rect 73158 636304 73214 636313
rect 73158 636239 73214 636248
rect 73002 634902 73108 634930
rect 74276 634916 74304 637055
rect 75564 634916 75592 644535
rect 76852 634916 76880 644671
rect 79414 638752 79470 638761
rect 79414 638687 79470 638696
rect 78126 638344 78182 638353
rect 78126 638279 78182 638288
rect 78140 634916 78168 638279
rect 79428 634916 79456 638687
rect 80716 634916 80744 644807
rect 82818 638344 82874 638353
rect 82818 638279 82874 638288
rect 83278 638344 83334 638353
rect 83278 638279 83334 638288
rect 81438 638208 81494 638217
rect 81438 638143 81494 638152
rect 81452 637838 81480 638143
rect 81440 637832 81492 637838
rect 81440 637774 81492 637780
rect 81990 637664 82046 637673
rect 82832 637634 82860 638279
rect 81990 637599 82046 637608
rect 82820 637628 82872 637634
rect 82004 634916 82032 637599
rect 82820 637570 82872 637576
rect 83292 634916 83320 638279
rect 84580 634916 84608 644943
rect 91112 644502 91140 645079
rect 91100 644496 91152 644502
rect 91100 644438 91152 644444
rect 88982 640112 89038 640121
rect 88982 640047 89038 640056
rect 88246 639840 88302 639849
rect 88246 639775 88302 639784
rect 88260 639334 88288 639775
rect 88996 639538 89024 640047
rect 89718 639840 89774 639849
rect 89718 639775 89774 639784
rect 88984 639532 89036 639538
rect 88984 639474 89036 639480
rect 88248 639328 88300 639334
rect 88248 639270 88300 639276
rect 87142 639160 87198 639169
rect 87142 639095 87198 639104
rect 86866 638616 86922 638625
rect 86866 638551 86922 638560
rect 85854 638480 85910 638489
rect 85854 638415 85910 638424
rect 85868 634916 85896 638415
rect 86880 638110 86908 638551
rect 86868 638104 86920 638110
rect 86868 638046 86920 638052
rect 87156 634916 87184 639095
rect 88800 639056 88852 639062
rect 88800 638998 88852 639004
rect 88812 634930 88840 638998
rect 88458 634902 88840 634930
rect 89732 634916 89760 639775
rect 91008 638988 91060 638994
rect 91008 638930 91060 638936
rect 91020 634916 91048 638930
rect 92308 634916 92336 645079
rect 109038 639976 109094 639985
rect 109038 639911 109094 639920
rect 110326 639976 110382 639985
rect 110326 639911 110382 639920
rect 107566 639840 107622 639849
rect 107566 639775 107622 639784
rect 106188 639260 106240 639266
rect 106188 639202 106240 639208
rect 106200 639169 106228 639202
rect 107580 639198 107608 639775
rect 109052 639606 109080 639911
rect 109040 639600 109092 639606
rect 109040 639542 109092 639548
rect 107568 639192 107620 639198
rect 106186 639160 106242 639169
rect 106186 639095 106242 639104
rect 106462 639160 106518 639169
rect 107568 639134 107620 639140
rect 106462 639095 106518 639104
rect 105174 639024 105230 639033
rect 105174 638959 105230 638968
rect 102598 638888 102654 638897
rect 102598 638823 102654 638832
rect 102138 638344 102194 638353
rect 102138 638279 102194 638288
rect 102152 637702 102180 638279
rect 102140 637696 102192 637702
rect 102140 637638 102192 637644
rect 98734 636032 98790 636041
rect 98734 635967 98790 635976
rect 92480 635384 92532 635390
rect 92480 635326 92532 635332
rect 92492 635089 92520 635326
rect 95148 635248 95200 635254
rect 95146 635216 95148 635225
rect 95200 635216 95202 635225
rect 95146 635151 95202 635160
rect 92478 635080 92534 635089
rect 92478 635015 92534 635024
rect 93766 635080 93822 635089
rect 93766 635015 93822 635024
rect 98092 635044 98144 635050
rect 93780 634930 93808 635015
rect 98092 634986 98144 634992
rect 96528 634976 96580 634982
rect 93610 634902 93808 634930
rect 94870 634944 94926 634953
rect 96186 634924 96528 634930
rect 98104 634953 98132 634986
rect 96186 634918 96580 634924
rect 98090 634944 98146 634953
rect 96186 634902 96568 634918
rect 94870 634879 94926 634888
rect 98748 634916 98776 635967
rect 99380 635316 99432 635322
rect 99380 635258 99432 635264
rect 99392 635089 99420 635258
rect 99378 635080 99434 635089
rect 99378 635015 99434 635024
rect 100022 634944 100078 634953
rect 98090 634879 98146 634888
rect 101338 634914 101720 634930
rect 102612 634916 102640 638823
rect 104808 635112 104860 635118
rect 104254 635080 104310 635089
rect 104808 635054 104860 635060
rect 104254 635015 104310 635024
rect 104268 634930 104296 635015
rect 104820 634953 104848 635054
rect 101338 634908 101732 634914
rect 101338 634902 101680 634908
rect 100022 634879 100078 634888
rect 97828 634846 97856 634877
rect 103914 634902 104296 634930
rect 104806 634944 104862 634953
rect 105188 634916 105216 638959
rect 106476 634916 106504 639095
rect 108304 637492 108356 637498
rect 108304 637434 108356 637440
rect 108316 637129 108344 637434
rect 108302 637120 108358 637129
rect 108302 637055 108358 637064
rect 107750 636304 107806 636313
rect 107750 636239 107806 636248
rect 107764 634916 107792 636239
rect 109130 636032 109186 636041
rect 109130 635967 109186 635976
rect 109038 635216 109094 635225
rect 109144 635186 109172 635967
rect 109038 635151 109094 635160
rect 109132 635180 109184 635186
rect 109052 634916 109080 635151
rect 109132 635122 109184 635128
rect 110340 634916 110368 639911
rect 111614 638616 111670 638625
rect 111614 638551 111670 638560
rect 110420 637764 110472 637770
rect 110420 637706 110472 637712
rect 110432 637673 110460 637706
rect 110418 637664 110474 637673
rect 110418 637599 110474 637608
rect 111628 634916 111656 638551
rect 112916 634916 112944 646439
rect 114190 645960 114246 645969
rect 114190 645895 114246 645904
rect 114204 634916 114232 645895
rect 115492 634916 115520 646575
rect 115860 646202 115888 646711
rect 116122 646640 116178 646649
rect 116122 646575 116178 646584
rect 115848 646196 115900 646202
rect 115848 646138 115900 646144
rect 116136 645969 116164 646575
rect 116122 645960 116178 645969
rect 116122 645895 116178 645904
rect 131118 645280 131174 645289
rect 131118 645215 131174 645224
rect 132222 645280 132278 645289
rect 132222 645215 132278 645224
rect 131132 644570 131160 645215
rect 131120 644564 131172 644570
rect 131120 644506 131172 644512
rect 126886 644192 126942 644201
rect 126886 644127 126942 644136
rect 124126 644056 124182 644065
rect 124126 643991 124182 644000
rect 125782 644056 125838 644065
rect 125782 643991 125838 644000
rect 123206 643920 123262 643929
rect 123206 643855 123262 643864
rect 118698 638752 118754 638761
rect 118698 638687 118754 638696
rect 118712 637974 118740 638687
rect 119342 638208 119398 638217
rect 119342 638143 119398 638152
rect 118700 637968 118752 637974
rect 118700 637910 118752 637916
rect 117964 637424 118016 637430
rect 117964 637366 118016 637372
rect 117228 637356 117280 637362
rect 117228 637298 117280 637304
rect 117240 636993 117268 637298
rect 117226 636984 117282 636993
rect 117226 636919 117282 636928
rect 116766 636848 116822 636857
rect 116766 636783 116822 636792
rect 116780 634916 116808 636783
rect 117976 636313 118004 637366
rect 118054 636848 118110 636857
rect 118054 636783 118110 636792
rect 117962 636304 118018 636313
rect 117962 636239 118018 636248
rect 118068 634916 118096 636783
rect 119356 634916 119384 638143
rect 121458 637528 121514 637537
rect 121458 637463 121514 637472
rect 121472 636818 121500 637463
rect 121460 636812 121512 636818
rect 121460 636754 121512 636760
rect 121918 636440 121974 636449
rect 121918 636375 121974 636384
rect 121932 634916 121960 636375
rect 123220 634916 123248 643855
rect 124140 643346 124168 643991
rect 124128 643340 124180 643346
rect 124128 643282 124180 643288
rect 125508 636880 125560 636886
rect 125508 636822 125560 636828
rect 125520 636585 125548 636822
rect 125506 636576 125562 636585
rect 125690 636576 125746 636585
rect 125506 636511 125562 636520
rect 125612 636534 125690 636562
rect 125612 636426 125640 636534
rect 125690 636511 125746 636520
rect 124968 636398 125640 636426
rect 124968 634930 124996 636398
rect 124522 634902 124996 634930
rect 125796 634916 125824 643991
rect 126900 643482 126928 644127
rect 126888 643476 126940 643482
rect 126888 643418 126940 643424
rect 127622 641472 127678 641481
rect 127622 641407 127678 641416
rect 127070 641200 127126 641209
rect 127070 641135 127126 641144
rect 127084 634916 127112 641135
rect 127636 640830 127664 641407
rect 127624 640824 127676 640830
rect 127624 640766 127676 640772
rect 129738 638480 129794 638489
rect 129738 638415 129794 638424
rect 129752 638042 129780 638415
rect 129740 638036 129792 638042
rect 129740 637978 129792 637984
rect 130934 637664 130990 637673
rect 130934 637599 130990 637608
rect 128358 637256 128414 637265
rect 128358 637191 128414 637200
rect 128372 637022 128400 637191
rect 128360 637016 128412 637022
rect 128360 636958 128412 636964
rect 128452 636948 128504 636954
rect 128452 636890 128504 636896
rect 128464 636721 128492 636890
rect 128450 636712 128506 636721
rect 128450 636647 128506 636656
rect 128818 636712 128874 636721
rect 128818 636647 128874 636656
rect 128832 634930 128860 636647
rect 129646 636304 129702 636313
rect 129646 636239 129702 636248
rect 128386 634902 128860 634930
rect 129660 634916 129688 636239
rect 130948 634916 130976 637599
rect 132236 634916 132264 645215
rect 133878 636712 133934 636721
rect 133878 636647 133934 636656
rect 104806 634879 104862 634888
rect 101680 634850 101732 634856
rect 97816 634840 97868 634846
rect 97474 634788 97816 634794
rect 97474 634782 97868 634788
rect 97474 634766 97856 634782
rect 133892 634545 133920 636647
rect 133878 634536 133934 634545
rect 133878 634471 133934 634480
rect 120621 634208 120630 634264
rect 120686 634208 120695 634264
rect 59266 632224 59322 632233
rect 59266 632159 59322 632168
rect 59174 630048 59230 630057
rect 59174 629983 59230 629992
rect 58806 618080 58862 618089
rect 58806 618015 58862 618024
rect 58714 607200 58770 607209
rect 58714 607135 58770 607144
rect 58530 601760 58586 601769
rect 58530 601695 58586 601704
rect 58622 571296 58678 571305
rect 58622 571231 58678 571240
rect 58438 529816 58494 529825
rect 58438 529751 58494 529760
rect 58636 529281 58664 571231
rect 58728 559201 58756 607135
rect 58820 559745 58848 618015
rect 58990 616992 59046 617001
rect 58990 616927 59046 616936
rect 58898 613728 58954 613737
rect 58898 613663 58954 613672
rect 58806 559736 58862 559745
rect 58806 559671 58862 559680
rect 58714 559192 58770 559201
rect 58714 559127 58770 559136
rect 58806 558104 58862 558113
rect 58806 558039 58862 558048
rect 58622 529272 58678 529281
rect 58622 529207 58678 529216
rect 58624 525904 58676 525910
rect 58624 525846 58676 525852
rect 58440 521552 58492 521558
rect 58440 521494 58492 521500
rect 57980 520464 58032 520470
rect 57980 520406 58032 520412
rect 57886 513904 57942 513913
rect 57886 513839 57942 513848
rect 57992 513330 58020 520406
rect 57980 513324 58032 513330
rect 57980 513266 58032 513272
rect 57888 511964 57940 511970
rect 57888 511906 57940 511912
rect 57796 507884 57848 507890
rect 57796 507826 57848 507832
rect 57704 500948 57756 500954
rect 57704 500890 57756 500896
rect 57612 499044 57664 499050
rect 57612 498986 57664 498992
rect 57532 498902 57744 498930
rect 57612 498840 57664 498846
rect 57518 498808 57574 498817
rect 57612 498782 57664 498788
rect 57518 498743 57574 498752
rect 57532 498137 57560 498743
rect 57518 498128 57574 498137
rect 57518 498063 57574 498072
rect 57518 496360 57574 496369
rect 57518 496295 57574 496304
rect 57532 492697 57560 496295
rect 57518 492688 57574 492697
rect 57518 492623 57574 492632
rect 57520 491632 57572 491638
rect 57520 491574 57572 491580
rect 57532 437753 57560 491574
rect 57624 486713 57652 498782
rect 57716 496330 57744 498902
rect 57704 496324 57756 496330
rect 57704 496266 57756 496272
rect 57702 496224 57758 496233
rect 57702 496159 57758 496168
rect 57716 491065 57744 496159
rect 57702 491056 57758 491065
rect 57702 490991 57758 491000
rect 57808 488646 57836 507826
rect 57796 488640 57848 488646
rect 57796 488582 57848 488588
rect 57704 488572 57756 488578
rect 57704 488514 57756 488520
rect 57610 486704 57666 486713
rect 57610 486639 57666 486648
rect 57518 437744 57574 437753
rect 57518 437679 57574 437688
rect 57716 429214 57744 488514
rect 57704 429208 57756 429214
rect 57704 429150 57756 429156
rect 57520 400920 57572 400926
rect 57520 400862 57572 400868
rect 57532 390114 57560 400862
rect 57520 390108 57572 390114
rect 57520 390050 57572 390056
rect 57428 366648 57480 366654
rect 57428 366590 57480 366596
rect 57900 361214 57928 511906
rect 57980 509924 58032 509930
rect 57980 509866 58032 509872
rect 57992 493338 58020 509866
rect 58452 503674 58480 521494
rect 58532 513324 58584 513330
rect 58532 513266 58584 513272
rect 58544 504422 58572 513266
rect 58636 511290 58664 525846
rect 58716 519036 58768 519042
rect 58716 518978 58768 518984
rect 58624 511284 58676 511290
rect 58624 511226 58676 511232
rect 58728 507890 58756 518978
rect 58716 507884 58768 507890
rect 58716 507826 58768 507832
rect 58532 504416 58584 504422
rect 58532 504358 58584 504364
rect 58440 503668 58492 503674
rect 58440 503610 58492 503616
rect 58624 503124 58676 503130
rect 58624 503066 58676 503072
rect 58072 500948 58124 500954
rect 58072 500890 58124 500896
rect 57980 493332 58032 493338
rect 57980 493274 58032 493280
rect 58084 488578 58112 500890
rect 58072 488572 58124 488578
rect 58072 488514 58124 488520
rect 58532 429208 58584 429214
rect 58532 429150 58584 429156
rect 58544 390182 58572 429150
rect 58532 390176 58584 390182
rect 58532 390118 58584 390124
rect 58636 361282 58664 503066
rect 58716 494760 58768 494766
rect 58716 494702 58768 494708
rect 58624 361276 58676 361282
rect 58624 361218 58676 361224
rect 57888 361208 57940 361214
rect 57888 361150 57940 361156
rect 57336 358284 57388 358290
rect 57336 358226 57388 358232
rect 58728 355706 58756 494702
rect 58820 491201 58848 558039
rect 58912 529145 58940 613663
rect 59004 544377 59032 616927
rect 59726 608288 59782 608297
rect 59726 608223 59782 608232
rect 59634 569120 59690 569129
rect 59634 569055 59690 569064
rect 59266 565856 59322 565865
rect 59188 565814 59266 565842
rect 59188 557534 59216 565814
rect 59266 565791 59322 565800
rect 59542 561436 59598 561445
rect 59542 561371 59598 561380
rect 59556 560318 59584 561371
rect 59544 560312 59596 560318
rect 59544 560254 59596 560260
rect 59268 558680 59320 558686
rect 59268 558622 59320 558628
rect 59280 557841 59308 558622
rect 59266 557832 59322 557841
rect 59266 557767 59322 557776
rect 59188 557506 59308 557534
rect 59176 553376 59228 553382
rect 59176 553318 59228 553324
rect 59188 552673 59216 553318
rect 59174 552664 59230 552673
rect 59174 552599 59230 552608
rect 59174 551440 59230 551449
rect 59174 551375 59230 551384
rect 59082 548312 59138 548321
rect 59082 548247 59138 548256
rect 58990 544368 59046 544377
rect 58990 544303 59046 544312
rect 58990 534440 59046 534449
rect 58990 534375 59046 534384
rect 58898 529136 58954 529145
rect 58898 529071 58954 529080
rect 58900 523728 58952 523734
rect 58900 523670 58952 523676
rect 58806 491192 58862 491201
rect 58806 491127 58862 491136
rect 58808 488640 58860 488646
rect 58808 488582 58860 488588
rect 58716 355700 58768 355706
rect 58716 355642 58768 355648
rect 57244 355632 57296 355638
rect 57244 355574 57296 355580
rect 58820 355434 58848 488582
rect 58912 429049 58940 523670
rect 59004 430137 59032 534375
rect 58990 430128 59046 430137
rect 58990 430063 59046 430072
rect 58898 429040 58954 429049
rect 58898 428975 58954 428984
rect 59096 427961 59124 548247
rect 59082 427952 59138 427961
rect 59082 427887 59138 427896
rect 59188 423609 59216 551375
rect 59280 538937 59308 557506
rect 59648 554033 59676 569055
rect 59634 554024 59690 554033
rect 59634 553959 59690 553968
rect 59740 548593 59768 608223
rect 59818 606112 59874 606121
rect 59818 606047 59874 606056
rect 59832 605834 59860 606047
rect 59832 605806 59952 605834
rect 59818 602848 59874 602857
rect 59818 602783 59874 602792
rect 59726 548584 59782 548593
rect 59726 548519 59782 548528
rect 59266 538928 59322 538937
rect 59266 538863 59322 538872
rect 59832 536761 59860 602783
rect 59818 536752 59874 536761
rect 59818 536687 59874 536696
rect 59636 532704 59688 532710
rect 59636 532646 59688 532652
rect 59648 531593 59676 532646
rect 59924 532545 59952 605806
rect 134524 591388 134576 591394
rect 134524 591330 134576 591336
rect 60740 560312 60792 560318
rect 60646 560280 60702 560289
rect 60740 560254 60792 560260
rect 60646 560215 60702 560224
rect 60660 559298 60688 560215
rect 60648 559292 60700 559298
rect 60648 559234 60700 559240
rect 60004 554668 60056 554674
rect 60004 554610 60056 554616
rect 60016 553761 60044 554610
rect 60002 553752 60058 553761
rect 60002 553687 60058 553696
rect 60096 549976 60148 549982
rect 60096 549918 60148 549924
rect 59910 532536 59966 532545
rect 59910 532471 59966 532480
rect 59634 531584 59690 531593
rect 59634 531519 59690 531528
rect 59820 527604 59872 527610
rect 59820 527546 59872 527552
rect 59268 527536 59320 527542
rect 59268 527478 59320 527484
rect 59280 521014 59308 527478
rect 59634 527232 59690 527241
rect 59634 527167 59690 527176
rect 59452 526448 59504 526454
rect 59452 526390 59504 526396
rect 59360 521620 59412 521626
rect 59360 521562 59412 521568
rect 59268 521008 59320 521014
rect 59268 520950 59320 520956
rect 59268 520668 59320 520674
rect 59268 520610 59320 520616
rect 59280 519489 59308 520610
rect 59266 519480 59322 519489
rect 59266 519415 59322 519424
rect 59372 516186 59400 521562
rect 59464 521558 59492 526390
rect 59544 522980 59596 522986
rect 59544 522922 59596 522928
rect 59452 521552 59504 521558
rect 59452 521494 59504 521500
rect 59452 520600 59504 520606
rect 59452 520542 59504 520548
rect 59360 516180 59412 516186
rect 59360 516122 59412 516128
rect 59464 511970 59492 520542
rect 59452 511964 59504 511970
rect 59452 511906 59504 511912
rect 59556 509234 59584 522922
rect 59648 521234 59676 527167
rect 59728 526380 59780 526386
rect 59728 526322 59780 526328
rect 59740 521558 59768 526322
rect 59832 522442 59860 527546
rect 60002 523016 60058 523025
rect 59924 522974 60002 523002
rect 59820 522436 59872 522442
rect 59820 522378 59872 522384
rect 59728 521552 59780 521558
rect 59728 521494 59780 521500
rect 59648 521206 59768 521234
rect 59636 521076 59688 521082
rect 59636 521018 59688 521024
rect 59648 520198 59676 521018
rect 59740 520674 59768 521206
rect 59820 520940 59872 520946
rect 59820 520882 59872 520888
rect 59728 520668 59780 520674
rect 59728 520610 59780 520616
rect 59728 520396 59780 520402
rect 59728 520338 59780 520344
rect 59636 520192 59688 520198
rect 59636 520134 59688 520140
rect 59740 520033 59768 520338
rect 59832 520198 59860 520882
rect 59820 520192 59872 520198
rect 59820 520134 59872 520140
rect 59726 520024 59782 520033
rect 59726 519959 59782 519968
rect 59818 519888 59874 519897
rect 59818 519823 59874 519832
rect 59832 518265 59860 519823
rect 59924 519466 59952 522974
rect 60002 522951 60058 522960
rect 60004 520668 60056 520674
rect 60004 520610 60056 520616
rect 60016 519586 60044 520610
rect 60004 519580 60056 519586
rect 60004 519522 60056 519528
rect 59924 519438 60044 519466
rect 59818 518256 59874 518265
rect 59818 518191 59874 518200
rect 59556 509206 59952 509234
rect 59360 505164 59412 505170
rect 59360 505106 59412 505112
rect 59372 503690 59400 505106
rect 59280 503662 59400 503690
rect 59820 503668 59872 503674
rect 59174 423600 59230 423609
rect 59174 423535 59230 423544
rect 59280 361350 59308 503662
rect 59820 503610 59872 503616
rect 59832 500206 59860 503610
rect 59820 500200 59872 500206
rect 59820 500142 59872 500148
rect 59924 390697 59952 509206
rect 60016 500585 60044 519438
rect 60108 517993 60136 549918
rect 60752 534954 60780 560254
rect 61384 556844 61436 556850
rect 61384 556786 61436 556792
rect 60832 553104 60884 553110
rect 60832 553046 60884 553052
rect 60844 552401 60872 553046
rect 60830 552392 60886 552401
rect 60830 552327 60886 552336
rect 60832 539572 60884 539578
rect 60832 539514 60884 539520
rect 60844 538801 60872 539514
rect 60830 538792 60886 538801
rect 60830 538727 60886 538736
rect 60740 534948 60792 534954
rect 60740 534890 60792 534896
rect 60188 530324 60240 530330
rect 60188 530266 60240 530272
rect 60200 520470 60228 530266
rect 60280 530052 60332 530058
rect 60280 529994 60332 530000
rect 60188 520464 60240 520470
rect 60188 520406 60240 520412
rect 60188 520124 60240 520130
rect 60188 520066 60240 520072
rect 60094 517984 60150 517993
rect 60094 517919 60150 517928
rect 60200 505345 60228 520066
rect 60186 505336 60242 505345
rect 60186 505271 60242 505280
rect 60188 504416 60240 504422
rect 60188 504358 60240 504364
rect 60096 501628 60148 501634
rect 60096 501570 60148 501576
rect 60002 500576 60058 500585
rect 60002 500511 60058 500520
rect 60108 500426 60136 501570
rect 60016 500398 60136 500426
rect 59910 390688 59966 390697
rect 59910 390623 59966 390632
rect 59268 361344 59320 361350
rect 59268 361286 59320 361292
rect 58808 355428 58860 355434
rect 58808 355370 58860 355376
rect 56140 352912 56192 352918
rect 56140 352854 56192 352860
rect 55864 350192 55916 350198
rect 55864 350134 55916 350140
rect 50620 347200 50672 347206
rect 50620 347142 50672 347148
rect 47952 347132 48004 347138
rect 47952 347074 48004 347080
rect 60016 342922 60044 500398
rect 60200 500290 60228 504358
rect 60108 500262 60228 500290
rect 60108 355774 60136 500262
rect 60188 500200 60240 500206
rect 60188 500142 60240 500148
rect 60200 358358 60228 500142
rect 60292 497185 60320 529994
rect 61108 529236 61160 529242
rect 61108 529178 61160 529184
rect 60832 527944 60884 527950
rect 60832 527886 60884 527892
rect 60556 527468 60608 527474
rect 60556 527410 60608 527416
rect 60372 525836 60424 525842
rect 60372 525778 60424 525784
rect 60278 497176 60334 497185
rect 60278 497111 60334 497120
rect 60280 496324 60332 496330
rect 60280 496266 60332 496272
rect 60292 364274 60320 496266
rect 60384 391678 60412 525778
rect 60568 521490 60596 527410
rect 60740 524952 60792 524958
rect 60740 524894 60792 524900
rect 60752 523274 60780 524894
rect 60660 523246 60780 523274
rect 60556 521484 60608 521490
rect 60556 521426 60608 521432
rect 60556 520396 60608 520402
rect 60556 520338 60608 520344
rect 60464 520192 60516 520198
rect 60464 520134 60516 520140
rect 60372 391672 60424 391678
rect 60372 391614 60424 391620
rect 60280 364268 60332 364274
rect 60280 364210 60332 364216
rect 60476 361418 60504 520134
rect 60464 361412 60516 361418
rect 60464 361354 60516 361360
rect 60188 358352 60240 358358
rect 60188 358294 60240 358300
rect 60096 355768 60148 355774
rect 60096 355710 60148 355716
rect 60568 353122 60596 520338
rect 60660 520062 60688 523246
rect 60740 523184 60792 523190
rect 60740 523126 60792 523132
rect 60752 522374 60780 523126
rect 60844 522986 60872 527886
rect 60832 522980 60884 522986
rect 60832 522922 60884 522928
rect 60740 522368 60792 522374
rect 60740 522310 60792 522316
rect 61120 522050 61148 529178
rect 61396 524414 61424 556786
rect 61488 539209 61516 560116
rect 61566 552664 61622 552673
rect 61566 552599 61622 552608
rect 61474 539200 61530 539209
rect 61474 539135 61530 539144
rect 61580 529242 61608 552599
rect 62500 535129 62528 560116
rect 63512 549001 63540 560116
rect 63592 558612 63644 558618
rect 63592 558554 63644 558560
rect 63604 558113 63632 558554
rect 64524 558249 64552 560116
rect 64510 558240 64566 558249
rect 64510 558175 64566 558184
rect 63590 558104 63646 558113
rect 63590 558039 63646 558048
rect 63498 548992 63554 549001
rect 63498 548927 63554 548936
rect 62486 535120 62542 535129
rect 62486 535055 62542 535064
rect 63592 534744 63644 534750
rect 63592 534686 63644 534692
rect 63604 534074 63632 534686
rect 63512 534046 63632 534074
rect 62856 531276 62908 531282
rect 62856 531218 62908 531224
rect 62764 530188 62816 530194
rect 62764 530130 62816 530136
rect 61568 529236 61620 529242
rect 61568 529178 61620 529184
rect 61568 527672 61620 527678
rect 61568 527614 61620 527620
rect 60752 522022 61148 522050
rect 61304 524386 61424 524414
rect 60648 520056 60700 520062
rect 60648 519998 60700 520004
rect 60646 519888 60702 519897
rect 60752 519874 60780 522022
rect 60924 521960 60976 521966
rect 60924 521902 60976 521908
rect 60832 521892 60884 521898
rect 60832 521834 60884 521840
rect 60702 519846 60780 519874
rect 60646 519823 60702 519832
rect 60646 519616 60702 519625
rect 60844 519602 60872 521834
rect 60702 519574 60872 519602
rect 60936 519586 60964 521902
rect 61108 521892 61160 521898
rect 61108 521834 61160 521840
rect 61120 520266 61148 521834
rect 61108 520260 61160 520266
rect 61108 520202 61160 520208
rect 61200 520260 61252 520266
rect 61200 520202 61252 520208
rect 60924 519580 60976 519586
rect 60646 519551 60702 519560
rect 60924 519522 60976 519528
rect 60832 519512 60884 519518
rect 61212 519466 61240 520202
rect 60884 519460 61240 519466
rect 60832 519454 61240 519460
rect 60844 519438 61240 519454
rect 60646 519344 60702 519353
rect 60702 519302 60872 519330
rect 60646 519279 60702 519288
rect 60844 519194 60872 519302
rect 61304 519194 61332 524386
rect 60844 519166 61332 519194
rect 60648 519104 60700 519110
rect 61580 519058 61608 527614
rect 61660 527400 61712 527406
rect 61660 527342 61712 527348
rect 61672 520470 61700 527342
rect 62028 527128 62080 527134
rect 62028 527070 62080 527076
rect 62040 526697 62068 527070
rect 62026 526688 62082 526697
rect 62026 526623 62082 526632
rect 61844 526312 61896 526318
rect 61844 526254 61896 526260
rect 61750 526144 61806 526153
rect 61750 526079 61806 526088
rect 61660 520464 61712 520470
rect 61660 520406 61712 520412
rect 61764 520130 61792 526079
rect 61856 521082 61884 526254
rect 62028 524884 62080 524890
rect 62028 524826 62080 524832
rect 61844 521076 61896 521082
rect 61844 521018 61896 521024
rect 61842 520296 61898 520305
rect 61842 520231 61844 520240
rect 61896 520231 61898 520240
rect 61844 520202 61896 520208
rect 62040 520198 62068 524826
rect 62776 520946 62804 530130
rect 62868 521626 62896 531218
rect 63512 529938 63540 534046
rect 65536 533225 65564 560116
rect 66548 547641 66576 560116
rect 67560 551721 67588 560116
rect 68282 558240 68338 558249
rect 68282 558175 68338 558184
rect 67546 551712 67602 551721
rect 67546 551647 67602 551656
rect 67548 547868 67600 547874
rect 67548 547810 67600 547816
rect 66534 547632 66590 547641
rect 66534 547567 66590 547576
rect 67560 546961 67588 547810
rect 67546 546952 67602 546961
rect 67546 546887 67602 546896
rect 66260 536784 66312 536790
rect 66260 536726 66312 536732
rect 66272 534074 66300 536726
rect 66180 534046 66300 534074
rect 65522 533216 65578 533225
rect 65522 533151 65578 533160
rect 66180 531350 66208 534046
rect 66168 531344 66220 531350
rect 66168 531286 66220 531292
rect 63420 529910 63540 529938
rect 63420 525842 63448 529910
rect 63408 525836 63460 525842
rect 63408 525778 63460 525784
rect 68296 524249 68324 558175
rect 68572 537849 68600 560116
rect 68558 537840 68614 537849
rect 68558 537775 68614 537784
rect 69020 536784 69072 536790
rect 69020 536726 69072 536732
rect 69032 534750 69060 536726
rect 69020 534744 69072 534750
rect 69020 534686 69072 534692
rect 69020 525768 69072 525774
rect 69020 525710 69072 525716
rect 69032 525065 69060 525710
rect 69584 525609 69612 560116
rect 70400 525700 70452 525706
rect 70400 525642 70452 525648
rect 69570 525600 69626 525609
rect 69570 525535 69626 525544
rect 69018 525056 69074 525065
rect 69018 524991 69074 525000
rect 70412 524929 70440 525642
rect 70596 525337 70624 560116
rect 71608 543425 71636 560116
rect 72424 543720 72476 543726
rect 72424 543662 72476 543668
rect 71594 543416 71650 543425
rect 71594 543351 71650 543360
rect 72436 536926 72464 543662
rect 72620 542065 72648 560116
rect 72606 542056 72662 542065
rect 72606 541991 72662 542000
rect 73632 540705 73660 560116
rect 74644 546281 74672 560116
rect 74630 546272 74686 546281
rect 74630 546207 74686 546216
rect 75656 545057 75684 560116
rect 75920 550588 75972 550594
rect 75920 550530 75972 550536
rect 75828 546372 75880 546378
rect 75828 546314 75880 546320
rect 75840 545601 75868 546314
rect 75826 545592 75882 545601
rect 75826 545527 75882 545536
rect 75932 545306 75960 550530
rect 75748 545278 75960 545306
rect 75642 545048 75698 545057
rect 75642 544983 75698 544992
rect 75748 543794 75776 545278
rect 75828 545080 75880 545086
rect 75828 545022 75880 545028
rect 75840 544649 75868 545022
rect 75826 544640 75882 544649
rect 75826 544575 75882 544584
rect 75736 543788 75788 543794
rect 75736 543730 75788 543736
rect 73618 540696 73674 540705
rect 73618 540631 73674 540640
rect 73160 540252 73212 540258
rect 73160 540194 73212 540200
rect 72424 536920 72476 536926
rect 72424 536862 72476 536868
rect 73172 536858 73200 540194
rect 73160 536852 73212 536858
rect 73160 536794 73212 536800
rect 76668 536353 76696 560116
rect 77300 546508 77352 546514
rect 77300 546450 77352 546456
rect 77312 540258 77340 546450
rect 77300 540252 77352 540258
rect 77300 540194 77352 540200
rect 76654 536344 76710 536353
rect 76654 536279 76710 536288
rect 70582 525328 70638 525337
rect 70582 525263 70638 525272
rect 71964 524952 72016 524958
rect 70398 524920 70454 524929
rect 71964 524894 72016 524900
rect 70398 524855 70454 524864
rect 71872 524476 71924 524482
rect 71872 524418 71924 524424
rect 68928 524340 68980 524346
rect 68928 524282 68980 524288
rect 68282 524240 68338 524249
rect 68282 524175 68338 524184
rect 68940 523433 68968 524282
rect 69664 523592 69716 523598
rect 69664 523534 69716 523540
rect 68926 523424 68982 523433
rect 68926 523359 68982 523368
rect 68928 523048 68980 523054
rect 68928 522990 68980 522996
rect 68940 522442 68968 522990
rect 69676 522578 69704 523534
rect 71780 523456 71832 523462
rect 71780 523398 71832 523404
rect 70400 522640 70452 522646
rect 70400 522582 70452 522588
rect 69388 522572 69440 522578
rect 69388 522514 69440 522520
rect 69664 522572 69716 522578
rect 69664 522514 69716 522520
rect 68928 522436 68980 522442
rect 68928 522378 68980 522384
rect 67364 522300 67416 522306
rect 67364 522242 67416 522248
rect 62856 521620 62908 521626
rect 62856 521562 62908 521568
rect 62764 520940 62816 520946
rect 62764 520882 62816 520888
rect 62120 520464 62172 520470
rect 62120 520406 62172 520412
rect 62028 520192 62080 520198
rect 62132 520169 62160 520406
rect 62028 520134 62080 520140
rect 62118 520160 62174 520169
rect 61752 520124 61804 520130
rect 67376 520146 67404 522242
rect 68376 522232 68428 522238
rect 68376 522174 68428 522180
rect 68388 520146 68416 522174
rect 69400 520146 69428 522514
rect 70412 520146 70440 522582
rect 71792 522306 71820 523398
rect 71780 522300 71832 522306
rect 71780 522242 71832 522248
rect 71884 521014 71912 524418
rect 71872 521008 71924 521014
rect 71872 520950 71924 520956
rect 71976 520946 72004 524894
rect 77680 523977 77708 560116
rect 78588 554804 78640 554810
rect 78588 554746 78640 554752
rect 78600 550594 78628 554746
rect 78588 550588 78640 550594
rect 78588 550530 78640 550536
rect 78692 549137 78720 560116
rect 79600 549908 79652 549914
rect 79600 549850 79652 549856
rect 79324 549228 79376 549234
rect 79324 549170 79376 549176
rect 78678 549128 78734 549137
rect 78678 549063 78734 549072
rect 79336 548457 79364 549170
rect 79322 548448 79378 548457
rect 79322 548383 79378 548392
rect 79612 546514 79640 549850
rect 79600 546508 79652 546514
rect 79600 546450 79652 546456
rect 79704 540977 79732 560116
rect 80060 550588 80112 550594
rect 80060 550530 80112 550536
rect 80072 550089 80100 550530
rect 80716 550225 80744 560116
rect 81440 552016 81492 552022
rect 81440 551958 81492 551964
rect 81452 551449 81480 551958
rect 81438 551440 81494 551449
rect 81438 551375 81494 551384
rect 81728 551177 81756 560116
rect 81714 551168 81770 551177
rect 81714 551103 81770 551112
rect 80702 550216 80758 550225
rect 80702 550151 80758 550160
rect 80058 550080 80114 550089
rect 80058 550015 80114 550024
rect 82740 543697 82768 560116
rect 82726 543688 82782 543697
rect 82726 543623 82782 543632
rect 82820 542360 82872 542366
rect 83752 542337 83780 560116
rect 82820 542302 82872 542308
rect 83738 542328 83794 542337
rect 82832 541521 82860 542302
rect 83738 542263 83794 542272
rect 82818 541512 82874 541521
rect 82818 541447 82874 541456
rect 79690 540968 79746 540977
rect 79690 540903 79746 540912
rect 84764 537305 84792 560116
rect 85776 539345 85804 560116
rect 86788 545601 86816 560116
rect 86868 556232 86920 556238
rect 86868 556174 86920 556180
rect 86880 554810 86908 556174
rect 86868 554804 86920 554810
rect 86868 554746 86920 554752
rect 86868 546304 86920 546310
rect 86868 546246 86920 546252
rect 86774 545592 86830 545601
rect 86774 545527 86830 545536
rect 86880 545465 86908 546246
rect 86866 545456 86922 545465
rect 86866 545391 86922 545400
rect 87800 544082 87828 560116
rect 88812 547777 88840 560116
rect 89628 558544 89680 558550
rect 89628 558486 89680 558492
rect 89640 556238 89668 558486
rect 89628 556232 89680 556238
rect 89628 556174 89680 556180
rect 88984 552220 89036 552226
rect 88984 552162 89036 552168
rect 88996 549914 89024 552162
rect 88984 549908 89036 549914
rect 88984 549850 89036 549856
rect 88984 547800 89036 547806
rect 88798 547768 88854 547777
rect 88984 547742 89036 547748
rect 88798 547703 88854 547712
rect 88996 546825 89024 547742
rect 88982 546816 89038 546825
rect 88982 546751 89038 546760
rect 88248 545012 88300 545018
rect 88248 544954 88300 544960
rect 88260 544241 88288 544954
rect 88246 544232 88302 544241
rect 88430 544232 88486 544241
rect 88246 544167 88302 544176
rect 88352 544190 88430 544218
rect 88352 544082 88380 544190
rect 88430 544167 88486 544176
rect 87800 544054 88380 544082
rect 88616 539640 88668 539646
rect 88616 539582 88668 539588
rect 86868 539504 86920 539510
rect 86868 539446 86920 539452
rect 85762 539336 85818 539345
rect 85762 539271 85818 539280
rect 86880 538665 86908 539446
rect 86866 538656 86922 538665
rect 86866 538591 86922 538600
rect 85488 538212 85540 538218
rect 85488 538154 85540 538160
rect 84750 537296 84806 537305
rect 84750 537231 84806 537240
rect 85500 537169 85528 538154
rect 85486 537160 85542 537169
rect 85486 537095 85542 537104
rect 84568 536852 84620 536858
rect 84568 536794 84620 536800
rect 83556 532772 83608 532778
rect 83556 532714 83608 532720
rect 80794 528048 80850 528057
rect 80624 528006 80794 528034
rect 78588 524272 78640 524278
rect 78588 524214 78640 524220
rect 77666 523968 77722 523977
rect 77666 523903 77722 523912
rect 78600 523297 78628 524214
rect 78586 523288 78642 523297
rect 78586 523223 78642 523232
rect 77484 522164 77536 522170
rect 77484 522106 77536 522112
rect 73344 521280 73396 521286
rect 73344 521222 73396 521228
rect 71964 520940 72016 520946
rect 71964 520882 72016 520888
rect 71320 520872 71372 520878
rect 71320 520814 71372 520820
rect 71332 520146 71360 520814
rect 72332 520328 72384 520334
rect 72332 520270 72384 520276
rect 72344 520146 72372 520270
rect 73356 520146 73384 521222
rect 74448 521212 74500 521218
rect 74448 521154 74500 521160
rect 74460 520146 74488 521154
rect 76472 520804 76524 520810
rect 76472 520746 76524 520752
rect 75368 520736 75420 520742
rect 75368 520678 75420 520684
rect 75380 520146 75408 520678
rect 76484 520146 76512 520746
rect 77496 520146 77524 522106
rect 78496 522096 78548 522102
rect 78496 522038 78548 522044
rect 78508 520146 78536 522038
rect 79416 521688 79468 521694
rect 79416 521630 79468 521636
rect 79428 520146 79456 521630
rect 80624 520146 80652 528006
rect 80794 527983 80850 527992
rect 82728 525836 82780 525842
rect 82728 525778 82780 525784
rect 81624 521688 81676 521694
rect 81624 521630 81676 521636
rect 81636 520146 81664 521630
rect 82740 520146 82768 525778
rect 67376 520118 67420 520146
rect 68388 520118 68432 520146
rect 69400 520118 69444 520146
rect 70412 520118 70456 520146
rect 71332 520118 71468 520146
rect 72344 520118 72480 520146
rect 73356 520118 73492 520146
rect 74460 520118 74504 520146
rect 75380 520118 75516 520146
rect 76484 520118 76528 520146
rect 77496 520118 77540 520146
rect 78508 520118 78552 520146
rect 79428 520118 79564 520146
rect 62118 520095 62174 520104
rect 61752 520066 61804 520072
rect 67392 519860 67420 520118
rect 68404 519860 68432 520118
rect 69416 519860 69444 520118
rect 70428 519860 70456 520118
rect 71440 519860 71468 520118
rect 72452 519860 72480 520118
rect 73464 519860 73492 520118
rect 74476 519860 74504 520118
rect 75488 519860 75516 520118
rect 76500 519860 76528 520118
rect 77512 519860 77540 520118
rect 78524 519860 78552 520118
rect 79536 519860 79564 520118
rect 80548 520118 80652 520146
rect 81560 520118 81664 520146
rect 82572 520118 82768 520146
rect 83568 520146 83596 532714
rect 84580 520146 84608 536794
rect 85580 535492 85632 535498
rect 85580 535434 85632 535440
rect 85592 520146 85620 535434
rect 87696 524476 87748 524482
rect 87696 524418 87748 524424
rect 86684 520328 86736 520334
rect 86684 520270 86736 520276
rect 86696 520146 86724 520270
rect 87708 520146 87736 524418
rect 83568 520118 83612 520146
rect 84580 520118 84624 520146
rect 85592 520118 85636 520146
rect 80548 519860 80576 520118
rect 81560 519860 81588 520118
rect 82572 519860 82600 520118
rect 83584 519860 83612 520118
rect 84596 519860 84624 520118
rect 85608 519860 85636 520118
rect 86620 520118 86724 520146
rect 87632 520118 87736 520146
rect 88628 520146 88656 539582
rect 89720 536784 89772 536790
rect 89720 536726 89772 536732
rect 89732 535945 89760 536726
rect 89718 535936 89774 535945
rect 89718 535871 89774 535880
rect 89824 534585 89852 560116
rect 90640 546508 90692 546514
rect 90640 546450 90692 546456
rect 89810 534576 89866 534585
rect 89810 534511 89866 534520
rect 89628 522368 89680 522374
rect 89628 522310 89680 522316
rect 89640 520146 89668 522310
rect 90652 520146 90680 546450
rect 90836 536489 90864 560116
rect 91192 559564 91244 559570
rect 91192 559506 91244 559512
rect 91204 558550 91232 559506
rect 91192 558544 91244 558550
rect 91192 558486 91244 558492
rect 91100 556912 91152 556918
rect 91100 556854 91152 556860
rect 91112 552226 91140 556854
rect 91100 552220 91152 552226
rect 91100 552162 91152 552168
rect 91652 542428 91704 542434
rect 91652 542370 91704 542376
rect 91100 540932 91152 540938
rect 91100 540874 91152 540880
rect 91112 540025 91140 540874
rect 91098 540016 91154 540025
rect 91098 539951 91154 539960
rect 90822 536480 90878 536489
rect 90822 536415 90878 536424
rect 91664 520146 91692 542370
rect 91848 540161 91876 560116
rect 92480 550452 92532 550458
rect 92480 550394 92532 550400
rect 92492 549817 92520 550394
rect 92860 550089 92888 560116
rect 92846 550080 92902 550089
rect 92846 550015 92902 550024
rect 92478 549808 92534 549817
rect 92478 549743 92534 549752
rect 93676 547936 93728 547942
rect 93676 547878 93728 547884
rect 92664 541000 92716 541006
rect 92664 540942 92716 540948
rect 92020 540252 92072 540258
rect 92020 540194 92072 540200
rect 91834 540152 91890 540161
rect 91834 540087 91890 540096
rect 92032 528554 92060 540194
rect 91756 528526 92060 528554
rect 91756 527882 91784 528526
rect 91744 527876 91796 527882
rect 91744 527818 91796 527824
rect 92676 520146 92704 540942
rect 93688 520146 93716 547878
rect 93872 529553 93900 560116
rect 94688 543788 94740 543794
rect 94688 543730 94740 543736
rect 93858 529544 93914 529553
rect 93858 529479 93914 529488
rect 94700 520146 94728 543730
rect 94884 528873 94912 560116
rect 95148 529780 95200 529786
rect 95148 529722 95200 529728
rect 95056 529712 95108 529718
rect 95056 529654 95108 529660
rect 94870 528864 94926 528873
rect 94870 528799 94926 528808
rect 95068 528737 95096 529654
rect 95160 529009 95188 529722
rect 95896 529689 95924 560116
rect 96528 529848 96580 529854
rect 96528 529790 96580 529796
rect 95882 529680 95938 529689
rect 95882 529615 95938 529624
rect 95514 529544 95570 529553
rect 95514 529479 95570 529488
rect 95146 529000 95202 529009
rect 95146 528935 95202 528944
rect 95528 528873 95556 529479
rect 96540 529417 96568 529790
rect 96526 529408 96582 529417
rect 96526 529343 96582 529352
rect 96908 529242 96936 560116
rect 97828 560102 97934 560130
rect 97828 553217 97856 560102
rect 98644 553240 98696 553246
rect 97814 553208 97870 553217
rect 98644 553182 98696 553188
rect 97814 553143 97870 553152
rect 97908 553172 97960 553178
rect 97908 553114 97960 553120
rect 97920 553081 97948 553114
rect 97906 553072 97962 553081
rect 97906 553007 97962 553016
rect 98656 552265 98684 553182
rect 98932 553081 98960 560116
rect 98918 553072 98974 553081
rect 98918 553007 98974 553016
rect 98642 552256 98698 552265
rect 98642 552191 98698 552200
rect 99380 550520 99432 550526
rect 99380 550462 99432 550468
rect 99392 549681 99420 550462
rect 99944 550361 99972 560116
rect 99930 550352 99986 550361
rect 99930 550287 99986 550296
rect 99378 549672 99434 549681
rect 99378 549607 99434 549616
rect 100760 539436 100812 539442
rect 100760 539378 100812 539384
rect 100772 538529 100800 539378
rect 100758 538520 100814 538529
rect 100758 538455 100814 538464
rect 100760 535424 100812 535430
rect 100760 535366 100812 535372
rect 100772 534449 100800 535366
rect 100956 535265 100984 560116
rect 101968 538529 101996 560116
rect 101954 538520 102010 538529
rect 101954 538455 102010 538464
rect 100942 535256 100998 535265
rect 100942 535191 100998 535200
rect 100758 534440 100814 534449
rect 100758 534375 100814 534384
rect 96896 529236 96948 529242
rect 96896 529178 96948 529184
rect 95514 528864 95570 528873
rect 95514 528799 95570 528808
rect 95054 528728 95110 528737
rect 95054 528663 95110 528672
rect 102980 527785 103008 560116
rect 103992 539073 104020 560116
rect 104900 558204 104952 558210
rect 104900 558146 104952 558152
rect 104912 556918 104940 558146
rect 104900 556912 104952 556918
rect 104900 556854 104952 556860
rect 104806 539472 104862 539481
rect 104806 539407 104862 539416
rect 103978 539064 104034 539073
rect 103978 538999 104034 539008
rect 104820 538558 104848 539407
rect 104808 538552 104860 538558
rect 104808 538494 104860 538500
rect 102966 527776 103022 527785
rect 102966 527711 103022 527720
rect 97908 527672 97960 527678
rect 97908 527614 97960 527620
rect 95608 526108 95660 526114
rect 95608 526050 95660 526056
rect 95620 520146 95648 526050
rect 97724 525020 97776 525026
rect 97724 524962 97776 524968
rect 96620 521144 96672 521150
rect 96620 521086 96672 521092
rect 96632 520146 96660 521086
rect 97736 520146 97764 524962
rect 97920 522510 97948 527614
rect 105004 526289 105032 560116
rect 106016 533905 106044 560116
rect 107028 540841 107056 560116
rect 107568 540864 107620 540870
rect 107014 540832 107070 540841
rect 107568 540806 107620 540812
rect 107014 540767 107070 540776
rect 107580 539889 107608 540806
rect 107566 539880 107622 539889
rect 107566 539815 107622 539824
rect 108040 535401 108068 560116
rect 109052 538214 109080 560116
rect 109052 538186 109264 538214
rect 109038 538112 109094 538121
rect 109038 538047 109094 538056
rect 109052 537198 109080 538047
rect 109040 537192 109092 537198
rect 109040 537134 109092 537140
rect 109040 536716 109092 536722
rect 109040 536658 109092 536664
rect 109052 535673 109080 536658
rect 109236 535945 109264 538186
rect 110064 537985 110092 560116
rect 111076 549273 111104 560116
rect 112088 551993 112116 560116
rect 112074 551984 112130 551993
rect 111800 551948 111852 551954
rect 112074 551919 112130 551928
rect 111800 551890 111852 551896
rect 111812 551313 111840 551890
rect 111798 551304 111854 551313
rect 111798 551239 111854 551248
rect 111062 549264 111118 549273
rect 111062 549199 111118 549208
rect 110420 549160 110472 549166
rect 110420 549102 110472 549108
rect 110432 548321 110460 549102
rect 110418 548312 110474 548321
rect 110418 548247 110474 548256
rect 110050 537976 110106 537985
rect 110050 537911 110106 537920
rect 109222 535936 109278 535945
rect 109222 535871 109278 535880
rect 109038 535664 109094 535673
rect 109038 535599 109094 535608
rect 108026 535392 108082 535401
rect 108026 535327 108082 535336
rect 108302 534848 108358 534857
rect 108302 534783 108358 534792
rect 108316 534410 108344 534783
rect 108304 534404 108356 534410
rect 108304 534346 108356 534352
rect 106188 534064 106240 534070
rect 106188 534006 106240 534012
rect 106002 533896 106058 533905
rect 106002 533831 106058 533840
rect 106200 533361 106228 534006
rect 106186 533352 106242 533361
rect 106186 533287 106242 533296
rect 105820 528624 105872 528630
rect 105820 528566 105872 528572
rect 104990 526280 105046 526289
rect 104990 526215 105046 526224
rect 101680 524816 101732 524822
rect 101680 524758 101732 524764
rect 99748 524748 99800 524754
rect 99748 524690 99800 524696
rect 98736 523320 98788 523326
rect 98736 523262 98788 523268
rect 97908 522504 97960 522510
rect 97908 522446 97960 522452
rect 98748 520146 98776 523262
rect 99760 520146 99788 524690
rect 100760 524612 100812 524618
rect 100760 524554 100812 524560
rect 100772 520146 100800 524554
rect 101692 520146 101720 524758
rect 102692 524680 102744 524686
rect 102692 524622 102744 524628
rect 102704 520146 102732 524622
rect 103796 523388 103848 523394
rect 103796 523330 103848 523336
rect 103808 520146 103836 523330
rect 104716 523252 104768 523258
rect 104716 523194 104768 523200
rect 104728 520146 104756 523194
rect 105832 520146 105860 528566
rect 113100 527105 113128 560116
rect 114112 552401 114140 560116
rect 114466 553344 114522 553353
rect 114466 553279 114522 553288
rect 114098 552392 114154 552401
rect 114098 552327 114154 552336
rect 114480 552158 114508 553279
rect 114468 552152 114520 552158
rect 114468 552094 114520 552100
rect 115124 534041 115152 560116
rect 116136 537169 116164 560116
rect 116122 537160 116178 537169
rect 116122 537095 116178 537104
rect 117148 535673 117176 560116
rect 117228 538144 117280 538150
rect 117228 538086 117280 538092
rect 117240 537033 117268 538086
rect 117226 537024 117282 537033
rect 117226 536959 117282 536968
rect 117228 536648 117280 536654
rect 117228 536590 117280 536596
rect 117240 535809 117268 536590
rect 117226 535800 117282 535809
rect 117226 535735 117282 535744
rect 117134 535664 117190 535673
rect 117134 535599 117190 535608
rect 115110 534032 115166 534041
rect 115110 533967 115166 533976
rect 115848 533996 115900 534002
rect 115848 533938 115900 533944
rect 115860 533089 115888 533938
rect 115846 533080 115902 533089
rect 115846 533015 115902 533024
rect 113086 527096 113142 527105
rect 111800 527060 111852 527066
rect 113086 527031 113142 527040
rect 111800 527002 111852 527008
rect 106186 526960 106242 526969
rect 106186 526895 106242 526904
rect 106200 526794 106228 526895
rect 106188 526788 106240 526794
rect 106188 526730 106240 526736
rect 111812 526561 111840 527002
rect 111798 526552 111854 526561
rect 111798 526487 111854 526496
rect 112904 526380 112956 526386
rect 112904 526322 112956 526328
rect 109776 526244 109828 526250
rect 109776 526186 109828 526192
rect 108764 526176 108816 526182
rect 108764 526118 108816 526124
rect 107844 522028 107896 522034
rect 107844 521970 107896 521976
rect 106832 520668 106884 520674
rect 106832 520610 106884 520616
rect 106844 520146 106872 520610
rect 107856 520146 107884 521970
rect 108776 520146 108804 526118
rect 109788 520146 109816 526186
rect 110788 526040 110840 526046
rect 110788 525982 110840 525988
rect 110800 520146 110828 525982
rect 111800 522572 111852 522578
rect 111800 522514 111852 522520
rect 111812 520146 111840 522514
rect 112916 520146 112944 526322
rect 114928 526312 114980 526318
rect 114928 526254 114980 526260
rect 113916 520532 113968 520538
rect 113916 520474 113968 520480
rect 113928 520146 113956 520474
rect 114940 520146 114968 526254
rect 116860 525972 116912 525978
rect 116860 525914 116912 525920
rect 115940 521824 115992 521830
rect 115940 521766 115992 521772
rect 115952 520146 115980 521766
rect 116872 520146 116900 525914
rect 117964 525564 118016 525570
rect 117964 525506 118016 525512
rect 117976 524793 118004 525506
rect 118160 524929 118188 560116
rect 119172 551857 119200 560116
rect 119158 551848 119214 551857
rect 118700 551812 118752 551818
rect 119158 551783 119214 551792
rect 118700 551754 118752 551760
rect 118712 551041 118740 551754
rect 118698 551032 118754 551041
rect 118698 550967 118754 550976
rect 120078 528048 120134 528057
rect 120078 527983 120134 527992
rect 120092 527882 120120 527983
rect 120184 527921 120212 560116
rect 121196 528057 121224 560116
rect 121460 528556 121512 528562
rect 121460 528498 121512 528504
rect 121182 528048 121238 528057
rect 121182 527983 121238 527992
rect 120170 527912 120226 527921
rect 120080 527876 120132 527882
rect 120170 527847 120226 527856
rect 120080 527818 120132 527824
rect 121472 527649 121500 528498
rect 122208 528465 122236 560116
rect 122194 528456 122250 528465
rect 122194 528391 122250 528400
rect 123220 528329 123248 560116
rect 124232 538214 124260 560116
rect 124864 539368 124916 539374
rect 124864 539310 124916 539316
rect 124232 538186 124628 538214
rect 123206 528320 123262 528329
rect 123206 528255 123262 528264
rect 124128 527672 124180 527678
rect 121458 527640 121514 527649
rect 124128 527614 124180 527620
rect 121458 527575 121514 527584
rect 123944 527604 123996 527610
rect 123944 527546 123996 527552
rect 122932 527332 122984 527338
rect 122932 527274 122984 527280
rect 120906 527232 120962 527241
rect 120962 527190 121040 527218
rect 120906 527167 120962 527176
rect 118146 524920 118202 524929
rect 118146 524855 118202 524864
rect 117962 524784 118018 524793
rect 117962 524719 118018 524728
rect 117872 523116 117924 523122
rect 117872 523058 117924 523064
rect 117884 520146 117912 523058
rect 118884 522436 118936 522442
rect 118884 522378 118936 522384
rect 118896 520146 118924 522378
rect 119896 520600 119948 520606
rect 119896 520542 119948 520548
rect 119908 520146 119936 520542
rect 121012 520146 121040 527190
rect 122012 524884 122064 524890
rect 122012 524826 122064 524832
rect 122024 520146 122052 524826
rect 122944 520146 122972 527274
rect 123956 520146 123984 527546
rect 124140 527377 124168 527614
rect 124600 527377 124628 538186
rect 124876 527950 124904 539310
rect 124864 527944 124916 527950
rect 124864 527886 124916 527892
rect 125244 527649 125272 560116
rect 126256 545465 126284 560116
rect 126888 546236 126940 546242
rect 126888 546178 126940 546184
rect 126242 545456 126298 545465
rect 126242 545391 126298 545400
rect 126900 545329 126928 546178
rect 126886 545320 126942 545329
rect 126886 545255 126942 545264
rect 127268 543561 127296 560116
rect 128280 557122 128308 560116
rect 128268 557116 128320 557122
rect 128268 557058 128320 557064
rect 128728 543720 128780 543726
rect 128728 543662 128780 543668
rect 127624 543652 127676 543658
rect 127624 543594 127676 543600
rect 127254 543552 127310 543561
rect 127254 543487 127310 543496
rect 127636 542881 127664 543594
rect 127622 542872 127678 542881
rect 127622 542807 127678 542816
rect 128360 542224 128412 542230
rect 128360 542166 128412 542172
rect 128372 541385 128400 542166
rect 128358 541376 128414 541385
rect 128358 541311 128414 541320
rect 128740 539374 128768 543662
rect 129292 541521 129320 560116
rect 129740 542156 129792 542162
rect 129740 542098 129792 542104
rect 129278 541512 129334 541521
rect 129278 541447 129334 541456
rect 129752 541249 129780 542098
rect 130304 541657 130332 560116
rect 131118 550624 131174 550633
rect 131118 550559 131174 550568
rect 131132 549438 131160 550559
rect 131316 550497 131344 560116
rect 131302 550488 131358 550497
rect 131302 550423 131358 550432
rect 131120 549432 131172 549438
rect 131120 549374 131172 549380
rect 131120 544944 131172 544950
rect 132328 544921 132356 560116
rect 131120 544886 131172 544892
rect 132314 544912 132370 544921
rect 131132 544105 131160 544886
rect 132314 544847 132370 544856
rect 131118 544096 131174 544105
rect 131118 544031 131174 544040
rect 130290 541648 130346 541657
rect 130290 541583 130346 541592
rect 129738 541240 129794 541249
rect 129738 541175 129794 541184
rect 128728 539368 128780 539374
rect 128728 539310 128780 539316
rect 125508 528488 125560 528494
rect 125508 528430 125560 528436
rect 125416 528352 125468 528358
rect 125416 528294 125468 528300
rect 125230 527640 125286 527649
rect 125230 527575 125286 527584
rect 125428 527513 125456 528294
rect 125520 528193 125548 528430
rect 133340 528222 133368 560116
rect 134536 543726 134564 591330
rect 135168 561672 135220 561678
rect 135168 561614 135220 561620
rect 135180 558210 135208 561614
rect 135168 558204 135220 558210
rect 135168 558146 135220 558152
rect 134524 543720 134576 543726
rect 134524 543662 134576 543668
rect 135166 530360 135222 530369
rect 135166 530295 135222 530304
rect 133328 528216 133380 528222
rect 125506 528184 125562 528193
rect 133328 528158 133380 528164
rect 125506 528119 125562 528128
rect 126980 527536 127032 527542
rect 125414 527504 125470 527513
rect 125048 527468 125100 527474
rect 126980 527478 127032 527484
rect 125414 527439 125470 527448
rect 125048 527410 125100 527416
rect 124126 527368 124182 527377
rect 124126 527303 124182 527312
rect 124586 527368 124642 527377
rect 124586 527303 124642 527312
rect 125060 520146 125088 527410
rect 125968 521960 126020 521966
rect 125968 521902 126020 521908
rect 125980 520146 126008 521902
rect 126992 520146 127020 527478
rect 132040 527400 132092 527406
rect 132040 527342 132092 527348
rect 130108 527196 130160 527202
rect 130108 527138 130160 527144
rect 129740 523524 129792 523530
rect 129740 523466 129792 523472
rect 129752 522442 129780 523466
rect 129740 522436 129792 522442
rect 129740 522378 129792 522384
rect 129096 521756 129148 521762
rect 129096 521698 129148 521704
rect 127992 520464 128044 520470
rect 127992 520406 128044 520412
rect 128004 520146 128032 520406
rect 129108 520146 129136 521698
rect 130120 520146 130148 527138
rect 131120 521892 131172 521898
rect 131120 521834 131172 521840
rect 131132 520146 131160 521834
rect 132052 520146 132080 527342
rect 133144 521008 133196 521014
rect 133144 520950 133196 520956
rect 133156 520146 133184 520950
rect 134064 520396 134116 520402
rect 134064 520338 134116 520344
rect 134076 520146 134104 520338
rect 135180 520146 135208 530295
rect 135916 526454 135944 700295
rect 137282 638752 137338 638761
rect 137204 638710 137282 638738
rect 135994 636984 136050 636993
rect 135994 636919 136050 636928
rect 136008 538665 136036 636919
rect 136178 636440 136234 636449
rect 136178 636375 136234 636384
rect 136088 602404 136140 602410
rect 136088 602346 136140 602352
rect 136100 591394 136128 602346
rect 136088 591388 136140 591394
rect 136088 591330 136140 591336
rect 136192 546961 136220 636375
rect 137204 634814 137232 638710
rect 137282 638687 137338 638696
rect 137284 638308 137336 638314
rect 137284 638250 137336 638256
rect 137296 638081 137324 638250
rect 137282 638072 137338 638081
rect 137282 638007 137338 638016
rect 137374 636712 137430 636721
rect 137374 636647 137430 636656
rect 137204 634786 137324 634814
rect 137296 620945 137324 634786
rect 137388 626249 137416 636647
rect 137374 626240 137430 626249
rect 137374 626175 137430 626184
rect 137282 620936 137338 620945
rect 137282 620871 137338 620880
rect 137466 618624 137522 618633
rect 137466 618559 137522 618568
rect 137282 611416 137338 611425
rect 137282 611351 137338 611360
rect 137190 575512 137246 575521
rect 137190 575447 137246 575456
rect 137098 572112 137154 572121
rect 137098 572047 137154 572056
rect 137112 555937 137140 572047
rect 137204 556170 137232 575447
rect 137192 556164 137244 556170
rect 137192 556106 137244 556112
rect 137192 556028 137244 556034
rect 137192 555970 137244 555976
rect 137098 555928 137154 555937
rect 137098 555863 137154 555872
rect 137204 554985 137232 555970
rect 137190 554976 137246 554985
rect 137190 554911 137246 554920
rect 136548 547732 136600 547738
rect 136548 547674 136600 547680
rect 136178 546952 136234 546961
rect 136178 546887 136234 546896
rect 136560 546689 136588 547674
rect 136546 546680 136602 546689
rect 136546 546615 136602 546624
rect 136548 539368 136600 539374
rect 136548 539310 136600 539316
rect 135994 538656 136050 538665
rect 135994 538591 136050 538600
rect 136560 538393 136588 539310
rect 136546 538384 136602 538393
rect 136546 538319 136602 538328
rect 137296 530602 137324 611351
rect 137374 606384 137430 606393
rect 137374 606319 137430 606328
rect 137388 531049 137416 606319
rect 137480 556306 137508 618559
rect 137650 608016 137706 608025
rect 137650 607951 137706 607960
rect 137558 604480 137614 604489
rect 137558 604415 137614 604424
rect 137468 556300 137520 556306
rect 137468 556242 137520 556248
rect 137468 556164 137520 556170
rect 137468 556106 137520 556112
rect 137480 555626 137508 556106
rect 137468 555620 137520 555626
rect 137468 555562 137520 555568
rect 137572 531321 137600 604415
rect 137664 555558 137692 607951
rect 137742 592512 137798 592521
rect 137742 592447 137798 592456
rect 137756 556986 137784 592447
rect 137744 556980 137796 556986
rect 137744 556922 137796 556928
rect 137744 556300 137796 556306
rect 137744 556242 137796 556248
rect 137652 555552 137704 555558
rect 137652 555494 137704 555500
rect 137756 550186 137784 556242
rect 137744 550180 137796 550186
rect 137744 550122 137796 550128
rect 137558 531312 137614 531321
rect 137558 531247 137614 531256
rect 137374 531040 137430 531049
rect 137374 530975 137430 530984
rect 137284 530596 137336 530602
rect 137284 530538 137336 530544
rect 137190 530496 137246 530505
rect 137190 530431 137246 530440
rect 136180 527264 136232 527270
rect 136180 527206 136232 527212
rect 135904 526448 135956 526454
rect 135904 526390 135956 526396
rect 136192 520146 136220 527206
rect 137204 520146 137232 530431
rect 137848 528426 137876 703520
rect 154132 700369 154160 703520
rect 163502 700496 163558 700505
rect 163502 700431 163558 700440
rect 154118 700360 154174 700369
rect 154118 700295 154174 700304
rect 163516 687177 163544 700431
rect 170324 700330 170352 703520
rect 202800 700505 202828 703520
rect 202786 700496 202842 700505
rect 202786 700431 202842 700440
rect 218992 700369 219020 703520
rect 235184 700369 235212 703520
rect 176934 700360 176990 700369
rect 170312 700324 170364 700330
rect 176934 700295 176990 700304
rect 218978 700360 219034 700369
rect 218978 700295 219034 700304
rect 235170 700360 235226 700369
rect 235170 700295 235226 700304
rect 170312 700266 170364 700272
rect 176948 698329 176976 700295
rect 173162 698320 173218 698329
rect 173162 698255 173218 698264
rect 176934 698320 176990 698329
rect 176934 698255 176990 698264
rect 173176 688537 173204 698255
rect 164422 688528 164478 688537
rect 164252 688486 164422 688514
rect 160098 687168 160154 687177
rect 160098 687103 160154 687112
rect 163502 687168 163558 687177
rect 163502 687103 163558 687112
rect 160112 685137 160140 687103
rect 164252 685930 164280 688486
rect 164422 688463 164478 688472
rect 173162 688528 173218 688537
rect 173162 688463 173218 688472
rect 267660 687954 267688 703520
rect 255964 687948 256016 687954
rect 255964 687890 256016 687896
rect 267648 687948 267700 687954
rect 267648 687890 267700 687896
rect 163700 685902 164280 685930
rect 158718 685128 158774 685137
rect 158718 685063 158774 685072
rect 160098 685128 160154 685137
rect 160098 685063 160154 685072
rect 158732 676274 158760 685063
rect 163700 677521 163728 685902
rect 162122 677512 162178 677521
rect 162122 677447 162178 677456
rect 163686 677512 163742 677521
rect 163686 677447 163742 677456
rect 158640 676246 158760 676274
rect 158640 674801 158668 676246
rect 153842 674792 153898 674801
rect 153842 674727 153898 674736
rect 158626 674792 158682 674801
rect 158626 674727 158682 674736
rect 153856 662561 153884 674727
rect 162136 667865 162164 677447
rect 255976 674830 256004 687890
rect 283852 687206 283880 703520
rect 300136 700398 300164 703520
rect 300124 700392 300176 700398
rect 300124 700334 300176 700340
rect 322204 700392 322256 700398
rect 322204 700334 322256 700340
rect 323582 700360 323638 700369
rect 283840 687200 283892 687206
rect 283840 687142 283892 687148
rect 286324 687200 286376 687206
rect 286324 687142 286376 687148
rect 250444 674824 250496 674830
rect 250444 674766 250496 674772
rect 255964 674824 256016 674830
rect 255964 674766 256016 674772
rect 158810 667856 158866 667865
rect 158810 667791 158866 667800
rect 162122 667856 162178 667865
rect 162122 667791 162178 667800
rect 158824 665825 158852 667791
rect 157338 665816 157394 665825
rect 157338 665751 157394 665760
rect 158810 665816 158866 665825
rect 158810 665751 158866 665760
rect 151082 662552 151138 662561
rect 151082 662487 151138 662496
rect 153842 662552 153898 662561
rect 153842 662487 153898 662496
rect 144184 657484 144236 657490
rect 144184 657426 144236 657432
rect 138664 644632 138716 644638
rect 138664 644574 138716 644580
rect 138676 637362 138704 644574
rect 138664 637356 138716 637362
rect 138664 637298 138716 637304
rect 142804 619608 142856 619614
rect 142804 619550 142856 619556
rect 141424 593360 141476 593366
rect 141424 593302 141476 593308
rect 137926 588432 137982 588441
rect 137926 588367 137982 588376
rect 137940 556918 137968 588367
rect 140044 583772 140096 583778
rect 140044 583714 140096 583720
rect 140056 561882 140084 583714
rect 140044 561876 140096 561882
rect 140044 561818 140096 561824
rect 141436 559570 141464 593302
rect 142816 586566 142844 619550
rect 142896 611380 142948 611386
rect 142896 611322 142948 611328
rect 142908 593366 142936 611322
rect 142896 593360 142948 593366
rect 142896 593302 142948 593308
rect 141516 586560 141568 586566
rect 141516 586502 141568 586508
rect 142804 586560 142856 586566
rect 142804 586502 142856 586508
rect 141528 583778 141556 586502
rect 141516 583772 141568 583778
rect 141516 583714 141568 583720
rect 141424 559564 141476 559570
rect 141424 559506 141476 559512
rect 137928 556912 137980 556918
rect 137928 556854 137980 556860
rect 144196 540258 144224 657426
rect 149702 649496 149758 649505
rect 149702 649431 149758 649440
rect 146208 645856 146260 645862
rect 146208 645798 146260 645804
rect 146220 641918 146248 645798
rect 144276 641912 144328 641918
rect 144276 641854 144328 641860
rect 146208 641912 146260 641918
rect 146208 641854 146260 641860
rect 144288 611386 144316 641854
rect 149716 640354 149744 649431
rect 151096 645930 151124 662487
rect 157352 657665 157380 665751
rect 250456 661774 250484 674766
rect 242440 661768 242492 661774
rect 242440 661710 242492 661716
rect 250444 661768 250496 661774
rect 250444 661710 250496 661716
rect 151174 657656 151230 657665
rect 151174 657591 151230 657600
rect 157338 657656 157394 657665
rect 157338 657591 157394 657600
rect 151188 649505 151216 657591
rect 242452 655518 242480 661710
rect 286336 657694 286364 687142
rect 322216 657762 322244 700334
rect 332520 700330 332548 703520
rect 323582 700295 323638 700304
rect 324964 700324 325016 700330
rect 322204 657756 322256 657762
rect 322204 657698 322256 657704
rect 286324 657688 286376 657694
rect 286324 657630 286376 657636
rect 294604 657688 294656 657694
rect 323596 657665 323624 700295
rect 324964 700266 325016 700272
rect 332508 700324 332560 700330
rect 332508 700266 332560 700272
rect 340144 700324 340196 700330
rect 340144 700266 340196 700272
rect 324976 657694 325004 700266
rect 340156 677550 340184 700266
rect 348804 686526 348832 703520
rect 348792 686520 348844 686526
rect 348792 686462 348844 686468
rect 358084 686520 358136 686526
rect 358084 686462 358136 686468
rect 358096 680406 358124 686462
rect 358084 680400 358136 680406
rect 358084 680342 358136 680348
rect 360844 680400 360896 680406
rect 360844 680342 360896 680348
rect 340144 677544 340196 677550
rect 340144 677486 340196 677492
rect 345664 677544 345716 677550
rect 345664 677486 345716 677492
rect 345676 660346 345704 677486
rect 360856 672110 360884 680342
rect 360844 672104 360896 672110
rect 360844 672046 360896 672052
rect 345664 660340 345716 660346
rect 345664 660282 345716 660288
rect 355968 660340 356020 660346
rect 355968 660282 356020 660288
rect 324964 657688 325016 657694
rect 294604 657630 294656 657636
rect 323582 657656 323638 657665
rect 239404 655512 239456 655518
rect 239404 655454 239456 655460
rect 242440 655512 242492 655518
rect 242440 655454 242492 655460
rect 178038 655072 178094 655081
rect 178038 655007 178094 655016
rect 177854 654936 177910 654945
rect 177854 654871 177910 654880
rect 177670 654800 177726 654809
rect 177670 654735 177726 654744
rect 156604 654560 156656 654566
rect 156604 654502 156656 654508
rect 151174 649496 151230 649505
rect 151174 649431 151230 649440
rect 151084 645924 151136 645930
rect 151084 645866 151136 645872
rect 153936 642252 153988 642258
rect 153936 642194 153988 642200
rect 148324 640348 148376 640354
rect 148324 640290 148376 640296
rect 149704 640348 149756 640354
rect 149704 640290 149756 640296
rect 148336 630698 148364 640290
rect 153842 639840 153898 639849
rect 153842 639775 153898 639784
rect 151084 634500 151136 634506
rect 151084 634442 151136 634448
rect 146944 630692 146996 630698
rect 146944 630634 146996 630640
rect 148324 630692 148376 630698
rect 148324 630634 148376 630640
rect 146956 621042 146984 630634
rect 144920 621036 144972 621042
rect 144920 620978 144972 620984
rect 146944 621036 146996 621042
rect 146944 620978 146996 620984
rect 144932 619614 144960 620978
rect 144920 619608 144972 619614
rect 144920 619550 144972 619556
rect 144276 611380 144328 611386
rect 144276 611322 144328 611328
rect 151096 547806 151124 634442
rect 151360 554804 151412 554810
rect 151360 554746 151412 554752
rect 151084 547800 151136 547806
rect 151084 547742 151136 547748
rect 148324 541068 148376 541074
rect 148324 541010 148376 541016
rect 144184 540252 144236 540258
rect 144184 540194 144236 540200
rect 138204 530188 138256 530194
rect 138204 530130 138256 530136
rect 137836 528420 137888 528426
rect 137836 528362 137888 528368
rect 138216 520146 138244 530130
rect 140228 530120 140280 530126
rect 140228 530062 140280 530068
rect 139400 523184 139452 523190
rect 139400 523126 139452 523132
rect 139412 522306 139440 523126
rect 139216 522300 139268 522306
rect 139216 522242 139268 522248
rect 139400 522300 139452 522306
rect 139400 522242 139452 522248
rect 139228 520146 139256 522242
rect 140240 520146 140268 530062
rect 147312 530052 147364 530058
rect 147312 529994 147364 530000
rect 144276 529984 144328 529990
rect 144276 529926 144328 529932
rect 143264 525904 143316 525910
rect 143264 525846 143316 525852
rect 142160 522436 142212 522442
rect 142160 522378 142212 522384
rect 141148 520940 141200 520946
rect 141148 520882 141200 520888
rect 141160 520146 141188 520882
rect 142172 520690 142200 522378
rect 142172 520662 142292 520690
rect 142264 520146 142292 520662
rect 143276 520146 143304 525846
rect 144288 520146 144316 529926
rect 144828 524544 144880 524550
rect 144828 524486 144880 524492
rect 144840 521966 144868 524486
rect 144828 521960 144880 521966
rect 144828 521902 144880 521908
rect 145472 521756 145524 521762
rect 145472 521698 145524 521704
rect 145484 520146 145512 521698
rect 146484 521076 146536 521082
rect 146484 521018 146536 521024
rect 146496 520146 146524 521018
rect 88628 520118 88672 520146
rect 89640 520118 89684 520146
rect 90652 520118 90696 520146
rect 91664 520118 91708 520146
rect 92676 520118 92720 520146
rect 93688 520118 93732 520146
rect 94700 520118 94744 520146
rect 95620 520118 95756 520146
rect 96632 520118 96768 520146
rect 97736 520118 97780 520146
rect 98748 520118 98792 520146
rect 99760 520118 99804 520146
rect 100772 520118 100816 520146
rect 101692 520118 101828 520146
rect 102704 520118 102840 520146
rect 103808 520118 103852 520146
rect 104728 520118 104864 520146
rect 105832 520118 105876 520146
rect 106844 520118 106888 520146
rect 107856 520118 107900 520146
rect 108776 520118 108912 520146
rect 109788 520118 109924 520146
rect 110800 520118 110936 520146
rect 111812 520118 111948 520146
rect 112916 520118 112960 520146
rect 113928 520118 113972 520146
rect 114940 520118 114984 520146
rect 115952 520118 115996 520146
rect 116872 520118 117008 520146
rect 117884 520118 118020 520146
rect 118896 520118 119032 520146
rect 119908 520118 120044 520146
rect 121012 520118 121056 520146
rect 122024 520118 122068 520146
rect 122944 520118 123080 520146
rect 123956 520118 124092 520146
rect 125060 520118 125104 520146
rect 125980 520118 126116 520146
rect 126992 520118 127128 520146
rect 128004 520118 128140 520146
rect 129108 520118 129152 520146
rect 130120 520118 130164 520146
rect 131132 520118 131176 520146
rect 132052 520118 132188 520146
rect 133156 520118 133200 520146
rect 134076 520118 134212 520146
rect 135180 520118 135224 520146
rect 136192 520118 136236 520146
rect 137204 520118 137248 520146
rect 138216 520118 138260 520146
rect 139228 520118 139272 520146
rect 140240 520118 140284 520146
rect 141160 520118 141296 520146
rect 142264 520118 142308 520146
rect 143276 520118 143320 520146
rect 144288 520118 144332 520146
rect 86620 519860 86648 520118
rect 87632 519860 87660 520118
rect 88644 519860 88672 520118
rect 89656 519860 89684 520118
rect 90668 519860 90696 520118
rect 91680 519860 91708 520118
rect 92692 519860 92720 520118
rect 93704 519860 93732 520118
rect 94716 519860 94744 520118
rect 95728 519860 95756 520118
rect 96740 519860 96768 520118
rect 97752 519860 97780 520118
rect 98764 519860 98792 520118
rect 99776 519860 99804 520118
rect 100788 519860 100816 520118
rect 101800 519860 101828 520118
rect 102812 519860 102840 520118
rect 103824 519860 103852 520118
rect 104836 519860 104864 520118
rect 105848 519860 105876 520118
rect 106860 519860 106888 520118
rect 107872 519860 107900 520118
rect 108884 519860 108912 520118
rect 109896 519860 109924 520118
rect 110908 519860 110936 520118
rect 111920 519860 111948 520118
rect 112932 519860 112960 520118
rect 113944 519860 113972 520118
rect 114956 519860 114984 520118
rect 115968 519860 115996 520118
rect 116980 519860 117008 520118
rect 117992 519860 118020 520118
rect 119004 519860 119032 520118
rect 120016 519860 120044 520118
rect 121028 519860 121056 520118
rect 122040 519860 122068 520118
rect 123052 519860 123080 520118
rect 124064 519860 124092 520118
rect 125076 519860 125104 520118
rect 126088 519860 126116 520118
rect 127100 519860 127128 520118
rect 128112 519860 128140 520118
rect 129124 519860 129152 520118
rect 130136 519860 130164 520118
rect 131148 519860 131176 520118
rect 132160 519860 132188 520118
rect 133172 519860 133200 520118
rect 134184 519860 134212 520118
rect 135196 519860 135224 520118
rect 136208 519860 136236 520118
rect 137220 519860 137248 520118
rect 138232 519860 138260 520118
rect 139244 519860 139272 520118
rect 140256 519860 140284 520118
rect 141268 519860 141296 520118
rect 142280 519860 142308 520118
rect 143292 519860 143320 520118
rect 144304 519860 144332 520118
rect 145316 520118 145512 520146
rect 146328 520118 146524 520146
rect 147324 520146 147352 529994
rect 148336 520146 148364 541010
rect 150348 522436 150400 522442
rect 150348 522378 150400 522384
rect 149244 521960 149296 521966
rect 149244 521902 149296 521908
rect 149256 520146 149284 521902
rect 150360 520146 150388 522378
rect 151372 520146 151400 554746
rect 153856 530641 153884 639775
rect 153948 550458 153976 642194
rect 154486 639976 154542 639985
rect 154486 639911 154542 639920
rect 154500 639402 154528 639911
rect 154488 639396 154540 639402
rect 154488 639338 154540 639344
rect 156616 557462 156644 654502
rect 176568 647352 176620 647358
rect 176566 647320 176568 647329
rect 176620 647320 176622 647329
rect 176566 647255 176622 647264
rect 176566 645960 176622 645969
rect 176566 645895 176568 645904
rect 176620 645895 176622 645904
rect 176568 645866 176620 645872
rect 177304 644836 177356 644842
rect 177304 644778 177356 644784
rect 176752 643544 176804 643550
rect 176752 643486 176804 643492
rect 176660 643408 176712 643414
rect 176660 643350 176712 643356
rect 176672 637430 176700 643350
rect 176764 637566 176792 643486
rect 176752 637560 176804 637566
rect 176752 637502 176804 637508
rect 177316 637498 177344 644778
rect 177580 640552 177632 640558
rect 177580 640494 177632 640500
rect 177592 640393 177620 640494
rect 177578 640384 177634 640393
rect 177578 640319 177634 640328
rect 177304 637492 177356 637498
rect 177304 637434 177356 637440
rect 176660 637424 176712 637430
rect 176660 637366 176712 637372
rect 175094 637256 175150 637265
rect 175094 637191 175150 637200
rect 173898 635624 173954 635633
rect 173898 635559 173954 635568
rect 156696 635520 156748 635526
rect 156696 635462 156748 635468
rect 156604 557456 156656 557462
rect 156604 557398 156656 557404
rect 156708 553110 156736 635462
rect 171968 634432 172020 634438
rect 171968 634374 172020 634380
rect 166354 626512 166410 626521
rect 166354 626447 166410 626456
rect 166262 623248 166318 623257
rect 166262 623183 166318 623192
rect 159364 613420 159416 613426
rect 159364 613362 159416 613368
rect 159376 602410 159404 613362
rect 164882 607744 164938 607753
rect 164882 607679 164938 607688
rect 163594 603664 163650 603673
rect 163594 603599 163650 603608
rect 159364 602404 159416 602410
rect 159364 602346 159416 602352
rect 162398 595232 162454 595241
rect 162398 595167 162454 595176
rect 162122 594688 162178 594697
rect 162122 594623 162178 594632
rect 159362 581632 159418 581641
rect 159362 581567 159418 581576
rect 156696 553104 156748 553110
rect 156696 553046 156748 553052
rect 153936 550452 153988 550458
rect 153936 550394 153988 550400
rect 158444 539708 158496 539714
rect 158444 539650 158496 539656
rect 156420 538416 156472 538422
rect 156420 538358 156472 538364
rect 154396 534200 154448 534206
rect 154396 534142 154448 534148
rect 153842 530632 153898 530641
rect 153842 530567 153898 530576
rect 152556 526176 152608 526182
rect 152556 526118 152608 526124
rect 152568 520146 152596 526118
rect 153384 522504 153436 522510
rect 153384 522446 153436 522452
rect 147324 520118 147368 520146
rect 148336 520118 148380 520146
rect 149256 520118 149392 520146
rect 150360 520118 150404 520146
rect 151372 520118 151416 520146
rect 145316 519860 145344 520118
rect 146328 519860 146356 520118
rect 147340 519860 147368 520118
rect 148352 519860 148380 520118
rect 149364 519860 149392 520118
rect 150376 519860 150404 520118
rect 151388 519860 151416 520118
rect 152400 520118 152596 520146
rect 153396 520146 153424 522446
rect 154408 520146 154436 534142
rect 155408 528624 155460 528630
rect 155408 528566 155460 528572
rect 155420 520146 155448 528566
rect 156432 520146 156460 538358
rect 157984 534132 158036 534138
rect 157984 534074 158036 534080
rect 157996 528358 158024 534074
rect 157984 528352 158036 528358
rect 157984 528294 158036 528300
rect 157340 522300 157392 522306
rect 157340 522242 157392 522248
rect 157352 520146 157380 522242
rect 158456 520146 158484 539650
rect 159376 527950 159404 581567
rect 159546 581224 159602 581233
rect 159546 581159 159602 581168
rect 159454 579728 159510 579737
rect 159454 579663 159510 579672
rect 159468 555257 159496 579663
rect 159454 555248 159510 555257
rect 159454 555183 159510 555192
rect 159560 552537 159588 581159
rect 159730 581088 159786 581097
rect 159730 581023 159786 581032
rect 159638 578504 159694 578513
rect 159638 578439 159694 578448
rect 159652 555529 159680 578439
rect 159744 556753 159772 581023
rect 159730 556744 159786 556753
rect 159730 556679 159786 556688
rect 159638 555520 159694 555529
rect 159638 555455 159694 555464
rect 159546 552528 159602 552537
rect 159546 552463 159602 552472
rect 161480 548004 161532 548010
rect 161480 547946 161532 547952
rect 160744 543312 160796 543318
rect 160744 543254 160796 543260
rect 160756 534138 160784 543254
rect 160744 534132 160796 534138
rect 160744 534074 160796 534080
rect 159364 527944 159416 527950
rect 159364 527886 159416 527892
rect 159640 525156 159692 525162
rect 159640 525098 159692 525104
rect 159652 520146 159680 525098
rect 160560 521824 160612 521830
rect 160560 521766 160612 521772
rect 160572 520146 160600 521766
rect 153396 520118 153440 520146
rect 154408 520118 154452 520146
rect 155420 520118 155464 520146
rect 156432 520118 156476 520146
rect 157352 520118 157488 520146
rect 158456 520118 158500 520146
rect 152400 519860 152428 520118
rect 153412 519860 153440 520118
rect 154424 519860 154452 520118
rect 155436 519860 155464 520118
rect 156448 519860 156476 520118
rect 157460 519860 157488 520118
rect 158472 519860 158500 520118
rect 159484 520118 159680 520146
rect 160496 520118 160600 520146
rect 161492 520146 161520 547946
rect 162136 530641 162164 594623
rect 162308 586628 162360 586634
rect 162308 586570 162360 586576
rect 162214 571840 162270 571849
rect 162214 571775 162270 571784
rect 162122 530632 162178 530641
rect 162122 530567 162178 530576
rect 162228 528154 162256 571775
rect 162320 559881 162348 586570
rect 162412 560561 162440 595167
rect 162490 592104 162546 592113
rect 162490 592039 162546 592048
rect 162398 560552 162454 560561
rect 162398 560487 162454 560496
rect 162504 560250 162532 592039
rect 163502 591424 163558 591433
rect 163502 591359 163558 591368
rect 162584 586560 162636 586566
rect 162584 586502 162636 586508
rect 162492 560244 162544 560250
rect 162492 560186 162544 560192
rect 162306 559872 162362 559881
rect 162306 559807 162362 559816
rect 162596 558657 162624 586502
rect 162766 576872 162822 576881
rect 162766 576807 162822 576816
rect 162674 576600 162730 576609
rect 162674 576535 162730 576544
rect 162582 558648 162638 558657
rect 162582 558583 162638 558592
rect 162688 555801 162716 576535
rect 162780 557025 162808 576807
rect 162766 557016 162822 557025
rect 162766 556951 162822 556960
rect 163516 556481 163544 591359
rect 163502 556472 163558 556481
rect 163502 556407 163558 556416
rect 162674 555792 162730 555801
rect 162674 555727 162730 555736
rect 162490 554840 162546 554849
rect 162490 554775 162546 554784
rect 162216 528148 162268 528154
rect 162216 528090 162268 528096
rect 162504 520146 162532 554775
rect 163504 550656 163556 550662
rect 163504 550598 163556 550604
rect 163516 520146 163544 550598
rect 163608 531185 163636 603599
rect 164896 555257 164924 607679
rect 164974 589656 165030 589665
rect 164974 589591 165030 589600
rect 164988 569702 165016 589591
rect 165158 588024 165214 588033
rect 165158 587959 165214 587968
rect 165068 579828 165120 579834
rect 165068 579770 165120 579776
rect 165080 569945 165108 579770
rect 165172 576854 165200 587959
rect 165172 576826 165292 576854
rect 165066 569936 165122 569945
rect 165066 569871 165122 569880
rect 164976 569696 165028 569702
rect 164976 569638 165028 569644
rect 164988 557433 165016 569638
rect 164974 557424 165030 557433
rect 164974 557359 165030 557368
rect 165080 555665 165108 569871
rect 165264 556617 165292 576826
rect 166170 569392 166226 569401
rect 166170 569327 166226 569336
rect 165528 560108 165580 560114
rect 165528 560050 165580 560056
rect 165250 556608 165306 556617
rect 165250 556543 165306 556552
rect 165540 556322 165568 560050
rect 166184 559609 166212 569327
rect 166170 559600 166226 559609
rect 166170 559535 166226 559544
rect 165448 556294 165568 556322
rect 165448 556073 165476 556294
rect 165526 556200 165582 556209
rect 165526 556135 165582 556144
rect 165434 556064 165490 556073
rect 165434 555999 165490 556008
rect 165066 555656 165122 555665
rect 165066 555591 165122 555600
rect 164882 555248 164938 555257
rect 164882 555183 164938 555192
rect 163594 531176 163650 531185
rect 163594 531111 163650 531120
rect 164146 531040 164202 531049
rect 164146 530975 164202 530984
rect 164160 530534 164188 530975
rect 164148 530528 164200 530534
rect 164148 530470 164200 530476
rect 164700 520464 164752 520470
rect 164700 520406 164752 520412
rect 164712 520146 164740 520406
rect 161492 520118 161536 520146
rect 162504 520118 162548 520146
rect 163516 520118 163560 520146
rect 159484 519860 159512 520118
rect 160496 519860 160524 520118
rect 161508 519860 161536 520118
rect 162520 519860 162548 520118
rect 163532 519860 163560 520118
rect 164544 520118 164740 520146
rect 165540 520146 165568 556135
rect 166172 547800 166224 547806
rect 166172 547742 166224 547748
rect 166184 546553 166212 547742
rect 166170 546544 166226 546553
rect 166170 546479 166226 546488
rect 166172 531276 166224 531282
rect 166172 531218 166224 531224
rect 166184 530233 166212 531218
rect 166170 530224 166226 530233
rect 166170 530159 166226 530168
rect 166276 528554 166304 623183
rect 166368 548554 166396 626447
rect 169022 624880 169078 624889
rect 169022 624815 169078 624824
rect 167642 624064 167698 624073
rect 167642 623999 167698 624008
rect 166446 605296 166502 605305
rect 166446 605231 166502 605240
rect 166356 548548 166408 548554
rect 166356 548490 166408 548496
rect 166460 530913 166488 605231
rect 166630 590608 166686 590617
rect 166630 590543 166686 590552
rect 166540 559020 166592 559026
rect 166540 558962 166592 558968
rect 166446 530904 166502 530913
rect 166446 530839 166502 530848
rect 166276 528526 166488 528554
rect 166460 521529 166488 528526
rect 166446 521520 166502 521529
rect 166264 521484 166316 521490
rect 166446 521455 166502 521464
rect 166264 521426 166316 521432
rect 166276 520713 166304 521426
rect 166262 520704 166318 520713
rect 166262 520639 166318 520648
rect 166552 520146 166580 558962
rect 166644 556617 166672 590543
rect 166906 582176 166962 582185
rect 166906 582111 166962 582120
rect 166920 581233 166948 582111
rect 166906 581224 166962 581233
rect 166906 581159 166962 581168
rect 166814 560280 166870 560289
rect 166814 560215 166870 560224
rect 166828 558958 166856 560215
rect 166816 558952 166868 558958
rect 166816 558894 166868 558900
rect 166630 556608 166686 556617
rect 166630 556543 166686 556552
rect 166920 547874 166948 581159
rect 166828 547846 166948 547874
rect 166828 546825 166856 547846
rect 166814 546816 166870 546825
rect 166814 546751 166870 546760
rect 166906 537568 166962 537577
rect 166906 537503 166962 537512
rect 166920 536926 166948 537503
rect 166908 536920 166960 536926
rect 166908 536862 166960 536868
rect 167552 534132 167604 534138
rect 167552 534074 167604 534080
rect 167092 521620 167144 521626
rect 167092 521562 167144 521568
rect 167000 521416 167052 521422
rect 167000 521358 167052 521364
rect 167012 521121 167040 521358
rect 166998 521112 167054 521121
rect 166998 521047 167054 521056
rect 167104 520849 167132 521562
rect 167090 520840 167146 520849
rect 167090 520775 167146 520784
rect 167564 520146 167592 534074
rect 167656 521665 167684 623999
rect 167826 622432 167882 622441
rect 167826 622367 167882 622376
rect 167734 589792 167790 589801
rect 167734 589727 167790 589736
rect 167748 557025 167776 589727
rect 167734 557016 167790 557025
rect 167734 556951 167790 556960
rect 167642 521656 167698 521665
rect 167642 521591 167698 521600
rect 167840 521393 167868 622367
rect 168286 585304 168342 585313
rect 168286 585239 168342 585248
rect 168102 585168 168158 585177
rect 168102 585103 168158 585112
rect 168012 560244 168064 560250
rect 168012 560186 168064 560192
rect 168024 557161 168052 560186
rect 168116 557297 168144 585103
rect 168300 558521 168328 585239
rect 168286 558512 168342 558521
rect 168286 558447 168342 558456
rect 168102 557288 168158 557297
rect 168102 557223 168158 557232
rect 168010 557152 168066 557161
rect 168010 557087 168066 557096
rect 168380 550384 168432 550390
rect 168380 550326 168432 550332
rect 168392 549545 168420 550326
rect 168378 549536 168434 549545
rect 168378 549471 168434 549480
rect 168380 536580 168432 536586
rect 168380 536522 168432 536528
rect 168392 535537 168420 536522
rect 168378 535528 168434 535537
rect 168378 535463 168434 535472
rect 168564 531480 168616 531486
rect 168564 531422 168616 531428
rect 168380 521552 168432 521558
rect 168380 521494 168432 521500
rect 167826 521384 167882 521393
rect 167826 521319 167882 521328
rect 168392 520577 168420 521494
rect 168378 520568 168434 520577
rect 168378 520503 168434 520512
rect 168576 520146 168604 531422
rect 169036 520849 169064 624815
rect 171782 619984 171838 619993
rect 171782 619919 171838 619928
rect 170494 600400 170550 600409
rect 170494 600335 170550 600344
rect 170402 598768 170458 598777
rect 170402 598703 170458 598712
rect 169390 591968 169446 591977
rect 169390 591903 169446 591912
rect 169114 573472 169170 573481
rect 169114 573407 169170 573416
rect 169128 562358 169156 573407
rect 169300 569832 169352 569838
rect 169220 569792 169300 569820
rect 169116 562352 169168 562358
rect 169116 562294 169168 562300
rect 169220 560386 169248 569792
rect 169300 569774 169352 569780
rect 169404 567194 169432 591903
rect 169574 590880 169630 590889
rect 169574 590815 169630 590824
rect 169484 586560 169536 586566
rect 169588 586514 169616 590815
rect 170310 588160 170366 588169
rect 170310 588095 170366 588104
rect 169536 586508 169616 586514
rect 169484 586502 169616 586508
rect 169496 586486 169616 586502
rect 169482 581088 169538 581097
rect 169482 581023 169538 581032
rect 169312 567166 169432 567194
rect 169208 560380 169260 560386
rect 169208 560322 169260 560328
rect 169220 556889 169248 560322
rect 169312 559858 169340 567166
rect 169390 559872 169446 559881
rect 169312 559830 169390 559858
rect 169390 559807 169446 559816
rect 169206 556880 169262 556889
rect 169206 556815 169262 556824
rect 169496 550633 169524 581023
rect 169588 558249 169616 586486
rect 169942 578504 169998 578513
rect 169942 578439 169998 578448
rect 169666 577824 169722 577833
rect 169666 577759 169722 577768
rect 169680 576881 169708 577759
rect 169666 576872 169722 576881
rect 169666 576807 169722 576816
rect 169574 558240 169630 558249
rect 169574 558175 169630 558184
rect 169482 550624 169538 550633
rect 169482 550559 169538 550568
rect 169680 536625 169708 576807
rect 169850 559736 169906 559745
rect 169850 559671 169906 559680
rect 169864 559502 169892 559671
rect 169852 559496 169904 559502
rect 169758 559464 169814 559473
rect 169852 559438 169904 559444
rect 169758 559399 169760 559408
rect 169812 559399 169814 559408
rect 169760 559370 169812 559376
rect 169760 549024 169812 549030
rect 169760 548966 169812 548972
rect 169772 548185 169800 548966
rect 169956 548321 169984 578439
rect 170128 562352 170180 562358
rect 170128 562294 170180 562300
rect 170140 557534 170168 562294
rect 170048 557506 170168 557534
rect 170048 555393 170076 557506
rect 170324 556345 170352 588095
rect 170310 556336 170366 556345
rect 170310 556271 170366 556280
rect 170034 555384 170090 555393
rect 170034 555319 170090 555328
rect 170048 552537 170076 555319
rect 170034 552528 170090 552537
rect 170034 552463 170090 552472
rect 169942 548312 169998 548321
rect 169942 548247 169998 548256
rect 169758 548176 169814 548185
rect 169758 548111 169814 548120
rect 169760 544876 169812 544882
rect 169760 544818 169812 544824
rect 169772 543969 169800 544818
rect 169758 543960 169814 543969
rect 169758 543895 169814 543904
rect 169760 540728 169812 540734
rect 169760 540670 169812 540676
rect 169772 539753 169800 540670
rect 169758 539744 169814 539753
rect 169758 539679 169814 539688
rect 169666 536616 169722 536625
rect 169666 536551 169722 536560
rect 169760 535356 169812 535362
rect 169760 535298 169812 535304
rect 169772 534313 169800 535298
rect 170416 534721 170444 598703
rect 170508 540569 170536 600335
rect 170586 599584 170642 599593
rect 170586 599519 170642 599528
rect 170600 544610 170628 599519
rect 170770 597952 170826 597961
rect 170770 597887 170826 597896
rect 170678 592240 170734 592249
rect 170678 592175 170734 592184
rect 170692 544649 170720 592175
rect 170784 552838 170812 597887
rect 171046 596864 171102 596873
rect 171046 596799 171102 596808
rect 170862 594144 170918 594153
rect 170862 594079 170918 594088
rect 170876 586634 170904 594079
rect 170864 586628 170916 586634
rect 170864 586570 170916 586576
rect 170876 586514 170904 586570
rect 170876 586486 170996 586514
rect 170968 559745 170996 586486
rect 171060 560017 171088 596799
rect 171138 574560 171194 574569
rect 171138 574495 171194 574504
rect 171152 569838 171180 574495
rect 171140 569832 171192 569838
rect 171140 569774 171192 569780
rect 171046 560008 171102 560017
rect 171046 559943 171102 559952
rect 170954 559736 171010 559745
rect 170954 559671 171010 559680
rect 170864 557048 170916 557054
rect 170864 556990 170916 556996
rect 170772 552832 170824 552838
rect 170772 552774 170824 552780
rect 170678 544640 170734 544649
rect 170588 544604 170640 544610
rect 170678 544575 170734 544584
rect 170588 544546 170640 544552
rect 170494 540560 170550 540569
rect 170494 540495 170550 540504
rect 170588 538348 170640 538354
rect 170588 538290 170640 538296
rect 170402 534712 170458 534721
rect 170402 534647 170458 534656
rect 169758 534304 169814 534313
rect 169758 534239 169814 534248
rect 169576 532840 169628 532846
rect 169576 532782 169628 532788
rect 169022 520840 169078 520849
rect 169022 520775 169078 520784
rect 169588 520146 169616 532782
rect 170600 520146 170628 538290
rect 170876 522306 170904 556990
rect 171796 536178 171824 619919
rect 171874 615088 171930 615097
rect 171874 615023 171930 615032
rect 171784 536172 171836 536178
rect 171784 536114 171836 536120
rect 171888 533526 171916 615023
rect 171980 613426 172008 634374
rect 173254 615904 173310 615913
rect 173254 615839 173310 615848
rect 171968 613420 172020 613426
rect 171968 613362 172020 613368
rect 173162 612640 173218 612649
rect 173162 612575 173218 612584
rect 171966 602032 172022 602041
rect 171966 601967 172022 601976
rect 171980 541822 172008 601967
rect 172058 601216 172114 601225
rect 172058 601151 172114 601160
rect 172072 547330 172100 601151
rect 172426 586392 172482 586401
rect 172426 586327 172482 586336
rect 172150 583264 172206 583273
rect 172150 583199 172206 583208
rect 172164 559337 172192 583199
rect 172440 576854 172468 586327
rect 172978 579728 173034 579737
rect 172978 579663 173034 579672
rect 172348 576826 172468 576854
rect 172244 560380 172296 560386
rect 172244 560322 172296 560328
rect 172150 559328 172206 559337
rect 172150 559263 172206 559272
rect 172256 551313 172284 560322
rect 172348 560250 172376 576826
rect 172428 569696 172480 569702
rect 172428 569638 172480 569644
rect 172336 560244 172388 560250
rect 172336 560186 172388 560192
rect 172348 555529 172376 560186
rect 172440 557161 172468 569638
rect 172886 561640 172942 561649
rect 172886 561575 172942 561584
rect 172426 557152 172482 557161
rect 172426 557087 172482 557096
rect 172334 555520 172390 555529
rect 172334 555455 172390 555464
rect 172428 551880 172480 551886
rect 172428 551822 172480 551828
rect 172242 551304 172298 551313
rect 172242 551239 172298 551248
rect 172440 550769 172468 551822
rect 172426 550760 172482 550769
rect 172426 550695 172482 550704
rect 172060 547324 172112 547330
rect 172060 547266 172112 547272
rect 172612 542496 172664 542502
rect 172612 542438 172664 542444
rect 171968 541816 172020 541822
rect 171968 541758 172020 541764
rect 172426 541784 172482 541793
rect 172426 541719 172482 541728
rect 172440 541210 172468 541719
rect 172428 541204 172480 541210
rect 172428 541146 172480 541152
rect 171876 533520 171928 533526
rect 171876 533462 171928 533468
rect 171692 523048 171744 523054
rect 171692 522990 171744 522996
rect 170864 522300 170916 522306
rect 170864 522242 170916 522248
rect 171704 520146 171732 522990
rect 165540 520118 165584 520146
rect 166552 520118 166596 520146
rect 167564 520118 167608 520146
rect 168576 520118 168620 520146
rect 169588 520118 169632 520146
rect 170600 520118 170644 520146
rect 164544 519860 164572 520118
rect 165556 519860 165584 520118
rect 166568 519860 166596 520118
rect 167580 519860 167608 520118
rect 168592 519860 168620 520118
rect 169604 519860 169632 520118
rect 170616 519860 170644 520118
rect 171628 520118 171732 520146
rect 172624 520146 172652 542438
rect 172900 537538 172928 561575
rect 172992 560561 173020 579663
rect 173070 575104 173126 575113
rect 173070 575039 173126 575048
rect 172978 560552 173034 560561
rect 172978 560487 173034 560496
rect 172978 559328 173034 559337
rect 172978 559263 173034 559272
rect 172992 558657 173020 559263
rect 172978 558648 173034 558657
rect 172978 558583 173034 558592
rect 173084 554985 173112 575039
rect 173070 554976 173126 554985
rect 173070 554911 173126 554920
rect 172888 537532 172940 537538
rect 172888 537474 172940 537480
rect 173176 529378 173204 612575
rect 173268 543114 173296 615839
rect 173438 614272 173494 614281
rect 173438 614207 173494 614216
rect 173346 602848 173402 602857
rect 173346 602783 173402 602792
rect 173256 543108 173308 543114
rect 173256 543050 173308 543056
rect 173360 530505 173388 602783
rect 173452 545970 173480 614207
rect 173912 596873 173940 635559
rect 174726 634808 174782 634817
rect 174726 634743 174782 634752
rect 174634 613456 174690 613465
rect 174634 613391 174690 613400
rect 174542 611008 174598 611017
rect 174542 610943 174598 610952
rect 173898 596864 173954 596873
rect 173898 596799 173954 596808
rect 173714 587616 173770 587625
rect 173714 587551 173770 587560
rect 173530 587344 173586 587353
rect 173530 587279 173586 587288
rect 173544 557433 173572 587279
rect 173728 579834 173756 587551
rect 173716 579828 173768 579834
rect 173716 579770 173768 579776
rect 173714 575648 173770 575657
rect 173714 575583 173770 575592
rect 173728 560114 173756 575583
rect 174450 574288 174506 574297
rect 174450 574223 174506 574232
rect 173806 569936 173862 569945
rect 173806 569871 173862 569880
rect 173716 560108 173768 560114
rect 173716 560050 173768 560056
rect 173728 557534 173756 560050
rect 173636 557506 173756 557534
rect 173530 557424 173586 557433
rect 173530 557359 173586 557368
rect 173636 549658 173664 557506
rect 173820 556050 173848 569871
rect 174266 558920 174322 558929
rect 174266 558855 174322 558864
rect 173728 556022 173848 556050
rect 173728 554577 173756 556022
rect 173808 554600 173860 554606
rect 173714 554568 173770 554577
rect 173808 554542 173860 554548
rect 173714 554503 173770 554512
rect 173820 553897 173848 554542
rect 173806 553888 173862 553897
rect 173806 553823 173862 553832
rect 174280 551410 174308 558855
rect 174464 555393 174492 574223
rect 174450 555384 174506 555393
rect 174450 555319 174506 555328
rect 174268 551404 174320 551410
rect 174268 551346 174320 551352
rect 173808 550452 173860 550458
rect 173808 550394 173860 550400
rect 173714 549672 173770 549681
rect 173636 549630 173714 549658
rect 173714 549607 173770 549616
rect 173820 549409 173848 550394
rect 173806 549400 173862 549409
rect 173806 549335 173862 549344
rect 173440 545964 173492 545970
rect 173440 545906 173492 545912
rect 174556 538898 174584 610943
rect 174648 554130 174676 613391
rect 174740 598505 174768 634743
rect 175108 615494 175136 637191
rect 176658 636848 176714 636857
rect 176658 636783 176714 636792
rect 176672 635769 176700 636783
rect 176658 635760 176714 635769
rect 176658 635695 176714 635704
rect 175186 634672 175242 634681
rect 175186 634607 175242 634616
rect 175200 633593 175228 634607
rect 175186 633584 175242 633593
rect 175186 633519 175242 633528
rect 177684 626793 177712 654735
rect 177762 636984 177818 636993
rect 177762 636919 177818 636928
rect 177776 630057 177804 636919
rect 177762 630048 177818 630057
rect 177762 629983 177818 629992
rect 177868 627881 177896 654871
rect 178052 654158 178080 655007
rect 178040 654152 178092 654158
rect 178040 654094 178092 654100
rect 189170 653576 189226 653585
rect 189170 653511 189226 653520
rect 184018 652352 184074 652361
rect 184018 652287 184074 652296
rect 178682 642560 178738 642569
rect 178682 642495 178738 642504
rect 178040 642320 178092 642326
rect 178040 642262 178092 642268
rect 178052 642161 178080 642262
rect 178038 642152 178094 642161
rect 178038 642087 178094 642096
rect 177948 642048 178000 642054
rect 177948 641990 178000 641996
rect 177960 641753 177988 641990
rect 177946 641744 178002 641753
rect 177946 641679 178002 641688
rect 177946 640384 178002 640393
rect 177946 640319 177948 640328
rect 178000 640319 178002 640328
rect 177948 640290 178000 640296
rect 177854 627872 177910 627881
rect 177854 627807 177910 627816
rect 177670 626784 177726 626793
rect 177670 626719 177726 626728
rect 177578 623520 177634 623529
rect 177578 623455 177634 623464
rect 175108 615466 175228 615494
rect 175200 610706 175228 615466
rect 177026 611416 177082 611425
rect 177026 611351 177082 611360
rect 175188 610700 175240 610706
rect 175188 610642 175240 610648
rect 175922 610192 175978 610201
rect 175922 610127 175978 610136
rect 174726 598496 174782 598505
rect 174726 598431 174782 598440
rect 174818 597136 174874 597145
rect 174818 597071 174874 597080
rect 174726 593872 174782 593881
rect 174726 593807 174782 593816
rect 174636 554124 174688 554130
rect 174636 554066 174688 554072
rect 174544 538892 174596 538898
rect 174544 538834 174596 538840
rect 174740 536246 174768 593807
rect 174832 548457 174860 597071
rect 174910 585712 174966 585721
rect 174910 585647 174966 585656
rect 174924 576858 174952 585647
rect 175186 585304 175242 585313
rect 175186 585239 175242 585248
rect 175094 585168 175150 585177
rect 175094 585103 175150 585112
rect 175108 582570 175136 585103
rect 175200 584361 175228 585239
rect 175830 584896 175886 584905
rect 175830 584831 175886 584840
rect 175186 584352 175242 584361
rect 175186 584287 175242 584296
rect 175108 582542 175228 582570
rect 174924 576830 175136 576858
rect 174910 572384 174966 572393
rect 174910 572319 174966 572328
rect 174924 558521 174952 572319
rect 175002 570208 175058 570217
rect 175002 570143 175058 570152
rect 174910 558512 174966 558521
rect 174910 558447 174966 558456
rect 174912 557116 174964 557122
rect 174912 557058 174964 557064
rect 174818 548448 174874 548457
rect 174818 548383 174874 548392
rect 174728 536240 174780 536246
rect 174728 536182 174780 536188
rect 173806 530904 173862 530913
rect 173806 530839 173862 530848
rect 173346 530496 173402 530505
rect 173346 530431 173402 530440
rect 173820 530194 173848 530839
rect 173808 530188 173860 530194
rect 173808 530130 173860 530136
rect 173164 529372 173216 529378
rect 173164 529314 173216 529320
rect 174636 528692 174688 528698
rect 174636 528634 174688 528640
rect 173808 525904 173860 525910
rect 173808 525846 173860 525852
rect 173820 520146 173848 525846
rect 172624 520118 172668 520146
rect 171628 519860 171656 520118
rect 172640 519860 172668 520118
rect 173652 520118 173848 520146
rect 174648 520146 174676 528634
rect 174924 522510 174952 557058
rect 175016 540682 175044 570143
rect 175108 556753 175136 576830
rect 175200 558385 175228 582542
rect 175554 571024 175610 571033
rect 175554 570959 175610 570968
rect 175462 560280 175518 560289
rect 175462 560215 175518 560224
rect 175186 558376 175242 558385
rect 175186 558311 175242 558320
rect 175094 556744 175150 556753
rect 175094 556679 175150 556688
rect 175188 556232 175240 556238
rect 175186 556200 175188 556209
rect 175240 556200 175242 556209
rect 175186 556135 175242 556144
rect 175188 548956 175240 548962
rect 175188 548898 175240 548904
rect 175200 547913 175228 548898
rect 175186 547904 175242 547913
rect 175186 547839 175242 547848
rect 175186 547224 175242 547233
rect 175186 547159 175242 547168
rect 175200 546582 175228 547159
rect 175188 546576 175240 546582
rect 175188 546518 175240 546524
rect 175016 540654 175320 540682
rect 175186 540560 175242 540569
rect 175292 540546 175320 540654
rect 175370 540560 175426 540569
rect 175292 540518 175370 540546
rect 175186 540495 175242 540504
rect 175370 540495 175426 540504
rect 175200 539850 175228 540495
rect 175188 539844 175240 539850
rect 175188 539786 175240 539792
rect 175476 532166 175504 560215
rect 175568 533497 175596 570959
rect 175740 560244 175792 560250
rect 175740 560186 175792 560192
rect 175752 559065 175780 560186
rect 175738 559056 175794 559065
rect 175738 558991 175794 559000
rect 175844 556889 175872 584831
rect 175830 556880 175886 556889
rect 175830 556815 175886 556824
rect 175830 556472 175886 556481
rect 175830 556407 175886 556416
rect 175844 556306 175872 556407
rect 175832 556300 175884 556306
rect 175832 556242 175884 556248
rect 175832 555484 175884 555490
rect 175832 555426 175884 555432
rect 175844 554849 175872 555426
rect 175830 554840 175886 554849
rect 175830 554775 175886 554784
rect 175832 551744 175884 551750
rect 175832 551686 175884 551692
rect 175844 550905 175872 551686
rect 175830 550896 175886 550905
rect 175830 550831 175886 550840
rect 175648 546644 175700 546650
rect 175648 546586 175700 546592
rect 175554 533488 175610 533497
rect 175554 533423 175610 533432
rect 175464 532160 175516 532166
rect 175464 532102 175516 532108
rect 174912 522504 174964 522510
rect 174912 522446 174964 522452
rect 175660 520146 175688 546586
rect 175936 537606 175964 610127
rect 176014 606112 176070 606121
rect 176014 606047 176070 606056
rect 176028 556073 176056 606047
rect 176290 595504 176346 595513
rect 176290 595439 176346 595448
rect 176198 583128 176254 583137
rect 176198 583063 176254 583072
rect 176106 579864 176162 579873
rect 176106 579799 176162 579808
rect 176014 556064 176070 556073
rect 176014 555999 176070 556008
rect 175924 537600 175976 537606
rect 175924 537542 175976 537548
rect 175922 536208 175978 536217
rect 175922 536143 175978 536152
rect 175936 535770 175964 536143
rect 175924 535764 175976 535770
rect 175924 535706 175976 535712
rect 175924 533928 175976 533934
rect 175924 533870 175976 533876
rect 175936 532953 175964 533870
rect 175922 532944 175978 532953
rect 175922 532879 175978 532888
rect 175922 531312 175978 531321
rect 175922 531247 175978 531256
rect 175936 530466 175964 531247
rect 176120 530913 176148 579799
rect 176212 536081 176240 583063
rect 176304 555801 176332 595439
rect 176566 588704 176622 588713
rect 176566 588639 176622 588648
rect 176580 588033 176608 588639
rect 176566 588024 176622 588033
rect 176566 587959 176622 587968
rect 176382 584352 176438 584361
rect 176382 584287 176438 584296
rect 176396 559337 176424 584287
rect 176474 582584 176530 582593
rect 176474 582519 176530 582528
rect 176382 559328 176438 559337
rect 176382 559263 176438 559272
rect 176290 555792 176346 555801
rect 176290 555727 176346 555736
rect 176488 551041 176516 582519
rect 176580 559473 176608 587959
rect 176566 559464 176622 559473
rect 176566 559399 176622 559408
rect 176474 551032 176530 551041
rect 176474 550967 176530 550976
rect 176566 549808 176622 549817
rect 176566 549743 176622 549752
rect 176580 549302 176608 549743
rect 176568 549296 176620 549302
rect 176568 549238 176620 549244
rect 176198 536072 176254 536081
rect 176198 536007 176254 536016
rect 176106 530904 176162 530913
rect 176106 530839 176162 530848
rect 175924 530460 175976 530466
rect 175924 530402 175976 530408
rect 177040 529310 177068 611351
rect 177302 609784 177358 609793
rect 177302 609719 177358 609728
rect 177210 607200 177266 607209
rect 177210 607135 177266 607144
rect 177118 569936 177174 569945
rect 177118 569871 177174 569880
rect 177132 533390 177160 569871
rect 177224 559570 177252 607135
rect 177212 559564 177264 559570
rect 177212 559506 177264 559512
rect 177316 558278 177344 609719
rect 177394 608560 177450 608569
rect 177394 608495 177450 608504
rect 177304 558272 177356 558278
rect 177304 558214 177356 558220
rect 177408 549914 177436 608495
rect 177486 601760 177542 601769
rect 177486 601695 177542 601704
rect 177396 549908 177448 549914
rect 177396 549850 177448 549856
rect 177500 544406 177528 601695
rect 177592 558210 177620 623455
rect 178696 621625 178724 642495
rect 183100 641912 183152 641918
rect 183100 641854 183152 641860
rect 179142 638480 179198 638489
rect 179142 638415 179198 638424
rect 179052 637900 179104 637906
rect 179052 637842 179104 637848
rect 179064 637673 179092 637842
rect 179050 637664 179106 637673
rect 179050 637599 179106 637608
rect 178958 635624 179014 635633
rect 178958 635559 179014 635568
rect 178774 633720 178830 633729
rect 178774 633655 178830 633664
rect 178682 621616 178738 621625
rect 178682 621551 178738 621560
rect 177854 610736 177910 610745
rect 177854 610671 177910 610680
rect 177670 607064 177726 607073
rect 177670 606999 177726 607008
rect 177580 558204 177632 558210
rect 177580 558146 177632 558152
rect 177488 544400 177540 544406
rect 177488 544342 177540 544348
rect 177684 540326 177712 606999
rect 177762 604480 177818 604489
rect 177762 604415 177818 604424
rect 177672 540320 177724 540326
rect 177672 540262 177724 540268
rect 177776 534750 177804 604415
rect 177764 534744 177816 534750
rect 177764 534686 177816 534692
rect 177120 533384 177172 533390
rect 177120 533326 177172 533332
rect 177868 529922 177896 610671
rect 178038 593056 178094 593065
rect 178038 592991 178094 593000
rect 178052 592113 178080 592991
rect 178038 592104 178094 592113
rect 178038 592039 178094 592048
rect 178590 584080 178646 584089
rect 178590 584015 178646 584024
rect 178498 573336 178554 573345
rect 178498 573271 178554 573280
rect 178406 568576 178462 568585
rect 178406 568511 178462 568520
rect 178420 562358 178448 568511
rect 178408 562352 178460 562358
rect 178408 562294 178460 562300
rect 178130 557016 178186 557025
rect 178130 556951 178186 556960
rect 178038 556608 178094 556617
rect 178038 556543 178094 556552
rect 178052 556374 178080 556543
rect 178144 556442 178172 556951
rect 178132 556436 178184 556442
rect 178132 556378 178184 556384
rect 178040 556368 178092 556374
rect 178040 556310 178092 556316
rect 178512 555665 178540 573271
rect 178604 557025 178632 584015
rect 178684 562352 178736 562358
rect 178684 562294 178736 562300
rect 178590 557016 178646 557025
rect 178590 556951 178646 556960
rect 178498 555656 178554 555665
rect 178498 555591 178554 555600
rect 178038 555248 178094 555257
rect 178038 555183 178094 555192
rect 178052 555014 178080 555183
rect 178040 555008 178092 555014
rect 178040 554950 178092 554956
rect 177946 554704 178002 554713
rect 177946 554639 178002 554648
rect 177960 553450 177988 554639
rect 178040 554532 178092 554538
rect 178040 554474 178092 554480
rect 178052 554169 178080 554474
rect 178038 554160 178094 554169
rect 178038 554095 178094 554104
rect 177948 553444 178000 553450
rect 177948 553386 178000 553392
rect 178040 549092 178092 549098
rect 178040 549034 178092 549040
rect 178052 548049 178080 549034
rect 178696 548865 178724 562294
rect 178682 548856 178738 548865
rect 178682 548791 178738 548800
rect 178038 548040 178094 548049
rect 178038 547975 178094 547984
rect 178040 542292 178092 542298
rect 178040 542234 178092 542240
rect 178052 541113 178080 542234
rect 178684 541136 178736 541142
rect 178038 541104 178094 541113
rect 178684 541078 178736 541084
rect 178038 541039 178094 541048
rect 177946 532672 178002 532681
rect 177946 532607 178002 532616
rect 177960 531418 177988 532607
rect 177948 531412 178000 531418
rect 177948 531354 178000 531360
rect 178224 531208 178276 531214
rect 178038 531176 178094 531185
rect 178224 531150 178276 531156
rect 178038 531111 178094 531120
rect 178132 531140 178184 531146
rect 178052 530262 178080 531111
rect 178132 531082 178184 531088
rect 178040 530256 178092 530262
rect 178040 530198 178092 530204
rect 178144 529961 178172 531082
rect 178236 530097 178264 531150
rect 178222 530088 178278 530097
rect 178222 530023 178278 530032
rect 178130 529952 178186 529961
rect 177856 529916 177908 529922
rect 178130 529887 178186 529896
rect 177856 529858 177908 529864
rect 177028 529304 177080 529310
rect 177028 529246 177080 529252
rect 177764 527264 177816 527270
rect 177764 527206 177816 527212
rect 176844 526448 176896 526454
rect 176844 526390 176896 526396
rect 176856 520146 176884 526390
rect 177776 520146 177804 527206
rect 178040 526992 178092 526998
rect 178040 526934 178092 526940
rect 178052 526425 178080 526934
rect 178038 526416 178094 526425
rect 178038 526351 178094 526360
rect 177946 525736 178002 525745
rect 177946 525671 178002 525680
rect 177960 524550 177988 525671
rect 177948 524544 178000 524550
rect 177948 524486 178000 524492
rect 177948 523524 178000 523530
rect 177948 523466 178000 523472
rect 177960 523433 177988 523466
rect 177946 523424 178002 523433
rect 177946 523359 178002 523368
rect 178040 522980 178092 522986
rect 178040 522922 178092 522928
rect 178052 522617 178080 522922
rect 178038 522608 178094 522617
rect 178038 522543 178094 522552
rect 174648 520118 174692 520146
rect 175660 520118 175704 520146
rect 173652 519860 173680 520118
rect 174664 519860 174692 520118
rect 175676 519860 175704 520118
rect 176688 520118 176884 520146
rect 177700 520118 177804 520146
rect 178696 520146 178724 541078
rect 178788 530890 178816 633655
rect 178972 600681 179000 635559
rect 179156 634817 179184 638415
rect 179326 636440 179382 636449
rect 179326 636375 179328 636384
rect 179380 636375 179382 636384
rect 179328 636346 179380 636352
rect 179972 636268 180024 636274
rect 179972 636210 180024 636216
rect 179234 635488 179290 635497
rect 179234 635423 179290 635432
rect 179142 634808 179198 634817
rect 179142 634743 179198 634752
rect 179142 633584 179198 633593
rect 179142 633519 179198 633528
rect 179052 610700 179104 610706
rect 179052 610642 179104 610648
rect 179064 601769 179092 610642
rect 179050 601760 179106 601769
rect 179050 601695 179106 601704
rect 178958 600672 179014 600681
rect 178958 600607 179014 600616
rect 179156 599593 179184 633519
rect 179142 599584 179198 599593
rect 179142 599519 179198 599528
rect 179248 597417 179276 635423
rect 179984 633457 180012 636210
rect 183112 634930 183140 641854
rect 184032 635202 184060 652287
rect 185306 652080 185362 652089
rect 185306 652015 185362 652024
rect 185320 635202 185348 652015
rect 187882 651400 187938 651409
rect 187882 651335 187938 651344
rect 186318 650448 186374 650457
rect 186318 650383 186374 650392
rect 186332 650078 186360 650383
rect 186594 650176 186650 650185
rect 186594 650111 186650 650120
rect 186320 650072 186372 650078
rect 186320 650014 186372 650020
rect 185674 635624 185730 635633
rect 185412 635582 185674 635610
rect 185412 635497 185440 635582
rect 185674 635559 185730 635568
rect 185398 635488 185454 635497
rect 185398 635423 185454 635432
rect 186608 635202 186636 650111
rect 186964 643748 187016 643754
rect 186964 643690 187016 643696
rect 182712 634902 183140 634930
rect 183986 635174 184060 635202
rect 185274 635174 185348 635202
rect 186562 635174 186636 635202
rect 183986 634916 184014 635174
rect 185274 634916 185302 635174
rect 186562 634916 186590 635174
rect 186976 634438 187004 643690
rect 187896 635202 187924 651335
rect 189184 635202 189212 653511
rect 190458 653440 190514 653449
rect 190458 653375 190514 653384
rect 190472 635202 190500 653375
rect 194322 653304 194378 653313
rect 194322 653239 194378 653248
rect 193128 640416 193180 640422
rect 193128 640358 193180 640364
rect 191746 637120 191802 637129
rect 187850 635174 187924 635202
rect 189138 635174 189212 635202
rect 190426 635174 190500 635202
rect 191668 637078 191746 637106
rect 191668 635202 191696 637078
rect 191746 637055 191802 637064
rect 191746 636848 191802 636857
rect 191746 636783 191802 636792
rect 191760 636342 191788 636783
rect 191748 636336 191800 636342
rect 191748 636278 191800 636284
rect 191668 635174 191742 635202
rect 187850 634916 187878 635174
rect 189138 634916 189166 635174
rect 190426 634916 190454 635174
rect 191714 634916 191742 635174
rect 193140 634930 193168 640358
rect 194336 635202 194364 653239
rect 227718 652352 227774 652361
rect 227718 652287 227774 652296
rect 211066 651944 211122 651953
rect 211066 651879 211122 651888
rect 208490 651808 208546 651817
rect 208490 651743 208546 651752
rect 207202 651536 207258 651545
rect 207202 651471 207258 651480
rect 205914 649768 205970 649777
rect 205914 649703 205970 649712
rect 205640 648848 205692 648854
rect 205640 648790 205692 648796
rect 199660 648712 199712 648718
rect 196898 648680 196954 648689
rect 196898 648615 196954 648624
rect 198738 648680 198794 648689
rect 205652 648689 205680 648790
rect 199660 648654 199712 648660
rect 200762 648680 200818 648689
rect 198738 648615 198740 648624
rect 195888 640688 195940 640694
rect 195888 640630 195940 640636
rect 193016 634902 193168 634930
rect 194290 635174 194364 635202
rect 194290 634916 194318 635174
rect 195900 634930 195928 640630
rect 196912 635202 196940 648615
rect 198792 648615 198794 648624
rect 198740 648586 198792 648592
rect 199672 644474 199700 648654
rect 200762 648615 200818 648624
rect 205638 648680 205694 648689
rect 205638 648615 205694 648624
rect 199488 644446 199700 644474
rect 198464 643136 198516 643142
rect 198464 643078 198516 643084
rect 195592 634902 195928 634930
rect 196866 635174 196940 635202
rect 196866 634916 196894 635174
rect 198476 634930 198504 643078
rect 199488 635202 199516 644446
rect 200776 635202 200804 648615
rect 203340 647420 203392 647426
rect 203340 647362 203392 647368
rect 202420 642116 202472 642122
rect 202420 642058 202472 642064
rect 198168 634902 198504 634930
rect 199442 635174 199516 635202
rect 200730 635174 200804 635202
rect 199442 634916 199470 635174
rect 200730 634916 200758 635174
rect 202432 634930 202460 642058
rect 203352 635202 203380 647362
rect 204628 645992 204680 645998
rect 204628 645934 204680 645940
rect 204640 635202 204668 645934
rect 205928 635202 205956 649703
rect 207216 635202 207244 651471
rect 208504 635202 208532 651743
rect 209780 646060 209832 646066
rect 209780 646002 209832 646008
rect 209792 635202 209820 646002
rect 211080 635202 211108 651879
rect 213826 651672 213882 651681
rect 214102 651672 214158 651681
rect 213826 651607 213882 651616
rect 213932 651630 214102 651658
rect 213840 651574 213868 651607
rect 213828 651568 213880 651574
rect 213828 651510 213880 651516
rect 213932 651386 213960 651630
rect 214102 651607 214158 651616
rect 227732 651438 227760 652287
rect 227810 652216 227866 652225
rect 227810 652151 227866 652160
rect 232976 652174 233372 652202
rect 213656 651358 213960 651386
rect 227720 651432 227772 651438
rect 227720 651374 227772 651380
rect 212446 650720 212502 650729
rect 212446 650655 212502 650664
rect 212354 650448 212410 650457
rect 212354 650383 212410 650392
rect 212368 635202 212396 650383
rect 212460 650146 212488 650655
rect 212448 650140 212500 650146
rect 212448 650082 212500 650088
rect 213656 635202 213684 651358
rect 226338 651128 226394 651137
rect 226338 651063 226394 651072
rect 214562 650992 214618 651001
rect 214562 650927 214618 650936
rect 214576 650214 214604 650927
rect 214930 650720 214986 650729
rect 214930 650655 214986 650664
rect 214564 650208 214616 650214
rect 214564 650150 214616 650156
rect 214944 635202 214972 650655
rect 226352 650282 226380 651063
rect 226522 650856 226578 650865
rect 226522 650791 226578 650800
rect 226340 650276 226392 650282
rect 226340 650218 226392 650224
rect 224222 649768 224278 649777
rect 224222 649703 224278 649712
rect 223946 649496 224002 649505
rect 223946 649431 224002 649440
rect 217508 647488 217560 647494
rect 217508 647430 217560 647436
rect 216588 642184 216640 642190
rect 216588 642126 216640 642132
rect 202032 634902 202460 634930
rect 203306 635174 203380 635202
rect 204594 635174 204668 635202
rect 205882 635174 205956 635202
rect 207170 635174 207244 635202
rect 208458 635174 208532 635202
rect 209746 635174 209820 635202
rect 211034 635174 211108 635202
rect 212322 635174 212396 635202
rect 213610 635174 213684 635202
rect 214898 635174 214972 635202
rect 203306 634916 203334 635174
rect 204594 634916 204622 635174
rect 205882 634916 205910 635174
rect 207170 634916 207198 635174
rect 208458 634916 208486 635174
rect 209746 634916 209774 635174
rect 211034 634916 211062 635174
rect 212322 634916 212350 635174
rect 213610 634916 213638 635174
rect 214898 634916 214926 635174
rect 216600 634930 216628 642126
rect 217520 635202 217548 647430
rect 218796 644768 218848 644774
rect 218796 644710 218848 644716
rect 218808 635202 218836 644710
rect 221740 643272 221792 643278
rect 221740 643214 221792 643220
rect 220360 639464 220412 639470
rect 220360 639406 220412 639412
rect 216200 634902 216628 634930
rect 217474 635174 217548 635202
rect 218762 635174 218836 635202
rect 217474 634916 217502 635174
rect 218762 634916 218790 635174
rect 220372 634930 220400 639406
rect 221752 634930 221780 643214
rect 222936 640756 222988 640762
rect 222936 640698 222988 640704
rect 222948 634930 222976 640698
rect 223960 635202 223988 649431
rect 224236 648786 224264 649703
rect 224224 648780 224276 648786
rect 224224 648722 224276 648728
rect 225512 643204 225564 643210
rect 225512 643146 225564 643152
rect 220064 634902 220400 634930
rect 221352 634902 221780 634930
rect 222640 634902 222976 634930
rect 223914 635174 223988 635202
rect 223914 634916 223942 635174
rect 225524 634930 225552 643146
rect 226536 635202 226564 650791
rect 227718 638888 227774 638897
rect 227718 638823 227774 638832
rect 227732 638246 227760 638823
rect 227720 638240 227772 638246
rect 227720 638182 227772 638188
rect 227824 635202 227852 652151
rect 231766 650584 231822 650593
rect 232042 650584 232098 650593
rect 231766 650519 231822 650528
rect 231872 650542 232042 650570
rect 231780 650350 231808 650519
rect 231768 650344 231820 650350
rect 231768 650286 231820 650292
rect 231872 650162 231900 650542
rect 232042 650519 232098 650528
rect 231688 650134 231900 650162
rect 230388 644700 230440 644706
rect 230388 644642 230440 644648
rect 227902 638344 227958 638353
rect 227902 638279 227958 638288
rect 227916 637537 227944 638279
rect 227902 637528 227958 637537
rect 227902 637463 227958 637472
rect 229466 636848 229522 636857
rect 229466 636783 229522 636792
rect 225216 634902 225552 634930
rect 226490 635174 226564 635202
rect 227778 635174 227852 635202
rect 226490 634916 226518 635174
rect 227778 634916 227806 635174
rect 229480 634930 229508 636783
rect 230400 635202 230428 644642
rect 231688 635202 231716 650134
rect 232976 635202 233004 652174
rect 233146 652080 233202 652089
rect 233344 652066 233372 652174
rect 233422 652080 233478 652089
rect 233344 652038 233422 652066
rect 233146 652015 233202 652024
rect 233422 652015 233478 652024
rect 233160 651506 233188 652015
rect 233148 651500 233200 651506
rect 233148 651442 233200 651448
rect 234618 648136 234674 648145
rect 234618 648071 234674 648080
rect 235538 648136 235594 648145
rect 235538 648071 235594 648080
rect 234632 647562 234660 648071
rect 234620 647556 234672 647562
rect 234620 647498 234672 647504
rect 234528 638376 234580 638382
rect 234528 638318 234580 638324
rect 229080 634902 229508 634930
rect 230354 635174 230428 635202
rect 231642 635174 231716 635202
rect 232930 635174 233004 635202
rect 230354 634916 230382 635174
rect 231642 634916 231670 635174
rect 232930 634916 232958 635174
rect 234540 634930 234568 638318
rect 235552 635202 235580 648071
rect 239416 643754 239444 655454
rect 294616 646542 294644 657630
rect 324964 657630 325016 657636
rect 323582 657591 323638 657600
rect 355980 654838 356008 660282
rect 364996 657830 365024 703520
rect 366364 672104 366416 672110
rect 366364 672046 366416 672052
rect 364984 657824 365036 657830
rect 364984 657766 365036 657772
rect 366376 656878 366404 672046
rect 366364 656872 366416 656878
rect 366364 656814 366416 656820
rect 371884 656872 371936 656878
rect 371884 656814 371936 656820
rect 355968 654832 356020 654838
rect 355968 654774 356020 654780
rect 366364 654832 366416 654838
rect 366364 654774 366416 654780
rect 359370 654664 359426 654673
rect 359370 654599 359426 654608
rect 356794 654528 356850 654537
rect 356794 654463 356850 654472
rect 305274 653712 305330 653721
rect 305274 653647 305330 653656
rect 294604 646536 294656 646542
rect 294604 646478 294656 646484
rect 304264 646536 304316 646542
rect 304264 646478 304316 646484
rect 240692 646128 240744 646134
rect 240692 646070 240744 646076
rect 239404 643748 239456 643754
rect 239404 643690 239456 643696
rect 237286 637392 237342 637401
rect 237208 637350 237286 637378
rect 235998 636984 236054 636993
rect 235998 636919 236054 636928
rect 236012 636614 236040 636919
rect 236000 636608 236052 636614
rect 236000 636550 236052 636556
rect 234232 634902 234568 634930
rect 235506 635174 235580 635202
rect 235506 634916 235534 635174
rect 237208 634930 237236 637350
rect 237286 637327 237342 637336
rect 240046 637120 240102 637129
rect 240046 637055 240102 637064
rect 237378 636576 237434 636585
rect 237378 636511 237434 636520
rect 239678 636576 239734 636585
rect 239678 636511 239734 636520
rect 236808 634902 237236 634930
rect 237392 634681 237420 636511
rect 238390 636440 238446 636449
rect 238390 636375 238446 636384
rect 238404 634930 238432 636375
rect 239692 634930 239720 636511
rect 240060 636478 240088 637055
rect 240048 636472 240100 636478
rect 240048 636414 240100 636420
rect 240704 635202 240732 646070
rect 261666 644056 261722 644065
rect 261666 643991 261722 644000
rect 259642 643920 259698 643929
rect 259642 643855 259698 643864
rect 251086 641336 251142 641345
rect 251086 641271 251142 641280
rect 249706 641064 249762 641073
rect 249706 640999 249762 641008
rect 249720 640898 249748 640999
rect 251100 640966 251128 641271
rect 259366 641064 259422 641073
rect 259366 640999 259422 641008
rect 251088 640960 251140 640966
rect 251088 640902 251140 640908
rect 249708 640892 249760 640898
rect 249708 640834 249760 640840
rect 249706 640384 249762 640393
rect 249706 640319 249762 640328
rect 242806 637392 242862 637401
rect 242806 637327 242862 637336
rect 242438 636984 242494 636993
rect 238096 634902 238432 634930
rect 239384 634902 239720 634930
rect 240658 635174 240732 635202
rect 242360 636942 242438 636970
rect 240658 634916 240686 635174
rect 242360 634930 242388 636942
rect 242438 636919 242494 636928
rect 242820 636682 242848 637327
rect 245014 637120 245070 637129
rect 244936 637078 245014 637106
rect 242808 636676 242860 636682
rect 242808 636618 242860 636624
rect 244936 634930 244964 637078
rect 245014 637055 245070 637064
rect 247130 637120 247186 637129
rect 247130 637055 247186 637064
rect 245568 636744 245620 636750
rect 245568 636686 245620 636692
rect 245580 636449 245608 636686
rect 247144 636585 247172 637055
rect 246946 636576 247002 636585
rect 246946 636511 246948 636520
rect 247000 636511 247002 636520
rect 247130 636576 247186 636585
rect 247130 636511 247186 636520
rect 246948 636482 247000 636488
rect 245566 636440 245622 636449
rect 245566 636375 245622 636384
rect 246118 636440 246174 636449
rect 246118 636375 246174 636384
rect 246132 634930 246160 636375
rect 249720 636313 249748 640319
rect 258722 638480 258778 638489
rect 258722 638415 258778 638424
rect 250902 638344 250958 638353
rect 258078 638344 258134 638353
rect 250958 638302 251036 638330
rect 250902 638279 250958 638288
rect 249706 636304 249762 636313
rect 249706 636239 249762 636248
rect 247592 635452 247644 635458
rect 247592 635394 247644 635400
rect 247604 634930 247632 635394
rect 249720 635202 249748 636239
rect 251008 635202 251036 638302
rect 258078 638279 258134 638288
rect 256606 638208 256662 638217
rect 252468 638172 252520 638178
rect 256606 638143 256662 638152
rect 252468 638114 252520 638120
rect 241960 634902 242388 634930
rect 244536 634902 244964 634930
rect 245824 634902 246160 634930
rect 247112 634902 247632 634930
rect 249674 635174 249748 635202
rect 250962 635174 251036 635202
rect 249674 634916 249702 635174
rect 250962 634916 250990 635174
rect 252480 634930 252508 638114
rect 255594 635760 255650 635769
rect 255594 635695 255650 635704
rect 252264 634902 252508 634930
rect 248372 634808 248428 634817
rect 248372 634743 248428 634752
rect 237378 634672 237434 634681
rect 237378 634607 237434 634616
rect 186964 634432 187016 634438
rect 186964 634374 187016 634380
rect 243211 634208 243220 634264
rect 243276 634208 243285 634264
rect 179970 633448 180026 633457
rect 179970 633383 180026 633392
rect 179234 597408 179290 597417
rect 179234 597343 179290 597352
rect 179970 594960 180026 594969
rect 179970 594895 180026 594904
rect 179050 593056 179106 593065
rect 179050 592991 179106 593000
rect 178866 580816 178922 580825
rect 178866 580751 178922 580760
rect 178880 531010 178908 580751
rect 178958 578368 179014 578377
rect 178958 578303 179014 578312
rect 178972 531049 179000 578303
rect 179064 560318 179092 592991
rect 179234 579184 179290 579193
rect 179234 579119 179290 579128
rect 179142 577552 179198 577561
rect 179142 577487 179198 577496
rect 179052 560312 179104 560318
rect 179052 560254 179104 560260
rect 179050 560144 179106 560153
rect 179050 560079 179106 560088
rect 179064 554198 179092 560079
rect 179052 554192 179104 554198
rect 179052 554134 179104 554140
rect 179156 531185 179184 577487
rect 179248 541793 179276 579119
rect 179326 576736 179382 576745
rect 179326 576671 179382 576680
rect 179878 576736 179934 576745
rect 179878 576671 179934 576680
rect 179234 541784 179290 541793
rect 179234 541719 179290 541728
rect 179340 531321 179368 576671
rect 179694 563612 179750 563621
rect 179694 563547 179750 563556
rect 179602 563136 179658 563145
rect 179602 563071 179658 563080
rect 179420 556504 179472 556510
rect 179420 556446 179472 556452
rect 179432 556345 179460 556446
rect 179418 556336 179474 556345
rect 179418 556271 179474 556280
rect 179418 556064 179474 556073
rect 179418 555999 179474 556008
rect 179432 555082 179460 555999
rect 179420 555076 179472 555082
rect 179420 555018 179472 555024
rect 179616 545766 179644 563071
rect 179604 545760 179656 545766
rect 179604 545702 179656 545708
rect 179708 541754 179736 563547
rect 179892 555257 179920 576671
rect 179984 557297 180012 594895
rect 254582 588704 254638 588713
rect 254582 588639 254638 588648
rect 254492 561060 254544 561066
rect 254492 561002 254544 561008
rect 253572 560652 253624 560658
rect 253572 560594 253624 560600
rect 253480 560516 253532 560522
rect 253480 560458 253532 560464
rect 246580 560448 246632 560454
rect 246284 560396 246580 560402
rect 246284 560390 246632 560396
rect 253018 560416 253074 560425
rect 246284 560374 246620 560390
rect 253018 560351 253074 560360
rect 245476 560312 245528 560318
rect 233422 560280 233478 560289
rect 245476 560254 245528 560260
rect 233422 560215 233478 560224
rect 216908 560144 216964 560153
rect 181502 559858 181530 560116
rect 182514 559858 182542 560116
rect 183526 559858 183554 560116
rect 184552 560102 184888 560130
rect 181502 559830 181576 559858
rect 182514 559830 182588 559858
rect 183526 559830 183600 559858
rect 180614 558920 180670 558929
rect 180614 558855 180670 558864
rect 180628 557598 180656 558855
rect 180706 558784 180762 558793
rect 180706 558719 180762 558728
rect 180720 557666 180748 558719
rect 180708 557660 180760 557666
rect 180708 557602 180760 557608
rect 180616 557592 180668 557598
rect 180616 557534 180668 557540
rect 179970 557288 180026 557297
rect 179970 557223 180026 557232
rect 179878 555248 179934 555257
rect 179878 555183 179934 555192
rect 180062 551440 180118 551449
rect 180062 551375 180118 551384
rect 180076 550730 180104 551375
rect 180064 550724 180116 550730
rect 180064 550666 180116 550672
rect 179696 541748 179748 541754
rect 179696 541690 179748 541696
rect 181548 541686 181576 559830
rect 182560 547194 182588 559830
rect 182548 547188 182600 547194
rect 182548 547130 182600 547136
rect 183572 545834 183600 559830
rect 184860 552702 184888 560102
rect 185550 559858 185578 560116
rect 186562 559858 186590 560116
rect 187574 559858 187602 560116
rect 188586 559858 188614 560116
rect 189612 560102 189948 560130
rect 185550 559830 185624 559858
rect 186562 559830 186636 559858
rect 187574 559830 187648 559858
rect 188586 559830 188660 559858
rect 184848 552696 184900 552702
rect 184848 552638 184900 552644
rect 185490 551440 185546 551449
rect 185490 551375 185546 551384
rect 185504 551041 185532 551375
rect 185490 551032 185546 551041
rect 185490 550967 185546 550976
rect 185596 547262 185624 559830
rect 185768 554872 185820 554878
rect 185768 554814 185820 554820
rect 185584 547256 185636 547262
rect 185584 547198 185636 547204
rect 183560 545828 183612 545834
rect 183560 545770 183612 545776
rect 181720 543856 181772 543862
rect 181720 543798 181772 543804
rect 181536 541680 181588 541686
rect 181536 541622 181588 541628
rect 179696 538280 179748 538286
rect 179696 538222 179748 538228
rect 179326 531312 179382 531321
rect 179326 531247 179382 531256
rect 179142 531176 179198 531185
rect 179142 531111 179198 531120
rect 178958 531040 179014 531049
rect 178868 531004 178920 531010
rect 178958 530975 179014 530984
rect 178868 530946 178920 530952
rect 178788 530862 179000 530890
rect 178868 530800 178920 530806
rect 178868 530742 178920 530748
rect 178880 526561 178908 530742
rect 178972 528554 179000 530862
rect 178972 528526 179092 528554
rect 178866 526552 178922 526561
rect 178866 526487 178922 526496
rect 179064 522889 179092 528526
rect 179050 522880 179106 522889
rect 179050 522815 179106 522824
rect 179708 520146 179736 538222
rect 180708 537056 180760 537062
rect 180708 536998 180760 537004
rect 180720 520146 180748 536998
rect 181732 520146 181760 543798
rect 184202 541648 184258 541657
rect 184202 541583 184258 541592
rect 183744 529984 183796 529990
rect 183744 529926 183796 529932
rect 182916 523116 182968 523122
rect 182916 523058 182968 523064
rect 182928 520146 182956 523058
rect 178696 520118 178740 520146
rect 179708 520118 179752 520146
rect 180720 520118 180764 520146
rect 181732 520118 181776 520146
rect 176688 519860 176716 520118
rect 177700 519860 177728 520118
rect 178712 519860 178740 520118
rect 179724 519860 179752 520118
rect 180736 519860 180764 520118
rect 181748 519860 181776 520118
rect 182760 520118 182956 520146
rect 183756 520146 183784 529926
rect 184216 522481 184244 541583
rect 184756 531344 184808 531350
rect 184756 531286 184808 531292
rect 184202 522472 184258 522481
rect 184202 522407 184258 522416
rect 184768 520146 184796 531286
rect 184848 522912 184900 522918
rect 184848 522854 184900 522860
rect 184860 521801 184888 522854
rect 184846 521792 184902 521801
rect 184846 521727 184902 521736
rect 185780 520146 185808 554814
rect 186608 536110 186636 559830
rect 187620 540394 187648 559830
rect 187792 546712 187844 546718
rect 187792 546654 187844 546660
rect 187608 540388 187660 540394
rect 187608 540330 187660 540336
rect 186596 536104 186648 536110
rect 186596 536046 186648 536052
rect 186872 525224 186924 525230
rect 186872 525166 186924 525172
rect 186884 520146 186912 525166
rect 183756 520118 183800 520146
rect 184768 520118 184812 520146
rect 185780 520118 185824 520146
rect 182760 519860 182788 520118
rect 183772 519860 183800 520118
rect 184784 519860 184812 520118
rect 185796 519860 185824 520118
rect 186808 520118 186912 520146
rect 187804 520146 187832 546654
rect 188632 533458 188660 559830
rect 189920 551342 189948 560102
rect 190610 559858 190638 560116
rect 191636 560102 191788 560130
rect 192648 560102 192984 560130
rect 190610 559830 190684 559858
rect 189908 551336 189960 551342
rect 189908 551278 189960 551284
rect 190656 540258 190684 559830
rect 191760 553110 191788 560102
rect 192956 554334 192984 560102
rect 193646 559858 193674 560116
rect 194658 559858 194686 560116
rect 195670 559858 195698 560116
rect 196682 559858 196710 560116
rect 197694 559858 197722 560116
rect 198706 559858 198734 560116
rect 199732 560102 199976 560130
rect 193646 559830 193720 559858
rect 194658 559830 194732 559858
rect 195670 559830 195744 559858
rect 196682 559830 196756 559858
rect 197694 559830 197768 559858
rect 198706 559830 198780 559858
rect 192944 554328 192996 554334
rect 192944 554270 192996 554276
rect 191748 553104 191800 553110
rect 191748 553046 191800 553052
rect 192852 545216 192904 545222
rect 192852 545158 192904 545164
rect 191104 543244 191156 543250
rect 191104 543186 191156 543192
rect 190644 540252 190696 540258
rect 190644 540194 190696 540200
rect 190828 536988 190880 536994
rect 190828 536930 190880 536936
rect 188620 533452 188672 533458
rect 188620 533394 188672 533400
rect 189908 527196 189960 527202
rect 189908 527138 189960 527144
rect 188988 520396 189040 520402
rect 188988 520338 189040 520344
rect 189000 520146 189028 520338
rect 189920 520146 189948 527138
rect 187804 520118 187848 520146
rect 186808 519860 186836 520118
rect 187820 519860 187848 520118
rect 188832 520118 189028 520146
rect 189844 520118 189948 520146
rect 190840 520146 190868 536930
rect 191116 521422 191144 543186
rect 191840 535560 191892 535566
rect 191840 535502 191892 535508
rect 191104 521416 191156 521422
rect 191104 521358 191156 521364
rect 191852 520146 191880 535502
rect 192864 520146 192892 545158
rect 193692 543046 193720 559830
rect 194704 543182 194732 559830
rect 194692 543176 194744 543182
rect 194692 543118 194744 543124
rect 193680 543040 193732 543046
rect 193680 542982 193732 542988
rect 195716 533594 195744 559830
rect 196728 545902 196756 559830
rect 196716 545896 196768 545902
rect 196716 545838 196768 545844
rect 197740 534818 197768 559830
rect 198752 548758 198780 559830
rect 199948 558346 199976 560102
rect 200730 559858 200758 560116
rect 201756 560102 202092 560130
rect 200730 559830 200804 559858
rect 199936 558340 199988 558346
rect 199936 558282 199988 558288
rect 198740 548752 198792 548758
rect 198740 548694 198792 548700
rect 200776 548622 200804 559830
rect 202064 557462 202092 560102
rect 202754 559858 202782 560116
rect 203780 560102 204116 560130
rect 202754 559830 202828 559858
rect 202052 557456 202104 557462
rect 202052 557398 202104 557404
rect 200764 548616 200816 548622
rect 200764 548558 200816 548564
rect 202800 544542 202828 559830
rect 204088 551478 204116 560102
rect 204778 559858 204806 560116
rect 205790 559858 205818 560116
rect 206802 559858 206830 560116
rect 207828 560102 208164 560130
rect 204778 559830 204852 559858
rect 205790 559830 205864 559858
rect 206802 559830 206876 559858
rect 204076 551472 204128 551478
rect 204076 551414 204128 551420
rect 202788 544536 202840 544542
rect 202788 544478 202840 544484
rect 204824 541657 204852 559830
rect 204810 541648 204866 541657
rect 204810 541583 204866 541592
rect 205836 537674 205864 559830
rect 206848 538966 206876 559830
rect 208136 552770 208164 560102
rect 208826 559858 208854 560116
rect 209838 559858 209866 560116
rect 210850 559858 210878 560116
rect 211862 559858 211890 560116
rect 212874 559858 212902 560116
rect 213886 559858 213914 560116
rect 214898 559858 214926 560116
rect 215910 559858 215938 560116
rect 216908 560079 216964 560088
rect 217934 559858 217962 560116
rect 218946 559858 218974 560116
rect 219958 559858 219986 560116
rect 220970 559858 220998 560116
rect 221982 559858 222010 560116
rect 222994 559858 223022 560116
rect 224006 559858 224034 560116
rect 225018 559858 225046 560116
rect 226030 559858 226058 560116
rect 227056 560102 227392 560130
rect 208826 559830 208900 559858
rect 209838 559830 209912 559858
rect 210850 559830 210924 559858
rect 211862 559830 211936 559858
rect 212874 559830 212948 559858
rect 213886 559830 213960 559858
rect 214898 559830 214972 559858
rect 215910 559830 215984 559858
rect 217934 559830 218008 559858
rect 218946 559830 219020 559858
rect 219958 559830 220032 559858
rect 220970 559830 221044 559858
rect 221982 559830 222056 559858
rect 222994 559830 223068 559858
rect 224006 559830 224080 559858
rect 225018 559830 225092 559858
rect 226030 559830 226104 559858
rect 208124 552764 208176 552770
rect 208124 552706 208176 552712
rect 208400 543652 208452 543658
rect 208400 543594 208452 543600
rect 208412 542745 208440 543594
rect 208872 542881 208900 559830
rect 209884 544474 209912 559830
rect 210896 550050 210924 559830
rect 210884 550044 210936 550050
rect 210884 549986 210936 549992
rect 211908 548690 211936 559830
rect 211896 548684 211948 548690
rect 211896 548626 211948 548632
rect 209872 544468 209924 544474
rect 209872 544410 209924 544416
rect 208858 542872 208914 542881
rect 208858 542807 208914 542816
rect 208398 542736 208454 542745
rect 208398 542671 208454 542680
rect 206836 538960 206888 538966
rect 206836 538902 206888 538908
rect 205824 537668 205876 537674
rect 205824 537610 205876 537616
rect 212920 534886 212948 559830
rect 213092 537124 213144 537130
rect 213092 537066 213144 537072
rect 212908 534880 212960 534886
rect 212908 534822 212960 534828
rect 197728 534812 197780 534818
rect 197728 534754 197780 534760
rect 211068 534336 211120 534342
rect 211068 534278 211120 534284
rect 209044 534268 209096 534274
rect 209044 534210 209096 534216
rect 195704 533588 195756 533594
rect 195704 533530 195756 533536
rect 194876 532908 194928 532914
rect 194876 532850 194928 532856
rect 193956 520940 194008 520946
rect 193956 520882 194008 520888
rect 193968 520146 193996 520882
rect 190840 520118 190884 520146
rect 191852 520118 191896 520146
rect 192864 520118 192908 520146
rect 188832 519860 188860 520118
rect 189844 519860 189872 520118
rect 190856 519860 190884 520118
rect 191868 519860 191896 520118
rect 192880 519860 192908 520118
rect 193892 520118 193996 520146
rect 194888 520146 194916 532850
rect 198924 531616 198976 531622
rect 198924 531558 198976 531564
rect 195888 530052 195940 530058
rect 195888 529994 195940 530000
rect 195900 520146 195928 529994
rect 198096 525972 198148 525978
rect 198096 525914 198148 525920
rect 197084 524680 197136 524686
rect 197084 524622 197136 524628
rect 197096 520146 197124 524622
rect 198108 520146 198136 525914
rect 194888 520118 194932 520146
rect 195900 520118 195944 520146
rect 193892 519860 193920 520118
rect 194904 519860 194932 520118
rect 195916 519860 195944 520118
rect 196928 520118 197124 520146
rect 197940 520118 198136 520146
rect 198936 520146 198964 531558
rect 208032 531548 208084 531554
rect 208032 531490 208084 531496
rect 202052 527400 202104 527406
rect 202052 527342 202104 527348
rect 200028 526040 200080 526046
rect 200028 525982 200080 525988
rect 200040 520146 200068 525982
rect 201040 524612 201092 524618
rect 201040 524554 201092 524560
rect 201052 520146 201080 524554
rect 202064 520146 202092 527342
rect 204168 527332 204220 527338
rect 204168 527274 204220 527280
rect 203064 523388 203116 523394
rect 203064 523330 203116 523336
rect 203076 520146 203104 523330
rect 204180 520146 204208 527274
rect 206192 523252 206244 523258
rect 206192 523194 206244 523200
rect 205180 521892 205232 521898
rect 205180 521834 205232 521840
rect 205192 520146 205220 521834
rect 206204 520146 206232 523194
rect 207204 520532 207256 520538
rect 207204 520474 207256 520480
rect 207216 520146 207244 520474
rect 198936 520118 198980 520146
rect 196928 519860 196956 520118
rect 197940 519860 197968 520118
rect 198952 519860 198980 520118
rect 199964 520118 200068 520146
rect 200976 520118 201080 520146
rect 201988 520118 202092 520146
rect 203000 520118 203104 520146
rect 204012 520118 204208 520146
rect 205024 520118 205220 520146
rect 206036 520118 206232 520146
rect 207048 520118 207244 520146
rect 208044 520146 208072 531490
rect 209056 520146 209084 534210
rect 210056 528760 210108 528766
rect 210056 528702 210108 528708
rect 210068 520146 210096 528702
rect 211080 520146 211108 534278
rect 212080 530120 212132 530126
rect 212080 530062 212132 530068
rect 212092 520146 212120 530062
rect 213104 520146 213132 537066
rect 213932 529446 213960 559830
rect 214104 531684 214156 531690
rect 214104 531626 214156 531632
rect 213920 529440 213972 529446
rect 213920 529382 213972 529388
rect 214116 520146 214144 531626
rect 214944 526969 214972 559830
rect 215116 532976 215168 532982
rect 215116 532918 215168 532924
rect 214930 526960 214986 526969
rect 214564 526924 214616 526930
rect 214930 526895 214986 526904
rect 214564 526866 214616 526872
rect 214576 526153 214604 526866
rect 214562 526144 214618 526153
rect 214562 526079 214618 526088
rect 215128 520146 215156 532918
rect 215956 532681 215984 559830
rect 216680 559632 216732 559638
rect 216680 559574 216732 559580
rect 216692 559201 216720 559574
rect 216678 559192 216734 559201
rect 216678 559127 216734 559136
rect 216680 544808 216732 544814
rect 216680 544750 216732 544756
rect 216692 543833 216720 544750
rect 217980 544105 218008 559830
rect 218152 545148 218204 545154
rect 218152 545090 218204 545096
rect 217966 544096 218022 544105
rect 217966 544031 218022 544040
rect 216678 543824 216734 543833
rect 216678 543759 216734 543768
rect 218060 540796 218112 540802
rect 218060 540738 218112 540744
rect 217140 539776 217192 539782
rect 217140 539718 217192 539724
rect 216128 535696 216180 535702
rect 216128 535638 216180 535644
rect 215942 532672 215998 532681
rect 215300 532636 215352 532642
rect 215942 532607 215998 532616
rect 215300 532578 215352 532584
rect 215312 531457 215340 532578
rect 215298 531448 215354 531457
rect 215298 531383 215354 531392
rect 216140 520146 216168 535638
rect 217152 520146 217180 539718
rect 218072 539617 218100 540738
rect 218058 539608 218114 539617
rect 218058 539543 218114 539552
rect 218164 520146 218192 545090
rect 218992 540297 219020 559830
rect 219164 553512 219216 553518
rect 219164 553454 219216 553460
rect 218978 540288 219034 540297
rect 218978 540223 219034 540232
rect 219176 520146 219204 553454
rect 220004 520713 220032 559830
rect 220176 554940 220228 554946
rect 220176 554882 220228 554888
rect 219990 520704 220046 520713
rect 219990 520639 220046 520648
rect 220188 520146 220216 554882
rect 220728 521416 220780 521422
rect 220728 521358 220780 521364
rect 220740 520441 220768 521358
rect 221016 521121 221044 559830
rect 221188 549364 221240 549370
rect 221188 549306 221240 549312
rect 221002 521112 221058 521121
rect 221002 521047 221058 521056
rect 220726 520432 220782 520441
rect 220726 520367 220782 520376
rect 221200 520146 221228 549306
rect 222028 539617 222056 559830
rect 222014 539608 222070 539617
rect 222014 539543 222070 539552
rect 222108 539300 222160 539306
rect 222108 539242 222160 539248
rect 222120 538257 222148 539242
rect 222106 538248 222162 538257
rect 222106 538183 222162 538192
rect 223040 533361 223068 559830
rect 224052 545329 224080 559830
rect 224224 550792 224276 550798
rect 224224 550734 224276 550740
rect 224132 546168 224184 546174
rect 224132 546110 224184 546116
rect 224144 546009 224172 546110
rect 224130 546000 224186 546009
rect 224130 545935 224186 545944
rect 224038 545320 224094 545329
rect 224038 545255 224094 545264
rect 223488 533860 223540 533866
rect 223488 533802 223540 533808
rect 223026 533352 223082 533361
rect 223026 533287 223082 533296
rect 223500 532817 223528 533802
rect 223486 532808 223542 532817
rect 223486 532743 223542 532752
rect 222384 524748 222436 524754
rect 222384 524690 222436 524696
rect 222108 521280 222160 521286
rect 222106 521248 222108 521257
rect 222160 521248 222162 521257
rect 222106 521183 222162 521192
rect 222396 520146 222424 524690
rect 223304 523320 223356 523326
rect 223304 523262 223356 523268
rect 223316 520146 223344 523262
rect 224130 523016 224186 523025
rect 224130 522951 224186 522960
rect 224144 522850 224172 522951
rect 224132 522844 224184 522850
rect 224132 522786 224184 522792
rect 208044 520118 208088 520146
rect 209056 520118 209100 520146
rect 210068 520118 210112 520146
rect 211080 520118 211124 520146
rect 212092 520118 212136 520146
rect 213104 520118 213148 520146
rect 214116 520118 214160 520146
rect 215128 520118 215172 520146
rect 216140 520118 216184 520146
rect 217152 520118 217196 520146
rect 218164 520118 218208 520146
rect 219176 520118 219220 520146
rect 220188 520118 220232 520146
rect 221200 520118 221244 520146
rect 199964 519860 199992 520118
rect 200976 519860 201004 520118
rect 201988 519860 202016 520118
rect 203000 519860 203028 520118
rect 204012 519860 204040 520118
rect 205024 519860 205052 520118
rect 206036 519860 206064 520118
rect 207048 519860 207076 520118
rect 208060 519860 208088 520118
rect 209072 519860 209100 520118
rect 210084 519860 210112 520118
rect 211096 519860 211124 520118
rect 212108 519860 212136 520118
rect 213120 519860 213148 520118
rect 214132 519860 214160 520118
rect 215144 519860 215172 520118
rect 216156 519860 216184 520118
rect 217168 519860 217196 520118
rect 218180 519860 218208 520118
rect 219192 519860 219220 520118
rect 220204 519860 220232 520118
rect 221216 519860 221244 520118
rect 222228 520118 222424 520146
rect 223240 520118 223344 520146
rect 224236 520146 224264 550734
rect 225064 538801 225092 559830
rect 226076 550118 226104 559830
rect 226246 558512 226302 558521
rect 226246 558447 226302 558456
rect 226064 550112 226116 550118
rect 226064 550054 226116 550060
rect 225510 539608 225566 539617
rect 225510 539543 225566 539552
rect 225050 538792 225106 538801
rect 225050 538727 225106 538736
rect 225524 538490 225552 539543
rect 225512 538484 225564 538490
rect 225512 538426 225564 538432
rect 224314 533216 224370 533225
rect 224314 533151 224370 533160
rect 224328 522209 224356 533151
rect 224960 525428 225012 525434
rect 224960 525370 225012 525376
rect 224972 524657 225000 525370
rect 225326 524920 225382 524929
rect 225326 524855 225382 524864
rect 224958 524648 225014 524657
rect 224958 524583 225014 524592
rect 224314 522200 224370 522209
rect 224314 522135 224370 522144
rect 225340 520146 225368 524855
rect 224236 520118 224280 520146
rect 222228 519860 222256 520118
rect 223240 519860 223268 520118
rect 224252 519860 224280 520118
rect 225264 520118 225368 520146
rect 226260 520146 226288 558447
rect 226338 555792 226394 555801
rect 226338 555727 226394 555736
rect 226352 555150 226380 555727
rect 226340 555144 226392 555150
rect 226340 555086 226392 555092
rect 227258 555112 227314 555121
rect 227258 555047 227314 555056
rect 227272 552537 227300 555047
rect 227364 553353 227392 560102
rect 228054 559858 228082 560116
rect 229080 560102 229232 560130
rect 230092 560102 230428 560130
rect 228054 559830 228128 559858
rect 227718 557424 227774 557433
rect 227718 557359 227774 557368
rect 227732 556578 227760 557359
rect 227720 556572 227772 556578
rect 227720 556514 227772 556520
rect 227350 553344 227406 553353
rect 227350 553279 227406 553288
rect 227258 552528 227314 552537
rect 227258 552463 227314 552472
rect 226982 539064 227038 539073
rect 226982 538999 227038 539008
rect 226996 523025 227024 538999
rect 226982 523016 227038 523025
rect 226982 522951 227038 522960
rect 226340 522708 226392 522714
rect 226340 522650 226392 522656
rect 226352 522073 226380 522650
rect 226338 522064 226394 522073
rect 226338 521999 226394 522008
rect 227272 520146 227300 552463
rect 228100 548729 228128 559830
rect 228270 556472 228326 556481
rect 228270 556407 228326 556416
rect 228284 551313 228312 556407
rect 228270 551304 228326 551313
rect 228270 551239 228326 551248
rect 228086 548720 228142 548729
rect 228086 548655 228142 548664
rect 227718 548448 227774 548457
rect 227718 548383 227774 548392
rect 227732 548146 227760 548383
rect 227720 548140 227772 548146
rect 227720 548082 227772 548088
rect 227720 522776 227772 522782
rect 227720 522718 227772 522724
rect 227732 521937 227760 522718
rect 227718 521928 227774 521937
rect 227718 521863 227774 521872
rect 228284 520146 228312 551239
rect 228362 549944 228418 549953
rect 228362 549879 228418 549888
rect 228376 522617 228404 549879
rect 229204 547874 229232 560102
rect 230400 557534 230428 560102
rect 231090 559858 231118 560116
rect 232102 559858 232130 560116
rect 233114 559858 233142 560116
rect 231090 559830 231164 559858
rect 232102 559830 232176 559858
rect 233114 559830 233188 559858
rect 230308 557506 230428 557534
rect 230202 557424 230258 557433
rect 230202 557359 230258 557368
rect 230216 555257 230244 557359
rect 230202 555248 230258 555257
rect 230124 555206 230202 555234
rect 229282 549808 229338 549817
rect 229282 549743 229338 549752
rect 229112 547846 229232 547874
rect 229112 528018 229140 547846
rect 229100 528012 229152 528018
rect 229100 527954 229152 527960
rect 228362 522608 228418 522617
rect 228362 522543 228418 522552
rect 229296 520146 229324 549743
rect 230124 547874 230152 555206
rect 230202 555183 230258 555192
rect 230202 553752 230258 553761
rect 230202 553687 230258 553696
rect 230216 549817 230244 553687
rect 230308 551290 230336 557506
rect 230388 556640 230440 556646
rect 230386 556608 230388 556617
rect 230440 556608 230442 556617
rect 230386 556543 230442 556552
rect 230388 554464 230440 554470
rect 230386 554432 230388 554441
rect 230440 554432 230442 554441
rect 230386 554367 230442 554376
rect 230386 551304 230442 551313
rect 230308 551262 230386 551290
rect 230386 551239 230442 551248
rect 230202 549808 230258 549817
rect 230202 549743 230258 549752
rect 230124 547846 230336 547874
rect 230308 520146 230336 547846
rect 231136 547233 231164 559830
rect 231768 558544 231820 558550
rect 231768 558486 231820 558492
rect 231214 558104 231270 558113
rect 231214 558039 231270 558048
rect 231228 557534 231256 558039
rect 231780 557705 231808 558486
rect 231766 557696 231822 557705
rect 231766 557631 231822 557640
rect 231228 557506 231348 557534
rect 231122 547224 231178 547233
rect 231122 547159 231178 547168
rect 231320 536625 231348 557506
rect 231766 547360 231822 547369
rect 231766 547295 231822 547304
rect 231780 546854 231808 547295
rect 231768 546848 231820 546854
rect 231768 546790 231820 546796
rect 231306 536616 231362 536625
rect 231306 536551 231362 536560
rect 231320 520146 231348 536551
rect 232148 528086 232176 559830
rect 232318 549808 232374 549817
rect 232318 549743 232374 549752
rect 232332 548321 232360 549743
rect 232318 548312 232374 548321
rect 232318 548247 232374 548256
rect 232136 528080 232188 528086
rect 232136 528022 232188 528028
rect 231768 527672 231820 527678
rect 231768 527614 231820 527620
rect 231780 521354 231808 527614
rect 231768 521348 231820 521354
rect 231768 521290 231820 521296
rect 232332 520146 232360 548247
rect 233160 536625 233188 559830
rect 233436 547874 233464 560215
rect 233698 560144 233754 560153
rect 233698 560079 233754 560088
rect 233712 559366 233740 560079
rect 234126 559858 234154 560116
rect 235138 559858 235166 560116
rect 236164 560102 236500 560130
rect 234126 559830 234200 559858
rect 235138 559830 235212 559858
rect 233700 559360 233752 559366
rect 233700 559302 233752 559308
rect 233344 547846 233464 547874
rect 233146 536616 233202 536625
rect 233146 536551 233202 536560
rect 233344 520146 233372 547846
rect 233884 526856 233936 526862
rect 233884 526798 233936 526804
rect 233896 526017 233924 526798
rect 234172 526697 234200 559830
rect 234342 555792 234398 555801
rect 234342 555727 234398 555736
rect 234356 550633 234384 555727
rect 234618 553344 234674 553353
rect 234618 553279 234674 553288
rect 234632 552090 234660 553279
rect 234620 552084 234672 552090
rect 234620 552026 234672 552032
rect 234342 550624 234398 550633
rect 234342 550559 234398 550568
rect 234158 526688 234214 526697
rect 234158 526623 234214 526632
rect 233882 526008 233938 526017
rect 233882 525943 233938 525952
rect 234356 520146 234384 550559
rect 235184 547369 235212 559830
rect 236366 558648 236422 558657
rect 236366 558583 236422 558592
rect 235354 552528 235410 552537
rect 235354 552463 235410 552472
rect 235170 547360 235226 547369
rect 235170 547295 235226 547304
rect 235368 546825 235396 552463
rect 235998 551576 236054 551585
rect 235998 551511 236054 551520
rect 236012 550866 236040 551511
rect 236000 550860 236052 550866
rect 236000 550802 236052 550808
rect 235354 546816 235410 546825
rect 235354 546751 235410 546760
rect 235368 520146 235396 546751
rect 235998 541648 236054 541657
rect 235998 541583 236054 541592
rect 236012 541278 236040 541583
rect 236000 541272 236052 541278
rect 236000 541214 236052 541220
rect 236380 520146 236408 558583
rect 236472 551041 236500 560102
rect 237162 559858 237190 560116
rect 238174 559858 238202 560116
rect 239186 559858 239214 560116
rect 240198 559858 240226 560116
rect 241210 559858 241238 560116
rect 242222 559858 242250 560116
rect 243234 559858 243262 560116
rect 244246 559858 244274 560116
rect 244462 559872 244518 559881
rect 237162 559830 237236 559858
rect 238174 559830 238248 559858
rect 239186 559830 239260 559858
rect 240198 559830 240272 559858
rect 241210 559830 241284 559858
rect 242222 559830 242296 559858
rect 243234 559830 243308 559858
rect 244246 559830 244320 559858
rect 236458 551032 236514 551041
rect 236458 550967 236514 550976
rect 237208 541657 237236 559830
rect 237378 559328 237434 559337
rect 237378 559263 237434 559272
rect 237194 541648 237250 541657
rect 237194 541583 237250 541592
rect 237392 520146 237420 559263
rect 238220 526969 238248 559830
rect 238390 558376 238446 558385
rect 238390 558311 238446 558320
rect 237470 526960 237526 526969
rect 237470 526895 237526 526904
rect 238206 526960 238262 526969
rect 238206 526895 238262 526904
rect 237484 526114 237512 526895
rect 237472 526108 237524 526114
rect 237472 526050 237524 526056
rect 238404 520146 238432 558311
rect 239232 543289 239260 559830
rect 240138 559464 240194 559473
rect 240138 559399 240194 559408
rect 240046 555520 240102 555529
rect 240046 555455 240102 555464
rect 240060 554713 240088 555455
rect 240152 554849 240180 559399
rect 240138 554840 240194 554849
rect 240138 554775 240194 554784
rect 239402 554704 239458 554713
rect 239402 554639 239458 554648
rect 240046 554704 240102 554713
rect 240046 554639 240102 554648
rect 239218 543280 239274 543289
rect 239218 543215 239274 543224
rect 239416 520146 239444 554639
rect 240048 554396 240100 554402
rect 240048 554338 240100 554344
rect 240060 553625 240088 554338
rect 240046 553616 240102 553625
rect 240046 553551 240102 553560
rect 240048 543584 240100 543590
rect 240048 543526 240100 543532
rect 240060 542609 240088 543526
rect 240046 542600 240102 542609
rect 240046 542535 240102 542544
rect 240244 523297 240272 559830
rect 240414 559192 240470 559201
rect 240414 559127 240470 559136
rect 240428 554577 240456 559127
rect 240414 554568 240470 554577
rect 240414 554503 240470 554512
rect 240230 523288 240286 523297
rect 240230 523223 240286 523232
rect 240428 520146 240456 554503
rect 241256 536217 241284 559830
rect 241426 556064 241482 556073
rect 241426 555999 241482 556008
rect 241440 554849 241468 555999
rect 241426 554840 241482 554849
rect 241426 554775 241482 554784
rect 241334 536616 241390 536625
rect 241334 536551 241390 536560
rect 241242 536208 241298 536217
rect 241242 536143 241298 536152
rect 241348 535634 241376 536551
rect 241336 535628 241388 535634
rect 241336 535570 241388 535576
rect 241336 524136 241388 524142
rect 241336 524078 241388 524084
rect 241348 523841 241376 524078
rect 241334 523832 241390 523841
rect 241334 523767 241390 523776
rect 241440 520146 241468 554775
rect 242268 543153 242296 559830
rect 242438 557152 242494 557161
rect 242438 557087 242494 557096
rect 242254 543144 242310 543153
rect 242254 543079 242310 543088
rect 242452 520146 242480 557087
rect 243280 549953 243308 559830
rect 243450 558784 243506 558793
rect 243450 558719 243506 558728
rect 243464 558249 243492 558719
rect 243450 558240 243506 558249
rect 243450 558175 243506 558184
rect 243266 549944 243322 549953
rect 243266 549879 243322 549888
rect 242806 542872 242862 542881
rect 242806 542807 242862 542816
rect 242820 542570 242848 542807
rect 242808 542564 242860 542570
rect 242808 542506 242860 542512
rect 243464 520146 243492 558175
rect 244292 557534 244320 559830
rect 245258 559858 245286 560116
rect 245488 560017 245516 560254
rect 248602 560144 248658 560153
rect 245474 560008 245530 560017
rect 245474 559943 245530 559952
rect 245258 559830 245332 559858
rect 244462 559807 244518 559816
rect 244292 557506 244412 557534
rect 244280 543516 244332 543522
rect 244280 543458 244332 543464
rect 244292 542473 244320 543458
rect 244384 542881 244412 557506
rect 244370 542872 244426 542881
rect 244370 542807 244426 542816
rect 244278 542464 244334 542473
rect 244278 542399 244334 542408
rect 244278 540288 244334 540297
rect 244278 540223 244334 540232
rect 244292 539986 244320 540223
rect 244280 539980 244332 539986
rect 244280 539922 244332 539928
rect 244476 520146 244504 559807
rect 245304 540025 245332 559830
rect 245290 540016 245346 540025
rect 245290 539951 245346 539960
rect 245488 520146 245516 559943
rect 247282 559858 247310 560116
rect 248294 559858 248322 560116
rect 248602 560079 248658 560088
rect 247282 559830 247356 559858
rect 248294 559830 248368 559858
rect 246394 559736 246450 559745
rect 246394 559671 246450 559680
rect 246408 558929 246436 559671
rect 246394 558920 246450 558929
rect 246394 558855 246450 558864
rect 245660 558476 245712 558482
rect 245660 558418 245712 558424
rect 245672 557569 245700 558418
rect 245658 557560 245714 557569
rect 246408 557534 246436 558855
rect 246408 557506 246528 557534
rect 245658 557495 245714 557504
rect 246304 546780 246356 546786
rect 246304 546722 246356 546728
rect 246316 525162 246344 546722
rect 246304 525156 246356 525162
rect 246304 525098 246356 525104
rect 246500 520146 246528 557506
rect 247130 557288 247186 557297
rect 247130 557223 247186 557232
rect 247144 555257 247172 557223
rect 247130 555248 247186 555257
rect 247040 555212 247092 555218
rect 247130 555183 247186 555192
rect 247040 555154 247092 555160
rect 247052 554985 247080 555154
rect 247038 554976 247094 554985
rect 247038 554911 247094 554920
rect 247038 540424 247094 540433
rect 247038 540359 247094 540368
rect 247052 539918 247080 540359
rect 247328 540297 247356 559830
rect 247498 555248 247554 555257
rect 247498 555183 247554 555192
rect 247314 540288 247370 540297
rect 247314 540223 247370 540232
rect 247040 539912 247092 539918
rect 247040 539854 247092 539860
rect 247040 526176 247092 526182
rect 247040 526118 247092 526124
rect 247052 525638 247080 526118
rect 247040 525632 247092 525638
rect 247040 525574 247092 525580
rect 247040 525496 247092 525502
rect 247040 525438 247092 525444
rect 247052 524521 247080 525438
rect 247038 524512 247094 524521
rect 247038 524447 247094 524456
rect 247512 520146 247540 555183
rect 248340 525065 248368 559830
rect 248616 557534 248644 560079
rect 249306 559858 249334 560116
rect 250318 559858 250346 560116
rect 251330 559858 251358 560116
rect 252342 559858 252370 560116
rect 249306 559830 249380 559858
rect 250318 559830 250392 559858
rect 251330 559830 251404 559858
rect 252342 559830 252416 559858
rect 248524 557506 248644 557534
rect 248524 553353 248552 557506
rect 248510 553344 248566 553353
rect 248510 553279 248566 553288
rect 248326 525056 248382 525065
rect 248326 524991 248382 525000
rect 248524 520146 248552 553279
rect 249352 526425 249380 559830
rect 249522 553888 249578 553897
rect 249522 553823 249578 553832
rect 249338 526416 249394 526425
rect 249338 526351 249394 526360
rect 249536 520146 249564 553823
rect 249706 552800 249762 552809
rect 249706 552735 249762 552744
rect 249720 552226 249748 552735
rect 249708 552220 249760 552226
rect 249708 552162 249760 552168
rect 250364 534857 250392 559830
rect 250534 557288 250590 557297
rect 250534 557223 250590 557232
rect 250444 557048 250496 557054
rect 250444 556990 250496 556996
rect 250456 544814 250484 556990
rect 250444 544808 250496 544814
rect 250444 544750 250496 544756
rect 250350 534848 250406 534857
rect 250350 534783 250406 534792
rect 249708 526720 249760 526726
rect 249708 526662 249760 526668
rect 249720 525881 249748 526662
rect 249706 525872 249762 525881
rect 249706 525807 249762 525816
rect 250548 520146 250576 557223
rect 251376 544785 251404 559830
rect 251824 558340 251876 558346
rect 251824 558282 251876 558288
rect 251546 557560 251602 557569
rect 251546 557495 251602 557504
rect 251362 544776 251418 544785
rect 251362 544711 251418 544720
rect 251088 535288 251140 535294
rect 251088 535230 251140 535236
rect 251100 534177 251128 535230
rect 251086 534168 251142 534177
rect 251086 534103 251142 534112
rect 251560 520146 251588 557495
rect 251836 544678 251864 558282
rect 251824 544672 251876 544678
rect 251824 544614 251876 544620
rect 252388 537577 252416 559830
rect 252558 559056 252614 559065
rect 252558 558991 252614 559000
rect 252466 557968 252522 557977
rect 252466 557903 252522 557912
rect 252480 557734 252508 557903
rect 252468 557728 252520 557734
rect 252468 557670 252520 557676
rect 252466 544096 252522 544105
rect 252466 544031 252522 544040
rect 252480 543930 252508 544031
rect 252468 543924 252520 543930
rect 252468 543866 252520 543872
rect 252468 538076 252520 538082
rect 252468 538018 252520 538024
rect 252374 537568 252430 537577
rect 252374 537503 252430 537512
rect 252480 536897 252508 538018
rect 252466 536888 252522 536897
rect 252466 536823 252522 536832
rect 251824 533044 251876 533050
rect 251824 532986 251876 532992
rect 251836 522442 251864 532986
rect 251824 522436 251876 522442
rect 251824 522378 251876 522384
rect 252572 520146 252600 558991
rect 253032 553110 253060 560351
rect 253354 559858 253382 560116
rect 253354 559830 253428 559858
rect 253020 553104 253072 553110
rect 253020 553046 253072 553052
rect 253202 552936 253258 552945
rect 253202 552871 253258 552880
rect 253216 552294 253244 552871
rect 253204 552288 253256 552294
rect 253204 552230 253256 552236
rect 253204 548072 253256 548078
rect 253204 548014 253256 548020
rect 253216 525230 253244 548014
rect 253400 539073 253428 559830
rect 253492 544882 253520 560458
rect 253584 554334 253612 560594
rect 254400 560584 254452 560590
rect 254400 560526 254452 560532
rect 254412 557462 254440 560526
rect 254400 557456 254452 557462
rect 254400 557398 254452 557404
rect 253572 554328 253624 554334
rect 253572 554270 253624 554276
rect 253570 552936 253626 552945
rect 253570 552871 253626 552880
rect 253480 544876 253532 544882
rect 253480 544818 253532 544824
rect 253386 539064 253442 539073
rect 253386 538999 253442 539008
rect 253204 525224 253256 525230
rect 253204 525166 253256 525172
rect 253202 522744 253258 522753
rect 253202 522679 253258 522688
rect 253216 522238 253244 522679
rect 253204 522232 253256 522238
rect 253204 522174 253256 522180
rect 253584 520146 253612 552871
rect 254504 548962 254532 561002
rect 254596 556073 254624 588639
rect 255042 577824 255098 577833
rect 255042 577759 255098 577768
rect 254950 576464 255006 576473
rect 254950 576399 255006 576408
rect 254766 575648 254822 575657
rect 254766 575583 254822 575592
rect 254676 560720 254728 560726
rect 254676 560662 254728 560668
rect 254582 556064 254638 556073
rect 254582 555999 254638 556008
rect 254492 548956 254544 548962
rect 254492 548898 254544 548904
rect 253938 546408 253994 546417
rect 253938 546343 253994 546352
rect 253952 545222 253980 546343
rect 253940 545216 253992 545222
rect 253940 545158 253992 545164
rect 253662 539200 253718 539209
rect 253662 539135 253718 539144
rect 253676 522073 253704 539135
rect 254582 538656 254638 538665
rect 254582 538591 254638 538600
rect 253662 522064 253718 522073
rect 253662 521999 253718 522008
rect 254596 520146 254624 538591
rect 254688 526794 254716 560662
rect 254780 553761 254808 575583
rect 254860 560652 254912 560658
rect 254860 560594 254912 560600
rect 254766 553752 254822 553761
rect 254766 553687 254822 553696
rect 254872 540734 254900 560594
rect 254964 557433 254992 576399
rect 255056 558113 255084 577759
rect 255226 574560 255282 574569
rect 255226 574495 255282 574504
rect 255134 573200 255190 573209
rect 255134 573135 255190 573144
rect 255042 558104 255098 558113
rect 255042 558039 255098 558048
rect 254950 557424 255006 557433
rect 254950 557359 255006 557368
rect 255044 556708 255096 556714
rect 255044 556650 255096 556656
rect 255056 543318 255084 556650
rect 255148 555121 255176 573135
rect 255240 556481 255268 574495
rect 255226 556472 255282 556481
rect 255226 556407 255282 556416
rect 255134 555112 255190 555121
rect 255134 555047 255190 555056
rect 255044 543312 255096 543318
rect 255044 543254 255096 543260
rect 254860 540728 254912 540734
rect 254860 540670 254912 540676
rect 254768 539980 254820 539986
rect 254768 539922 254820 539928
rect 254676 526788 254728 526794
rect 254676 526730 254728 526736
rect 254780 521014 254808 539922
rect 254860 531752 254912 531758
rect 254860 531694 254912 531700
rect 254872 522374 254900 531694
rect 254860 522368 254912 522374
rect 254860 522310 254912 522316
rect 254768 521008 254820 521014
rect 254768 520950 254820 520956
rect 255608 520146 255636 635695
rect 255962 633448 256018 633457
rect 255962 633383 256018 633392
rect 255976 600273 256004 633383
rect 255962 600264 256018 600273
rect 255962 600199 256018 600208
rect 255962 594144 256018 594153
rect 255962 594079 256018 594088
rect 255870 584352 255926 584361
rect 255870 584287 255926 584296
rect 255884 559337 255912 584287
rect 255870 559328 255926 559337
rect 255870 559263 255926 559272
rect 255976 558929 256004 594079
rect 256054 589792 256110 589801
rect 256054 589727 256110 589736
rect 255962 558920 256018 558929
rect 255962 558855 256018 558864
rect 256068 557161 256096 589727
rect 256422 587616 256478 587625
rect 256422 587551 256478 587560
rect 256330 585440 256386 585449
rect 256330 585375 256386 585384
rect 256238 582176 256294 582185
rect 256238 582111 256294 582120
rect 256146 578912 256202 578921
rect 256146 578847 256202 578856
rect 256054 557152 256110 557161
rect 256054 557087 256110 557096
rect 256160 549817 256188 578847
rect 256252 552537 256280 582111
rect 256344 558385 256372 585375
rect 256436 559201 256464 587551
rect 256514 569256 256570 569265
rect 256514 569191 256570 569200
rect 256422 559192 256478 559201
rect 256422 559127 256478 559136
rect 256330 558376 256386 558385
rect 256330 558311 256386 558320
rect 256528 553353 256556 569191
rect 256514 553344 256570 553353
rect 256514 553279 256570 553288
rect 256238 552528 256294 552537
rect 256238 552463 256294 552472
rect 256146 549808 256202 549817
rect 256146 549743 256202 549752
rect 256620 520146 256648 638143
rect 257986 598904 258042 598913
rect 257986 598839 258042 598848
rect 257710 575512 257766 575521
rect 257710 575447 257766 575456
rect 257526 572928 257582 572937
rect 257526 572863 257582 572872
rect 257540 558385 257568 572863
rect 257618 571840 257674 571849
rect 257618 571775 257674 571784
rect 257526 558376 257582 558385
rect 257526 558311 257582 558320
rect 257632 555529 257660 571775
rect 257724 559745 257752 575447
rect 257802 572792 257858 572801
rect 257802 572727 257858 572736
rect 257710 559736 257766 559745
rect 257710 559671 257766 559680
rect 257618 555520 257674 555529
rect 257618 555455 257674 555464
rect 257816 554441 257844 572727
rect 257894 572656 257950 572665
rect 257894 572591 257950 572600
rect 257802 554432 257858 554441
rect 257802 554367 257858 554376
rect 256700 554328 256752 554334
rect 256700 554270 256752 554276
rect 256712 553489 256740 554270
rect 256698 553480 256754 553489
rect 256698 553415 256754 553424
rect 256698 553344 256754 553353
rect 256698 553279 256754 553288
rect 256712 552945 256740 553279
rect 256698 552936 256754 552945
rect 256698 552871 256754 552880
rect 257908 530505 257936 572591
rect 258000 554577 258028 598839
rect 257986 554568 258042 554577
rect 257986 554503 258042 554512
rect 256698 530496 256754 530505
rect 256698 530431 256754 530440
rect 257894 530496 257950 530505
rect 257894 530431 257950 530440
rect 256712 530398 256740 530431
rect 256700 530392 256752 530398
rect 256700 530334 256752 530340
rect 256698 526688 256754 526697
rect 256698 526623 256754 526632
rect 256712 526182 256740 526623
rect 256700 526176 256752 526182
rect 256700 526118 256752 526124
rect 258092 524929 258120 638279
rect 258170 599584 258226 599593
rect 258170 599519 258226 599528
rect 258184 557569 258212 599519
rect 258736 598505 258764 638415
rect 259380 638353 259408 640999
rect 259366 638344 259422 638353
rect 259366 638279 259422 638288
rect 258906 635624 258962 635633
rect 258906 635559 258962 635568
rect 258722 598496 258778 598505
rect 258722 598431 258778 598440
rect 258736 596174 258764 598431
rect 258920 597417 258948 635559
rect 258906 597408 258962 597417
rect 258906 597343 258962 597352
rect 258644 596146 258764 596174
rect 258644 584610 258672 596146
rect 258644 584582 258856 584610
rect 258724 584452 258776 584458
rect 258724 584394 258776 584400
rect 258170 557560 258226 557569
rect 258170 557495 258226 557504
rect 258736 553897 258764 584394
rect 258828 557297 258856 584582
rect 258920 584458 258948 597343
rect 259090 595232 259146 595241
rect 259090 595167 259146 595176
rect 258908 584452 258960 584458
rect 258908 584394 258960 584400
rect 259104 582434 259132 595167
rect 259366 591968 259422 591977
rect 259366 591903 259422 591912
rect 258920 582406 259132 582434
rect 258814 557288 258870 557297
rect 258814 557223 258870 557232
rect 258920 555257 258948 582406
rect 259380 582374 259408 591903
rect 259012 582346 259408 582374
rect 259012 559881 259040 582346
rect 259090 561776 259146 561785
rect 259090 561711 259146 561720
rect 259184 561740 259236 561746
rect 258998 559872 259054 559881
rect 258998 559807 259054 559816
rect 259000 556980 259052 556986
rect 259000 556922 259052 556928
rect 258906 555248 258962 555257
rect 258906 555183 258962 555192
rect 258722 553888 258778 553897
rect 258722 553823 258778 553832
rect 258630 546952 258686 546961
rect 258630 546887 258686 546896
rect 258078 524920 258134 524929
rect 258078 524855 258134 524864
rect 257526 522880 257582 522889
rect 257582 522838 257660 522866
rect 257526 522815 257582 522824
rect 256698 522744 256754 522753
rect 256698 522679 256754 522688
rect 256712 521762 256740 522679
rect 256700 521756 256752 521762
rect 256700 521698 256752 521704
rect 257632 520146 257660 522838
rect 258644 520146 258672 546887
rect 259012 522374 259040 556922
rect 259104 533769 259132 561711
rect 259184 561682 259236 561688
rect 259196 543522 259224 561682
rect 259184 543516 259236 543522
rect 259184 543458 259236 543464
rect 259090 533760 259146 533769
rect 259090 533695 259146 533704
rect 259000 522368 259052 522374
rect 259000 522310 259052 522316
rect 259656 520146 259684 643855
rect 260194 637256 260250 637265
rect 260194 637191 260250 637200
rect 260104 617568 260156 617574
rect 260104 617510 260156 617516
rect 260116 556714 260144 617510
rect 260208 601769 260236 637191
rect 260286 635488 260342 635497
rect 260286 635423 260342 635432
rect 260194 601760 260250 601769
rect 260194 601695 260250 601704
rect 260104 556708 260156 556714
rect 260104 556650 260156 556656
rect 260208 553353 260236 601695
rect 260300 600681 260328 635423
rect 260654 634672 260710 634681
rect 260654 634607 260710 634616
rect 260286 600672 260342 600681
rect 260286 600607 260342 600616
rect 260300 559065 260328 600607
rect 260286 559056 260342 559065
rect 260286 558991 260342 559000
rect 260194 553344 260250 553353
rect 260194 553279 260250 553288
rect 260668 520146 260696 634607
rect 261680 520146 261708 643991
rect 297270 643784 297326 643793
rect 297270 643719 297326 643728
rect 294050 642968 294106 642977
rect 294050 642903 294106 642912
rect 294064 642462 294092 642903
rect 294052 642456 294104 642462
rect 293958 642424 294014 642433
rect 294052 642398 294104 642404
rect 293958 642359 293960 642368
rect 294012 642359 294014 642368
rect 293960 642330 294012 642336
rect 294786 642288 294842 642297
rect 294786 642223 294842 642232
rect 294602 642152 294658 642161
rect 294602 642087 294658 642096
rect 262678 641200 262734 641209
rect 262678 641135 262734 641144
rect 262692 520146 262720 641135
rect 291844 638376 291896 638382
rect 291844 638318 291896 638324
rect 287702 636848 287758 636857
rect 287702 636783 287758 636792
rect 285034 634808 285090 634817
rect 285034 634743 285090 634752
rect 263690 634536 263746 634545
rect 263690 634471 263746 634480
rect 263704 520146 263732 634471
rect 282184 619676 282236 619682
rect 282184 619618 282236 619624
rect 282196 617574 282224 619618
rect 282184 617568 282236 617574
rect 282184 617510 282236 617516
rect 284206 611552 284262 611561
rect 284206 611487 284262 611496
rect 280804 556980 280856 556986
rect 280804 556922 280856 556928
rect 271144 555620 271196 555626
rect 271144 555562 271196 555568
rect 270774 551712 270830 551721
rect 270774 551647 270830 551656
rect 266726 548992 266782 549001
rect 266726 548927 266782 548936
rect 264242 547632 264298 547641
rect 264242 547567 264298 547576
rect 264256 522889 264284 547567
rect 265714 535120 265770 535129
rect 265714 535055 265770 535064
rect 264242 522880 264298 522889
rect 264242 522815 264298 522824
rect 264610 522064 264666 522073
rect 264666 522022 264744 522050
rect 264610 521999 264666 522008
rect 264716 520146 264744 522022
rect 265728 520146 265756 535055
rect 266740 520146 266768 548927
rect 270222 537840 270278 537849
rect 270222 537775 270278 537784
rect 267738 524240 267794 524249
rect 267738 524175 267794 524184
rect 267752 520146 267780 524175
rect 270236 522889 270264 537775
rect 269670 522880 269726 522889
rect 270222 522880 270278 522889
rect 269726 522838 269804 522866
rect 269670 522815 269726 522824
rect 268750 522200 268806 522209
rect 268750 522135 268806 522144
rect 269026 522200 269082 522209
rect 269026 522135 269082 522144
rect 268764 520146 268792 522135
rect 269040 521830 269068 522135
rect 269028 521824 269080 521830
rect 269028 521766 269080 521772
rect 269776 520146 269804 522838
rect 270222 522815 270278 522824
rect 270788 520146 270816 551647
rect 271156 522442 271184 555562
rect 277858 546272 277914 546281
rect 277858 546207 277914 546216
rect 274822 543416 274878 543425
rect 274822 543351 274878 543360
rect 272706 525600 272762 525609
rect 272762 525558 272840 525586
rect 272706 525535 272762 525544
rect 271602 522880 271658 522889
rect 271970 522880 272026 522889
rect 271658 522838 271828 522866
rect 271602 522815 271658 522824
rect 271144 522436 271196 522442
rect 271144 522378 271196 522384
rect 271800 520146 271828 522838
rect 271970 522815 272026 522824
rect 271984 522209 272012 522815
rect 271970 522200 272026 522209
rect 271970 522135 272026 522144
rect 272812 520146 272840 525558
rect 273810 525328 273866 525337
rect 273810 525263 273866 525272
rect 273824 520146 273852 525263
rect 274836 520146 274864 543351
rect 275834 542056 275890 542065
rect 275834 541991 275890 542000
rect 275848 520146 275876 541991
rect 276846 540696 276902 540705
rect 276846 540631 276902 540640
rect 276860 520146 276888 540631
rect 277872 520146 277900 546207
rect 278870 545048 278926 545057
rect 278870 544983 278926 544992
rect 278884 520146 278912 544983
rect 279882 536344 279938 536353
rect 279882 536279 279938 536288
rect 279896 520146 279924 536279
rect 280816 531146 280844 556922
rect 283930 550216 283986 550225
rect 283930 550151 283986 550160
rect 281906 549128 281962 549137
rect 281906 549063 281962 549072
rect 280804 531140 280856 531146
rect 280804 531082 280856 531088
rect 280710 523968 280766 523977
rect 280766 523926 280936 523954
rect 280710 523903 280766 523912
rect 280908 520146 280936 523926
rect 281920 520146 281948 549063
rect 282918 540968 282974 540977
rect 282918 540903 282974 540912
rect 282932 520146 282960 540903
rect 283944 520146 283972 550151
rect 284220 546553 284248 611487
rect 284942 551168 284998 551177
rect 284942 551103 284998 551112
rect 284206 546544 284262 546553
rect 284206 546479 284262 546488
rect 284956 520146 284984 551103
rect 285048 534993 285076 634743
rect 286324 603152 286376 603158
rect 286324 603094 286376 603100
rect 285954 543688 286010 543697
rect 285954 543623 286010 543632
rect 285034 534984 285090 534993
rect 285034 534919 285090 534928
rect 285772 530324 285824 530330
rect 285772 530266 285824 530272
rect 285680 529644 285732 529650
rect 285680 529586 285732 529592
rect 285692 528601 285720 529586
rect 285678 528592 285734 528601
rect 285678 528527 285734 528536
rect 285784 526454 285812 530266
rect 285772 526448 285824 526454
rect 285772 526390 285824 526396
rect 285680 524816 285732 524822
rect 285680 524758 285732 524764
rect 285692 521082 285720 524758
rect 285680 521076 285732 521082
rect 285680 521018 285732 521024
rect 285968 520146 285996 543623
rect 286336 526726 286364 603094
rect 286966 542328 287022 542337
rect 286966 542263 287022 542272
rect 286324 526720 286376 526726
rect 286324 526662 286376 526668
rect 286980 520146 287008 542263
rect 287716 526454 287744 636783
rect 289084 618316 289136 618322
rect 289084 618258 289136 618264
rect 288346 578232 288402 578241
rect 288346 578167 288402 578176
rect 287796 560312 287848 560318
rect 287796 560254 287848 560260
rect 287808 531214 287836 560254
rect 288360 550225 288388 578167
rect 288346 550216 288402 550225
rect 288346 550151 288402 550160
rect 288990 539336 289046 539345
rect 288990 539271 289046 539280
rect 287978 537296 288034 537305
rect 287978 537231 288034 537240
rect 287796 531208 287848 531214
rect 287796 531150 287848 531156
rect 287704 526448 287756 526454
rect 287704 526390 287756 526396
rect 287992 520146 288020 537231
rect 288346 526960 288402 526969
rect 288346 526895 288402 526904
rect 288360 526250 288388 526895
rect 288348 526244 288400 526250
rect 288348 526186 288400 526192
rect 288346 520704 288402 520713
rect 288346 520639 288402 520648
rect 288360 520606 288388 520639
rect 288348 520600 288400 520606
rect 288348 520542 288400 520548
rect 289004 520146 289032 539271
rect 289096 528494 289124 618258
rect 291106 585168 291162 585177
rect 291106 585103 291162 585112
rect 289174 581224 289230 581233
rect 289174 581159 289230 581168
rect 289188 555801 289216 581159
rect 290922 581088 290978 581097
rect 290922 581023 290978 581032
rect 289266 580000 289322 580009
rect 289266 579935 289322 579944
rect 289280 560289 289308 579935
rect 289726 570208 289782 570217
rect 289726 570143 289782 570152
rect 289450 568032 289506 568041
rect 289450 567967 289506 567976
rect 289266 560280 289322 560289
rect 289266 560215 289322 560224
rect 289464 556209 289492 567967
rect 289634 564496 289690 564505
rect 289634 564431 289690 564440
rect 289542 563136 289598 563145
rect 289542 563071 289598 563080
rect 289450 556200 289506 556209
rect 289450 556135 289506 556144
rect 289174 555792 289230 555801
rect 289174 555727 289230 555736
rect 289556 552809 289584 563071
rect 289542 552800 289598 552809
rect 289542 552735 289598 552744
rect 289648 546038 289676 564431
rect 289740 549137 289768 570143
rect 289726 549128 289782 549137
rect 289726 549063 289782 549072
rect 289636 546032 289688 546038
rect 289636 545974 289688 545980
rect 290002 545592 290058 545601
rect 290002 545527 290058 545536
rect 289084 528488 289136 528494
rect 289084 528430 289136 528436
rect 290016 520146 290044 545527
rect 290830 544232 290886 544241
rect 290830 544167 290886 544176
rect 290844 538214 290872 544167
rect 290936 539345 290964 581023
rect 291014 580952 291070 580961
rect 291014 580887 291070 580896
rect 291028 542201 291056 580887
rect 291014 542192 291070 542201
rect 291014 542127 291070 542136
rect 290922 539336 290978 539345
rect 290922 539271 290978 539280
rect 290844 538186 291056 538214
rect 291028 520146 291056 538186
rect 291120 524113 291148 585103
rect 291750 572384 291806 572393
rect 291750 572319 291806 572328
rect 291764 558521 291792 572319
rect 291750 558512 291806 558521
rect 291750 558447 291806 558456
rect 291856 541890 291884 638318
rect 292028 637016 292080 637022
rect 292028 636958 292080 636964
rect 291934 622432 291990 622441
rect 291934 622367 291990 622376
rect 291948 554305 291976 622367
rect 292040 612746 292068 636958
rect 294616 624889 294644 642087
rect 294800 625705 294828 642223
rect 295982 638752 296038 638761
rect 295982 638687 296038 638696
rect 294786 625696 294842 625705
rect 294786 625631 294842 625640
rect 294602 624880 294658 624889
rect 294602 624815 294658 624824
rect 293224 616888 293276 616894
rect 293224 616830 293276 616836
rect 292028 612740 292080 612746
rect 292028 612682 292080 612688
rect 292210 596592 292266 596601
rect 292210 596527 292266 596536
rect 292026 590880 292082 590889
rect 292026 590815 292082 590824
rect 292040 558793 292068 590815
rect 292118 586664 292174 586673
rect 292118 586599 292174 586608
rect 292026 558784 292082 558793
rect 292026 558719 292082 558728
rect 292132 554713 292160 586599
rect 292224 569265 292252 596527
rect 292394 583264 292450 583273
rect 292394 583199 292450 583208
rect 292210 569256 292266 569265
rect 292210 569191 292266 569200
rect 292302 566944 292358 566953
rect 292302 566879 292358 566888
rect 292210 558784 292266 558793
rect 292210 558719 292266 558728
rect 292118 554704 292174 554713
rect 292118 554639 292174 554648
rect 291934 554296 291990 554305
rect 291934 554231 291990 554240
rect 292026 547768 292082 547777
rect 292026 547703 292082 547712
rect 291844 541884 291896 541890
rect 291844 541826 291896 541832
rect 291106 524104 291162 524113
rect 291106 524039 291162 524048
rect 291842 521112 291898 521121
rect 291842 521047 291898 521056
rect 291856 520674 291884 521047
rect 291844 520668 291896 520674
rect 291844 520610 291896 520616
rect 292040 520146 292068 547703
rect 292224 533633 292252 558719
rect 292316 551721 292344 566879
rect 292408 558657 292436 583199
rect 292486 562320 292542 562329
rect 292486 562255 292542 562264
rect 292394 558648 292450 558657
rect 292394 558583 292450 558592
rect 292302 551712 292358 551721
rect 292302 551647 292358 551656
rect 292500 543697 292528 562255
rect 293236 557054 293264 616830
rect 295246 601080 295302 601089
rect 295246 601015 295302 601024
rect 294602 593056 294658 593065
rect 294602 592991 294658 593000
rect 293774 568576 293830 568585
rect 293774 568511 293830 568520
rect 293316 558408 293368 558414
rect 293316 558350 293368 558356
rect 293224 557048 293276 557054
rect 293224 556990 293276 556996
rect 292486 543688 292542 543697
rect 292486 543623 292542 543632
rect 293038 534576 293094 534585
rect 293038 534511 293094 534520
rect 292210 533624 292266 533633
rect 292210 533559 292266 533568
rect 293052 520146 293080 534511
rect 293328 521286 293356 558350
rect 293788 555801 293816 568511
rect 293866 565856 293922 565865
rect 293866 565791 293922 565800
rect 293774 555792 293830 555801
rect 293774 555727 293830 555736
rect 293880 546553 293908 565791
rect 294052 560924 294104 560930
rect 294052 560866 294104 560872
rect 293960 560720 294012 560726
rect 293960 560662 294012 560668
rect 293972 558482 294000 560662
rect 293960 558476 294012 558482
rect 293960 558418 294012 558424
rect 294064 558346 294092 560866
rect 294616 560153 294644 592991
rect 295154 590608 295210 590617
rect 295154 590543 295210 590552
rect 295062 589248 295118 589257
rect 295062 589183 295118 589192
rect 294970 586528 295026 586537
rect 294970 586463 295026 586472
rect 294878 569936 294934 569945
rect 294878 569871 294934 569880
rect 294602 560144 294658 560153
rect 294602 560079 294658 560088
rect 294052 558340 294104 558346
rect 294052 558282 294104 558288
rect 294892 552945 294920 569871
rect 294984 559881 295012 586463
rect 294970 559872 295026 559881
rect 294970 559807 295026 559816
rect 294878 552936 294934 552945
rect 294878 552871 294934 552880
rect 295076 547777 295104 589183
rect 295062 547768 295118 547777
rect 295062 547703 295118 547712
rect 293866 546544 293922 546553
rect 293866 546479 293922 546488
rect 295062 540152 295118 540161
rect 295062 540087 295118 540096
rect 294050 536480 294106 536489
rect 294050 536415 294106 536424
rect 293316 521280 293368 521286
rect 293316 521222 293368 521228
rect 294064 520146 294092 536415
rect 295076 520146 295104 540087
rect 295168 538665 295196 590543
rect 295154 538656 295210 538665
rect 295154 538591 295210 538600
rect 295260 535129 295288 601015
rect 295246 535120 295302 535129
rect 295246 535055 295302 535064
rect 295996 522345 296024 638687
rect 296166 636712 296222 636721
rect 296166 636647 296222 636656
rect 296074 550080 296130 550089
rect 296074 550015 296130 550024
rect 295982 522336 296038 522345
rect 295982 522271 296038 522280
rect 296088 520146 296116 550015
rect 296180 522209 296208 636647
rect 297284 633321 297312 643719
rect 297914 643512 297970 643521
rect 297914 643447 297970 643456
rect 297730 643376 297786 643385
rect 297730 643311 297786 643320
rect 297546 642696 297602 642705
rect 297546 642631 297602 642640
rect 297456 636948 297508 636954
rect 297456 636890 297508 636896
rect 297364 636880 297416 636886
rect 297364 636822 297416 636828
rect 297270 633312 297326 633321
rect 297270 633247 297326 633256
rect 297376 623529 297404 636822
rect 297362 623520 297418 623529
rect 297362 623455 297418 623464
rect 297362 621344 297418 621353
rect 297362 621279 297418 621288
rect 296626 597544 296682 597553
rect 296626 597479 296682 597488
rect 296534 596184 296590 596193
rect 296534 596119 296590 596128
rect 296548 587217 296576 596119
rect 296534 587208 296590 587217
rect 296534 587143 296590 587152
rect 296534 586392 296590 586401
rect 296534 586327 296590 586336
rect 296548 577425 296576 586327
rect 296534 577416 296590 577425
rect 296534 577351 296590 577360
rect 296534 576736 296590 576745
rect 296534 576671 296590 576680
rect 296548 567497 296576 576671
rect 296534 567488 296590 567497
rect 296534 567423 296590 567432
rect 296534 567080 296590 567089
rect 296534 567015 296590 567024
rect 296548 557841 296576 567015
rect 296534 557832 296590 557841
rect 296534 557767 296590 557776
rect 296534 557288 296590 557297
rect 296534 557223 296590 557232
rect 296548 550225 296576 557223
rect 296534 550216 296590 550225
rect 296534 550151 296590 550160
rect 296640 525473 296668 597479
rect 296718 587208 296774 587217
rect 296718 587143 296774 587152
rect 296732 586537 296760 587143
rect 296718 586528 296774 586537
rect 296718 586463 296774 586472
rect 297376 536654 297404 621279
rect 297468 617001 297496 636890
rect 297560 628969 297588 642631
rect 297638 640928 297694 640937
rect 297638 640863 297694 640872
rect 297546 628960 297602 628969
rect 297546 628895 297602 628904
rect 297652 627881 297680 640863
rect 297744 631145 297772 643311
rect 297822 635488 297878 635497
rect 297822 635423 297878 635432
rect 297730 631136 297786 631145
rect 297730 631071 297786 631080
rect 297638 627872 297694 627881
rect 297638 627807 297694 627816
rect 297836 626793 297864 635423
rect 297928 632233 297956 643447
rect 298098 642560 298154 642569
rect 298098 642495 298154 642504
rect 298006 640248 298062 640257
rect 298006 640183 298062 640192
rect 297914 632224 297970 632233
rect 297914 632159 297970 632168
rect 298020 630057 298048 640183
rect 298006 630048 298062 630057
rect 298006 629983 298062 629992
rect 297822 626784 297878 626793
rect 297822 626719 297878 626728
rect 298006 620256 298062 620265
rect 298006 620191 298062 620200
rect 298020 619682 298048 620191
rect 298008 619676 298060 619682
rect 298008 619618 298060 619624
rect 298006 619168 298062 619177
rect 298006 619103 298062 619112
rect 298020 618322 298048 619103
rect 298008 618316 298060 618322
rect 298008 618258 298060 618264
rect 298006 618080 298062 618089
rect 298006 618015 298062 618024
rect 297454 616992 297510 617001
rect 297454 616927 297510 616936
rect 298020 616894 298048 618015
rect 298008 616888 298060 616894
rect 298008 616830 298060 616836
rect 298006 613728 298062 613737
rect 297928 613686 298006 613714
rect 297546 609376 297602 609385
rect 297546 609311 297602 609320
rect 297454 608288 297510 608297
rect 297454 608223 297510 608232
rect 297468 551750 297496 608223
rect 297560 558550 297588 609311
rect 297638 606112 297694 606121
rect 297638 606047 297694 606056
rect 297652 560250 297680 606047
rect 297928 605834 297956 613686
rect 298006 613663 298062 613672
rect 298008 612740 298060 612746
rect 298008 612682 298060 612688
rect 298020 612649 298048 612682
rect 298006 612640 298062 612649
rect 298006 612575 298062 612584
rect 297928 605806 298048 605834
rect 297914 603936 297970 603945
rect 297914 603871 297970 603880
rect 297928 603158 297956 603871
rect 297916 603152 297968 603158
rect 297916 603094 297968 603100
rect 297730 569120 297786 569129
rect 297730 569055 297786 569064
rect 297640 560244 297692 560250
rect 297640 560186 297692 560192
rect 297548 558544 297600 558550
rect 297548 558486 297600 558492
rect 297744 557530 297772 569055
rect 297914 561368 297970 561377
rect 297914 561303 297970 561312
rect 297928 560930 297956 561303
rect 297916 560924 297968 560930
rect 297916 560866 297968 560872
rect 297732 557524 297784 557530
rect 297732 557466 297784 557472
rect 297456 551744 297508 551750
rect 297456 551686 297508 551692
rect 298020 542473 298048 605806
rect 298006 542464 298062 542473
rect 298006 542399 298062 542408
rect 297364 536648 297416 536654
rect 297364 536590 297416 536596
rect 298006 526280 298062 526289
rect 298006 526215 298062 526224
rect 296626 525464 296682 525473
rect 296626 525399 296682 525408
rect 296902 522336 296958 522345
rect 296958 522294 297128 522322
rect 296902 522271 296958 522280
rect 296166 522200 296222 522209
rect 296166 522135 296222 522144
rect 297100 520146 297128 522294
rect 298020 522073 298048 526215
rect 298006 522064 298062 522073
rect 298006 521999 298062 522008
rect 298112 520146 298140 642495
rect 304276 634545 304304 646478
rect 305288 634916 305316 653647
rect 324594 650312 324650 650321
rect 324594 650247 324650 650256
rect 314290 649360 314346 649369
rect 314290 649295 314346 649304
rect 309140 639600 309192 639606
rect 309140 639542 309192 639548
rect 310426 639568 310482 639577
rect 307850 639296 307906 639305
rect 307850 639231 307906 639240
rect 306564 636812 306616 636818
rect 306564 636754 306616 636760
rect 306576 634916 306604 636754
rect 307864 634916 307892 639231
rect 309152 634916 309180 639542
rect 310426 639503 310482 639512
rect 310440 634916 310468 639503
rect 313004 638308 313056 638314
rect 313004 638250 313056 638256
rect 311714 637800 311770 637809
rect 311714 637735 311770 637744
rect 311728 634916 311756 637735
rect 313016 634916 313044 638250
rect 314304 634916 314332 649295
rect 323306 642016 323362 642025
rect 323306 641951 323362 641960
rect 320732 640960 320784 640966
rect 320732 640902 320784 640908
rect 316866 640792 316922 640801
rect 316866 640727 316922 640736
rect 315578 640656 315634 640665
rect 315578 640591 315634 640600
rect 315592 634916 315620 640591
rect 316880 634916 316908 640727
rect 318156 639532 318208 639538
rect 318156 639474 318208 639480
rect 318168 634916 318196 639474
rect 319444 638104 319496 638110
rect 319444 638046 319496 638052
rect 319456 634916 319484 638046
rect 320744 634916 320772 640902
rect 322020 640892 322072 640898
rect 322020 640834 322072 640840
rect 322032 634916 322060 640834
rect 323320 634916 323348 641951
rect 324608 634916 324636 650247
rect 345202 649632 345258 649641
rect 345202 649567 345258 649576
rect 334898 649224 334954 649233
rect 334898 649159 334954 649168
rect 332322 648952 332378 648961
rect 332322 648887 332378 648896
rect 327170 648000 327226 648009
rect 327170 647935 327226 647944
rect 325884 646196 325936 646202
rect 325884 646138 325936 646144
rect 325896 634916 325924 646138
rect 327184 634916 327212 647935
rect 329746 647592 329802 647601
rect 329746 647527 329802 647536
rect 328458 643240 328514 643249
rect 328458 643175 328514 643184
rect 328472 634916 328500 643175
rect 329760 634916 329788 647527
rect 331036 640824 331088 640830
rect 331036 640766 331088 640772
rect 331048 634916 331076 640766
rect 332336 634916 332364 648887
rect 333610 647864 333666 647873
rect 333610 647799 333666 647808
rect 333624 634916 333652 647799
rect 334912 634916 334940 649159
rect 343914 649088 343970 649097
rect 343914 649023 343970 649032
rect 336186 647728 336242 647737
rect 336186 647663 336242 647672
rect 336200 634916 336228 647663
rect 341338 647456 341394 647465
rect 341338 647391 341394 647400
rect 338764 643476 338816 643482
rect 338764 643418 338816 643424
rect 337476 640620 337528 640626
rect 337476 640562 337528 640568
rect 337488 634916 337516 640562
rect 338776 634916 338804 643418
rect 340052 642456 340104 642462
rect 340052 642398 340104 642404
rect 340064 634916 340092 642398
rect 341352 634916 341380 647391
rect 342628 635384 342680 635390
rect 342628 635326 342680 635332
rect 342640 634916 342668 635326
rect 343928 634916 343956 649023
rect 345216 634916 345244 649567
rect 347778 648816 347834 648825
rect 347778 648751 347834 648760
rect 346492 642320 346544 642326
rect 346492 642262 346544 642268
rect 346504 634916 346532 642262
rect 347792 634916 347820 648751
rect 354220 647556 354272 647562
rect 354220 647498 354272 647504
rect 351644 644496 351696 644502
rect 351644 644438 351696 644444
rect 350356 641980 350408 641986
rect 350356 641922 350408 641928
rect 349068 640484 349120 640490
rect 349068 640426 349120 640432
rect 349080 634916 349108 640426
rect 350368 634916 350396 641922
rect 351656 634916 351684 644438
rect 352932 641844 352984 641850
rect 352932 641786 352984 641792
rect 352944 634916 352972 641786
rect 354232 634916 354260 647498
rect 355508 641776 355560 641782
rect 355508 641718 355560 641724
rect 355520 634916 355548 641718
rect 356808 634916 356836 654463
rect 358082 654392 358138 654401
rect 358082 654327 358138 654336
rect 358096 634916 358124 654327
rect 359384 634916 359412 654599
rect 363234 654256 363290 654265
rect 363234 654191 363290 654200
rect 360658 653032 360714 653041
rect 360658 652967 360714 652976
rect 360672 634916 360700 652967
rect 361948 651568 362000 651574
rect 361948 651510 362000 651516
rect 361960 634916 361988 651510
rect 363248 634916 363276 654191
rect 364522 652896 364578 652905
rect 364522 652831 364578 652840
rect 364536 634916 364564 652831
rect 366376 647222 366404 654774
rect 368388 654152 368440 654158
rect 368388 654094 368440 654100
rect 366364 647216 366416 647222
rect 366364 647158 366416 647164
rect 365812 643340 365864 643346
rect 365812 643282 365864 643288
rect 365824 634916 365852 643282
rect 367100 637832 367152 637838
rect 367100 637774 367152 637780
rect 367112 634916 367140 637774
rect 368400 634916 368428 654094
rect 371896 652050 371924 656814
rect 371884 652044 371936 652050
rect 371884 651986 371936 651992
rect 377404 652044 377456 652050
rect 377404 651986 377456 651992
rect 374368 650344 374420 650350
rect 374368 650286 374420 650292
rect 372252 647284 372304 647290
rect 372252 647226 372304 647232
rect 371884 647216 371936 647222
rect 371884 647158 371936 647164
rect 370962 641064 371018 641073
rect 370962 640999 371018 641008
rect 369674 640384 369730 640393
rect 369674 640319 369730 640328
rect 369688 636313 369716 640319
rect 369674 636304 369730 636313
rect 369674 636239 369730 636248
rect 369688 634916 369716 636239
rect 370976 634916 371004 640999
rect 304262 634536 304318 634545
rect 304262 634471 304318 634480
rect 371896 634438 371924 647158
rect 372264 634916 372292 647226
rect 371884 634432 371936 634438
rect 299662 634400 299718 634409
rect 299662 634335 299718 634344
rect 302698 634400 302754 634409
rect 371884 634374 371936 634380
rect 302698 634335 302754 634344
rect 299676 634001 299704 634335
rect 303977 634208 303986 634264
rect 304042 634208 304051 634264
rect 299662 633992 299718 634001
rect 299662 633927 299718 633936
rect 374380 625154 374408 650286
rect 375656 650276 375708 650282
rect 375656 650218 375708 650224
rect 374828 650208 374880 650214
rect 374828 650150 374880 650156
rect 374552 650140 374604 650146
rect 374552 650082 374604 650088
rect 374458 636304 374514 636313
rect 374458 636239 374514 636248
rect 374472 632641 374500 636239
rect 374458 632632 374514 632641
rect 374458 632567 374514 632576
rect 374380 625126 374500 625154
rect 374472 623665 374500 625126
rect 374564 625025 374592 650082
rect 374736 650072 374788 650078
rect 374736 650014 374788 650020
rect 374748 626249 374776 650014
rect 374734 626240 374790 626249
rect 374734 626175 374790 626184
rect 374550 625016 374606 625025
rect 374550 624951 374606 624960
rect 374840 624617 374868 650150
rect 375564 642252 375616 642258
rect 375564 642194 375616 642200
rect 375470 639840 375526 639849
rect 375470 639775 375526 639784
rect 375380 635520 375432 635526
rect 375380 635462 375432 635468
rect 374826 624608 374882 624617
rect 374826 624543 374882 624552
rect 374458 623656 374514 623665
rect 374458 623591 374514 623600
rect 374642 618488 374698 618497
rect 374642 618423 374698 618432
rect 374550 614000 374606 614009
rect 374550 613935 374606 613944
rect 374458 612096 374514 612105
rect 374458 612031 374514 612040
rect 299846 604480 299902 604489
rect 299846 604415 299902 604424
rect 299754 602984 299810 602993
rect 299754 602919 299810 602928
rect 299386 601896 299442 601905
rect 299386 601831 299442 601840
rect 299202 594824 299258 594833
rect 299202 594759 299258 594768
rect 299110 571160 299166 571169
rect 299110 571095 299166 571104
rect 299018 561776 299074 561785
rect 299018 561711 299074 561720
rect 298742 560552 298798 560561
rect 298742 560487 298798 560496
rect 298756 540705 298784 560487
rect 299032 560289 299060 561711
rect 299018 560280 299074 560289
rect 299018 560215 299074 560224
rect 299124 551177 299152 571095
rect 299110 551168 299166 551177
rect 299110 551103 299166 551112
rect 299216 543833 299244 594759
rect 299294 592104 299350 592113
rect 299294 592039 299350 592048
rect 299202 543824 299258 543833
rect 299202 543759 299258 543768
rect 299202 543688 299258 543697
rect 299202 543623 299258 543632
rect 299216 542638 299244 543623
rect 299204 542632 299256 542638
rect 299204 542574 299256 542580
rect 298742 540696 298798 540705
rect 298742 540631 298798 540640
rect 299308 537010 299336 592039
rect 299124 536982 299336 537010
rect 299124 528554 299152 536982
rect 299400 536874 299428 601831
rect 299664 561740 299716 561746
rect 299664 561682 299716 561688
rect 299572 561196 299624 561202
rect 299572 561138 299624 561144
rect 299584 560998 299612 561138
rect 299572 560992 299624 560998
rect 299572 560934 299624 560940
rect 299572 560448 299624 560454
rect 299572 560390 299624 560396
rect 299584 557534 299612 560390
rect 299676 560114 299704 561682
rect 299664 560108 299716 560114
rect 299664 560050 299716 560056
rect 299584 557506 299704 557534
rect 299676 546106 299704 557506
rect 299768 552537 299796 602919
rect 299754 552528 299810 552537
rect 299754 552463 299810 552472
rect 299664 546100 299716 546106
rect 299664 546042 299716 546048
rect 299308 536846 299428 536874
rect 299308 529417 299336 536846
rect 299386 536752 299442 536761
rect 299386 536687 299442 536696
rect 299400 535838 299428 536687
rect 299388 535832 299440 535838
rect 299388 535774 299440 535780
rect 299860 534585 299888 604415
rect 299938 597544 299994 597553
rect 299938 597479 299994 597488
rect 299846 534576 299902 534585
rect 299846 534511 299902 534520
rect 299386 529816 299442 529825
rect 299386 529751 299442 529760
rect 299294 529408 299350 529417
rect 299294 529343 299350 529352
rect 299400 528834 299428 529751
rect 299388 528828 299440 528834
rect 299388 528770 299440 528776
rect 299124 528526 299336 528554
rect 299308 528290 299336 528526
rect 299296 528284 299348 528290
rect 299296 528226 299348 528232
rect 299952 523433 299980 597479
rect 319364 560658 319746 560674
rect 319352 560652 319746 560658
rect 319404 560646 319746 560652
rect 319352 560594 319404 560600
rect 300584 560584 300636 560590
rect 300584 560526 300636 560532
rect 302238 560552 302294 560561
rect 300596 558346 300624 560526
rect 300676 560516 300728 560522
rect 302294 560510 302542 560538
rect 302238 560487 302294 560496
rect 300676 560458 300728 560464
rect 300688 558550 300716 560458
rect 305550 560280 305606 560289
rect 315408 560250 315698 560266
rect 305550 560215 305606 560224
rect 315396 560244 315698 560250
rect 315448 560238 315698 560244
rect 315396 560186 315448 560192
rect 318340 560176 318392 560182
rect 300676 558544 300728 558550
rect 300676 558486 300728 558492
rect 300584 558340 300636 558346
rect 300584 558282 300636 558288
rect 301516 536586 301544 560116
rect 303540 558414 303568 560116
rect 303528 558408 303580 558414
rect 303528 558350 303580 558356
rect 304552 550390 304580 560116
rect 306392 560114 306590 560130
rect 318392 560124 318734 560130
rect 318340 560118 318734 560124
rect 306380 560108 306590 560114
rect 306432 560102 306590 560108
rect 306380 560050 306432 560056
rect 307206 553208 307262 553217
rect 307206 553143 307262 553152
rect 304540 550384 304592 550390
rect 304540 550326 304592 550332
rect 301504 536580 301556 536586
rect 301504 536522 301556 536528
rect 306194 529680 306250 529689
rect 306194 529615 306250 529624
rect 305182 529000 305238 529009
rect 305182 528935 305238 528944
rect 302238 528864 302294 528873
rect 302238 528799 302294 528808
rect 299938 523424 299994 523433
rect 299938 523359 299994 523368
rect 302252 522345 302280 528799
rect 302238 522336 302294 522345
rect 302238 522271 302294 522280
rect 304078 522336 304134 522345
rect 304134 522294 304212 522322
rect 304078 522271 304134 522280
rect 303066 522200 303122 522209
rect 303618 522200 303674 522209
rect 303122 522158 303200 522186
rect 303066 522135 303122 522144
rect 301134 521656 301190 521665
rect 301134 521591 301190 521600
rect 300030 521520 300086 521529
rect 300086 521478 300164 521506
rect 300030 521455 300086 521464
rect 299018 521384 299074 521393
rect 299074 521342 299152 521370
rect 299018 521319 299074 521328
rect 299124 520146 299152 521342
rect 300136 520146 300164 521478
rect 301148 520146 301176 521591
rect 302054 520840 302110 520849
rect 302110 520798 302188 520826
rect 302054 520775 302110 520784
rect 302160 520146 302188 520798
rect 303172 520146 303200 522158
rect 303618 522135 303674 522144
rect 303632 521898 303660 522135
rect 303620 521892 303672 521898
rect 303620 521834 303672 521840
rect 304184 520146 304212 522294
rect 305196 520146 305224 528935
rect 306208 520146 306236 529615
rect 307220 520146 307248 553143
rect 307588 546174 307616 560116
rect 308218 553072 308274 553081
rect 308218 553007 308274 553016
rect 307576 546168 307628 546174
rect 307576 546110 307628 546116
rect 308232 520146 308260 553007
rect 308600 525434 308628 560116
rect 309230 550352 309286 550361
rect 309230 550287 309286 550296
rect 308588 525428 308640 525434
rect 308588 525370 308640 525376
rect 309244 520146 309272 550287
rect 309612 535294 309640 560116
rect 309600 535288 309652 535294
rect 309600 535230 309652 535236
rect 310242 535256 310298 535265
rect 310242 535191 310298 535200
rect 310256 520146 310284 535191
rect 310624 530777 310652 560116
rect 311254 538520 311310 538529
rect 311254 538455 311310 538464
rect 310610 530768 310666 530777
rect 310610 530703 310666 530712
rect 311268 520146 311296 538455
rect 311636 538082 311664 560116
rect 311624 538076 311676 538082
rect 311624 538018 311676 538024
rect 312174 527776 312230 527785
rect 312230 527734 312308 527762
rect 312174 527711 312230 527720
rect 312280 520146 312308 527734
rect 312648 521354 312676 560116
rect 313660 546242 313688 560116
rect 314672 558550 314700 560116
rect 314660 558544 314712 558550
rect 314660 558486 314712 558492
rect 313922 555928 313978 555937
rect 313922 555863 313978 555872
rect 313648 546236 313700 546242
rect 313648 546178 313700 546184
rect 313936 538214 313964 555863
rect 316696 542162 316724 560116
rect 317708 551818 317736 560116
rect 318352 560102 318734 560118
rect 317696 551812 317748 551818
rect 317696 551754 317748 551760
rect 320362 549264 320418 549273
rect 320362 549199 320418 549208
rect 316684 542156 316736 542162
rect 316684 542098 316736 542104
rect 316314 540832 316370 540841
rect 316314 540767 316370 540776
rect 313936 538186 314056 538214
rect 313188 530528 313240 530534
rect 313188 530470 313240 530476
rect 313200 522578 313228 530470
rect 313370 523152 313426 523161
rect 313370 523087 313426 523096
rect 313278 523016 313334 523025
rect 313278 522951 313334 522960
rect 313188 522572 313240 522578
rect 313188 522514 313240 522520
rect 313292 521694 313320 522951
rect 313280 521688 313332 521694
rect 313280 521630 313332 521636
rect 312636 521348 312688 521354
rect 312636 521290 312688 521296
rect 313384 520146 313412 523087
rect 314028 522345 314056 538186
rect 315302 533896 315358 533905
rect 315302 533831 315358 533840
rect 314014 522336 314070 522345
rect 314014 522271 314070 522280
rect 314290 522064 314346 522073
rect 314290 521999 314346 522008
rect 226260 520118 226304 520146
rect 227272 520118 227316 520146
rect 228284 520118 228328 520146
rect 229296 520118 229340 520146
rect 230308 520118 230352 520146
rect 231320 520118 231364 520146
rect 232332 520118 232376 520146
rect 233344 520118 233388 520146
rect 234356 520118 234400 520146
rect 235368 520118 235412 520146
rect 236380 520118 236424 520146
rect 237392 520118 237436 520146
rect 238404 520118 238448 520146
rect 239416 520118 239460 520146
rect 240428 520118 240472 520146
rect 241440 520118 241484 520146
rect 242452 520118 242496 520146
rect 243464 520118 243508 520146
rect 244476 520118 244520 520146
rect 245488 520118 245532 520146
rect 246500 520118 246544 520146
rect 247512 520118 247556 520146
rect 248524 520118 248568 520146
rect 249536 520118 249580 520146
rect 250548 520118 250592 520146
rect 251560 520118 251604 520146
rect 252572 520118 252616 520146
rect 253584 520118 253628 520146
rect 254596 520118 254640 520146
rect 255608 520118 255652 520146
rect 256620 520118 256664 520146
rect 257632 520118 257676 520146
rect 258644 520118 258688 520146
rect 259656 520118 259700 520146
rect 260668 520118 260712 520146
rect 261680 520118 261724 520146
rect 262692 520118 262736 520146
rect 263704 520118 263748 520146
rect 264716 520118 264760 520146
rect 265728 520118 265772 520146
rect 266740 520118 266784 520146
rect 267752 520118 267796 520146
rect 268764 520118 268808 520146
rect 269776 520118 269820 520146
rect 270788 520118 270832 520146
rect 271800 520118 271844 520146
rect 272812 520118 272856 520146
rect 273824 520118 273868 520146
rect 274836 520118 274880 520146
rect 275848 520118 275892 520146
rect 276860 520118 276904 520146
rect 277872 520118 277916 520146
rect 278884 520118 278928 520146
rect 279896 520118 279940 520146
rect 280908 520118 280952 520146
rect 281920 520118 281964 520146
rect 282932 520118 282976 520146
rect 283944 520118 283988 520146
rect 284956 520118 285000 520146
rect 285968 520118 286012 520146
rect 286980 520118 287024 520146
rect 287992 520118 288036 520146
rect 289004 520118 289048 520146
rect 290016 520118 290060 520146
rect 291028 520118 291072 520146
rect 292040 520118 292084 520146
rect 293052 520118 293096 520146
rect 294064 520118 294108 520146
rect 295076 520118 295120 520146
rect 296088 520118 296132 520146
rect 297100 520118 297144 520146
rect 298112 520118 298156 520146
rect 299124 520118 299168 520146
rect 300136 520118 300180 520146
rect 301148 520118 301192 520146
rect 302160 520118 302204 520146
rect 303172 520118 303216 520146
rect 304184 520118 304228 520146
rect 305196 520118 305240 520146
rect 306208 520118 306252 520146
rect 307220 520118 307264 520146
rect 308232 520118 308276 520146
rect 309244 520118 309288 520146
rect 310256 520118 310300 520146
rect 311268 520118 311312 520146
rect 312280 520118 312324 520146
rect 225264 519860 225292 520118
rect 226276 519860 226304 520118
rect 227288 519860 227316 520118
rect 228300 519860 228328 520118
rect 229312 519860 229340 520118
rect 230324 519860 230352 520118
rect 231336 519860 231364 520118
rect 232348 519860 232376 520118
rect 233360 519860 233388 520118
rect 234372 519860 234400 520118
rect 235384 519860 235412 520118
rect 236396 519860 236424 520118
rect 237408 519860 237436 520118
rect 238420 519860 238448 520118
rect 239432 519860 239460 520118
rect 240444 519860 240472 520118
rect 241456 519860 241484 520118
rect 242468 519860 242496 520118
rect 243480 519860 243508 520118
rect 244492 519860 244520 520118
rect 245504 519860 245532 520118
rect 246516 519860 246544 520118
rect 247528 519860 247556 520118
rect 248540 519860 248568 520118
rect 249552 519860 249580 520118
rect 250564 519860 250592 520118
rect 251576 519860 251604 520118
rect 252588 519860 252616 520118
rect 253600 519860 253628 520118
rect 254612 519860 254640 520118
rect 255624 519860 255652 520118
rect 256636 519860 256664 520118
rect 257648 519860 257676 520118
rect 258660 519860 258688 520118
rect 259672 519860 259700 520118
rect 260684 519860 260712 520118
rect 261696 519860 261724 520118
rect 262708 519860 262736 520118
rect 263720 519860 263748 520118
rect 264732 519860 264760 520118
rect 265744 519860 265772 520118
rect 266756 519860 266784 520118
rect 267768 519860 267796 520118
rect 268780 519860 268808 520118
rect 269792 519860 269820 520118
rect 270804 519860 270832 520118
rect 271816 519860 271844 520118
rect 272828 519860 272856 520118
rect 273840 519860 273868 520118
rect 274852 519860 274880 520118
rect 275864 519860 275892 520118
rect 276876 519860 276904 520118
rect 277888 519860 277916 520118
rect 278900 519860 278928 520118
rect 279912 519860 279940 520118
rect 280924 519860 280952 520118
rect 281936 519860 281964 520118
rect 282948 519860 282976 520118
rect 283960 519860 283988 520118
rect 284972 519860 285000 520118
rect 285984 519860 286012 520118
rect 286996 519860 287024 520118
rect 288008 519860 288036 520118
rect 289020 519860 289048 520118
rect 290032 519860 290060 520118
rect 291044 519860 291072 520118
rect 292056 519860 292084 520118
rect 293068 519860 293096 520118
rect 294080 519860 294108 520118
rect 295092 519860 295120 520118
rect 296104 519860 296132 520118
rect 297116 519860 297144 520118
rect 298128 519860 298156 520118
rect 299140 519860 299168 520118
rect 300152 519860 300180 520118
rect 301164 519860 301192 520118
rect 302176 519860 302204 520118
rect 303188 519860 303216 520118
rect 304200 519860 304228 520118
rect 305212 519860 305240 520118
rect 306224 519860 306252 520118
rect 307236 519860 307264 520118
rect 308248 519860 308276 520118
rect 309260 519860 309288 520118
rect 310272 519860 310300 520118
rect 311284 519860 311312 520118
rect 312296 519860 312324 520118
rect 313308 520118 313412 520146
rect 314304 520146 314332 521999
rect 315316 520146 315344 533831
rect 316328 520146 316356 540767
rect 319350 537976 319406 537985
rect 319350 537911 319406 537920
rect 318338 535936 318394 535945
rect 318338 535871 318394 535880
rect 317326 535392 317382 535401
rect 317326 535327 317382 535336
rect 317340 520146 317368 535327
rect 318352 520146 318380 535871
rect 319364 520146 319392 537911
rect 320376 520146 320404 549199
rect 320744 547738 320772 560116
rect 321374 551984 321430 551993
rect 321374 551919 321430 551928
rect 320732 547732 320784 547738
rect 320732 547674 320784 547680
rect 321388 520146 321416 551919
rect 321756 529718 321784 560116
rect 322768 558793 322796 560116
rect 322754 558784 322810 558793
rect 322754 558719 322810 558728
rect 323780 554674 323808 560116
rect 323768 554668 323820 554674
rect 323768 554610 323820 554616
rect 323398 552392 323454 552401
rect 323398 552327 323454 552336
rect 321744 529712 321796 529718
rect 321744 529654 321796 529660
rect 322386 527096 322442 527105
rect 322386 527031 322442 527040
rect 322400 520146 322428 527031
rect 323412 520146 323440 552327
rect 324792 544950 324820 560116
rect 324780 544944 324832 544950
rect 324780 544886 324832 544892
rect 325804 543590 325832 560116
rect 326816 553178 326844 560116
rect 326804 553172 326856 553178
rect 326804 553114 326856 553120
rect 327828 550526 327856 560116
rect 328458 551848 328514 551857
rect 328458 551783 328514 551792
rect 327816 550520 327868 550526
rect 327816 550462 327868 550468
rect 325792 543584 325844 543590
rect 325792 543526 325844 543532
rect 325422 537160 325478 537169
rect 325422 537095 325478 537104
rect 324410 534032 324466 534041
rect 324410 533967 324466 533976
rect 324424 520146 324452 533967
rect 325436 520146 325464 537095
rect 326434 535800 326490 535809
rect 326434 535735 326490 535744
rect 326448 520146 326476 535735
rect 327354 524784 327410 524793
rect 327410 524742 327488 524770
rect 327354 524719 327410 524728
rect 327460 520146 327488 524742
rect 328472 520146 328500 551783
rect 328840 542230 328868 560116
rect 329852 545018 329880 560116
rect 329840 545012 329892 545018
rect 329840 544954 329892 544960
rect 328828 542224 328880 542230
rect 328828 542166 328880 542172
rect 330864 538150 330892 560116
rect 331876 539374 331904 560116
rect 331956 556912 332008 556918
rect 331956 556854 332008 556860
rect 331864 539368 331916 539374
rect 331864 539310 331916 539316
rect 330852 538144 330904 538150
rect 330852 538086 330904 538092
rect 331494 528456 331550 528465
rect 331494 528391 331550 528400
rect 330390 528048 330446 528057
rect 330446 528006 330524 528034
rect 330390 527983 330446 527992
rect 329378 527912 329434 527921
rect 329434 527870 329512 527898
rect 329378 527847 329434 527856
rect 329484 520146 329512 527870
rect 330496 520146 330524 528006
rect 331508 520146 331536 528391
rect 331968 522170 331996 556854
rect 332888 534002 332916 560116
rect 332876 533996 332928 534002
rect 332876 533938 332928 533944
rect 333900 529786 333928 560116
rect 334912 535362 334940 560116
rect 335924 546310 335952 560116
rect 336936 552673 336964 560116
rect 336922 552664 336978 552673
rect 336922 552599 336978 552608
rect 335912 546304 335964 546310
rect 335912 546246 335964 546252
rect 335542 545456 335598 545465
rect 335542 545391 335598 545400
rect 334900 535356 334952 535362
rect 334900 535298 334952 535304
rect 333888 529780 333940 529786
rect 333888 529722 333940 529728
rect 332322 528320 332378 528329
rect 332378 528278 332548 528306
rect 332322 528255 332378 528264
rect 331956 522164 332008 522170
rect 331956 522106 332008 522112
rect 332520 520146 332548 528278
rect 334530 527640 334586 527649
rect 334530 527575 334586 527584
rect 333426 527368 333482 527377
rect 333482 527326 333560 527354
rect 333426 527303 333482 527312
rect 333532 520146 333560 527326
rect 334544 520146 334572 527575
rect 335556 520146 335584 545391
rect 336554 543552 336610 543561
rect 336554 543487 336610 543496
rect 336568 520146 336596 543487
rect 337948 533866 337976 560116
rect 338578 541512 338634 541521
rect 338578 541447 338634 541456
rect 337936 533860 337988 533866
rect 337936 533802 337988 533808
rect 337476 522504 337528 522510
rect 337476 522446 337528 522452
rect 337488 520146 337516 522446
rect 338592 520146 338620 541447
rect 338960 521490 338988 560116
rect 339972 533934 340000 560116
rect 340602 550488 340658 550497
rect 340602 550423 340658 550432
rect 339960 533928 340012 533934
rect 339960 533870 340012 533876
rect 339498 522472 339554 522481
rect 339554 522430 339632 522458
rect 339498 522407 339554 522416
rect 338948 521484 339000 521490
rect 338948 521426 339000 521432
rect 339604 520146 339632 522430
rect 340616 520146 340644 550423
rect 340984 539442 341012 560116
rect 341614 544912 341670 544921
rect 341614 544847 341670 544856
rect 340972 539436 341024 539442
rect 340972 539378 341024 539384
rect 341628 520146 341656 544847
rect 341996 527066 342024 560116
rect 343008 536722 343036 560116
rect 343640 552288 343692 552294
rect 343640 552230 343692 552236
rect 342996 536716 343048 536722
rect 342996 536658 343048 536664
rect 342904 530596 342956 530602
rect 342904 530538 342956 530544
rect 342628 528216 342680 528222
rect 342628 528158 342680 528164
rect 341984 527060 342036 527066
rect 341984 527002 342036 527008
rect 342640 520146 342668 528158
rect 342916 522510 342944 530538
rect 342904 522504 342956 522510
rect 342904 522446 342956 522452
rect 343652 520146 343680 552230
rect 344020 550594 344048 560116
rect 344652 552220 344704 552226
rect 344652 552162 344704 552168
rect 344008 550588 344060 550594
rect 344008 550530 344060 550536
rect 344664 520146 344692 552162
rect 345032 540870 345060 560116
rect 345662 554024 345718 554033
rect 345662 553959 345718 553968
rect 345020 540864 345072 540870
rect 345020 540806 345072 540812
rect 345676 520146 345704 553959
rect 346044 552022 346072 560116
rect 346676 557728 346728 557734
rect 346676 557670 346728 557676
rect 346032 552016 346084 552022
rect 346032 551958 346084 551964
rect 346688 520146 346716 557670
rect 347056 547874 347084 560116
rect 347136 555552 347188 555558
rect 347136 555494 347188 555500
rect 347044 547868 347096 547874
rect 347044 547810 347096 547816
rect 347148 522646 347176 555494
rect 348068 549030 348096 560116
rect 348056 549024 348108 549030
rect 348056 548966 348108 548972
rect 348700 534948 348752 534954
rect 348700 534890 348752 534896
rect 347686 529272 347742 529281
rect 347686 529207 347742 529216
rect 347136 522640 347188 522646
rect 347136 522582 347188 522588
rect 347700 520146 347728 529207
rect 348712 520146 348740 534890
rect 349080 525094 349108 560116
rect 350092 546378 350120 560116
rect 350080 546372 350132 546378
rect 350080 546314 350132 546320
rect 350722 544504 350778 544513
rect 350722 544439 350778 544448
rect 349710 543008 349766 543017
rect 349710 542943 349766 542952
rect 349068 525088 349120 525094
rect 349068 525030 349120 525036
rect 349724 520146 349752 542943
rect 350538 542872 350594 542881
rect 350538 542807 350594 542816
rect 350552 539481 350580 542807
rect 350538 539472 350594 539481
rect 350538 539407 350594 539416
rect 350736 520146 350764 544439
rect 351104 524210 351132 560116
rect 351736 552152 351788 552158
rect 351736 552094 351788 552100
rect 351092 524204 351144 524210
rect 351092 524146 351144 524152
rect 351748 520146 351776 552094
rect 352116 539510 352144 560116
rect 353128 558482 353156 560116
rect 353116 558476 353168 558482
rect 353116 558418 353168 558424
rect 354140 549166 354168 560116
rect 355152 558618 355180 560116
rect 355140 558612 355192 558618
rect 355140 558554 355192 558560
rect 354128 549160 354180 549166
rect 354128 549102 354180 549108
rect 354772 539912 354824 539918
rect 354772 539854 354824 539860
rect 352104 539504 352156 539510
rect 352104 539446 352156 539452
rect 352746 538928 352802 538937
rect 352746 538863 352802 538872
rect 352760 520146 352788 538863
rect 353760 535832 353812 535838
rect 353760 535774 353812 535780
rect 353772 520146 353800 535774
rect 354784 520146 354812 539854
rect 355784 535764 355836 535770
rect 355784 535706 355836 535712
rect 355796 520146 355824 535706
rect 356164 523734 356192 560116
rect 357176 558686 357204 560116
rect 357808 559632 357860 559638
rect 357808 559574 357860 559580
rect 357164 558680 357216 558686
rect 357164 558622 357216 558628
rect 356794 532536 356850 532545
rect 356794 532471 356850 532480
rect 356152 523728 356204 523734
rect 356152 523670 356204 523676
rect 356808 520146 356836 532471
rect 357820 520146 357848 559574
rect 358188 535430 358216 560116
rect 358818 548584 358874 548593
rect 358818 548519 358874 548528
rect 358176 535424 358228 535430
rect 358176 535366 358228 535372
rect 358832 520146 358860 548519
rect 359200 546446 359228 560116
rect 359830 547088 359886 547097
rect 359830 547023 359886 547032
rect 359188 546440 359240 546446
rect 359188 546382 359240 546388
rect 359844 520146 359872 547023
rect 360212 543658 360240 560116
rect 361224 558754 361252 560116
rect 361212 558748 361264 558754
rect 361212 558690 361264 558696
rect 360844 550860 360896 550866
rect 360844 550802 360896 550808
rect 360200 543652 360252 543658
rect 360200 543594 360252 543600
rect 360856 520146 360884 550802
rect 362236 543726 362264 560116
rect 362866 545864 362922 545873
rect 362866 545799 362922 545808
rect 362224 543720 362276 543726
rect 362224 543662 362276 543668
rect 361854 522608 361910 522617
rect 361854 522543 361910 522552
rect 361868 520146 361896 522543
rect 362880 520146 362908 545799
rect 363248 542366 363276 560116
rect 364260 545086 364288 560116
rect 364248 545080 364300 545086
rect 364248 545022 364300 545028
rect 363236 542360 363288 542366
rect 363236 542302 363288 542308
rect 363878 529136 363934 529145
rect 363878 529071 363934 529080
rect 363892 520146 363920 529071
rect 364892 528828 364944 528834
rect 364892 528770 364944 528776
rect 364904 520146 364932 528770
rect 365272 527134 365300 560116
rect 365904 546848 365956 546854
rect 365904 546790 365956 546796
rect 365260 527128 365312 527134
rect 365260 527070 365312 527076
rect 365916 520146 365944 546790
rect 366284 534070 366312 560116
rect 367296 558822 367324 560116
rect 367928 559496 367980 559502
rect 367928 559438 367980 559444
rect 367284 558816 367336 558822
rect 367284 558758 367336 558764
rect 366914 544368 366970 544377
rect 366914 544303 366970 544312
rect 366272 534064 366324 534070
rect 366272 534006 366324 534012
rect 366928 520146 366956 544303
rect 367940 520146 367968 559438
rect 368308 540938 368336 560116
rect 368940 559428 368992 559434
rect 368940 559370 368992 559376
rect 368296 540932 368348 540938
rect 368296 540874 368348 540880
rect 368952 520146 368980 559370
rect 369320 553314 369348 560116
rect 369952 559292 370004 559298
rect 369952 559234 370004 559240
rect 369308 553308 369360 553314
rect 369308 553250 369360 553256
rect 369124 522912 369176 522918
rect 369124 522854 369176 522860
rect 369136 522102 369164 522854
rect 369124 522096 369176 522102
rect 369124 522038 369176 522044
rect 369964 520146 369992 559234
rect 370332 536790 370360 560116
rect 370964 559224 371016 559230
rect 370964 559166 371016 559172
rect 370320 536784 370372 536790
rect 370320 536726 370372 536732
rect 370976 520146 371004 559166
rect 371344 539578 371372 560116
rect 371976 559156 372028 559162
rect 371976 559098 372028 559104
rect 371332 539572 371384 539578
rect 371332 539514 371384 539520
rect 371988 520146 372016 559098
rect 372356 558890 372384 560116
rect 373264 559088 373316 559094
rect 373264 559030 373316 559036
rect 372344 558884 372396 558890
rect 372344 558826 372396 558832
rect 372988 549432 373040 549438
rect 372988 549374 373040 549380
rect 373000 520146 373028 549374
rect 373276 522918 373304 559030
rect 373368 538218 373396 560116
rect 373356 538212 373408 538218
rect 373356 538154 373408 538160
rect 374092 530460 374144 530466
rect 374092 530402 374144 530408
rect 373264 522912 373316 522918
rect 373264 522854 373316 522860
rect 374000 522912 374052 522918
rect 374000 522854 374052 522860
rect 374012 520146 374040 522854
rect 374104 522034 374132 530402
rect 374472 526998 374500 612031
rect 374564 532642 374592 613935
rect 374656 551954 374684 618423
rect 374826 607336 374882 607345
rect 374826 607271 374882 607280
rect 374734 569936 374790 569945
rect 374734 569871 374790 569880
rect 374644 551948 374696 551954
rect 374644 551890 374696 551896
rect 374748 540802 374776 569871
rect 374736 540796 374788 540802
rect 374736 540738 374788 540744
rect 374552 532636 374604 532642
rect 374552 532578 374604 532584
rect 374840 531282 374868 607271
rect 375392 602857 375420 635462
rect 375484 606937 375512 639775
rect 375576 608569 375604 642194
rect 375668 621625 375696 650218
rect 377416 643346 377444 651986
rect 387154 646912 387210 646921
rect 387154 646847 387210 646856
rect 383106 645280 383162 645289
rect 383106 645215 383162 645224
rect 377404 643340 377456 643346
rect 377404 643282 377456 643288
rect 380532 643340 380584 643346
rect 380532 643282 380584 643288
rect 380070 642832 380126 642841
rect 380070 642767 380126 642776
rect 379058 640520 379114 640529
rect 379058 640455 379114 640464
rect 376852 639124 376904 639130
rect 376852 639066 376904 639072
rect 376760 634500 376812 634506
rect 376760 634442 376812 634448
rect 375654 621616 375710 621625
rect 375654 621551 375710 621560
rect 376206 619168 376262 619177
rect 376206 619103 376262 619112
rect 375746 617536 375802 617545
rect 375746 617471 375802 617480
rect 375654 611008 375710 611017
rect 375654 610943 375710 610952
rect 375562 608560 375618 608569
rect 375562 608495 375618 608504
rect 375470 606928 375526 606937
rect 375470 606863 375526 606872
rect 375562 603664 375618 603673
rect 375562 603599 375618 603608
rect 375378 602848 375434 602857
rect 375378 602783 375434 602792
rect 375012 538552 375064 538558
rect 375012 538494 375064 538500
rect 374828 531276 374880 531282
rect 374828 531218 374880 531224
rect 374460 526992 374512 526998
rect 374460 526934 374512 526940
rect 374092 522028 374144 522034
rect 374092 521970 374144 521976
rect 375024 520146 375052 538494
rect 375576 522102 375604 603599
rect 375668 532409 375696 610943
rect 375760 554062 375788 617471
rect 375838 613456 375894 613465
rect 375838 613391 375894 613400
rect 375852 554742 375880 613391
rect 375930 602032 375986 602041
rect 375930 601967 375986 601976
rect 375944 556850 375972 601967
rect 376022 597136 376078 597145
rect 376022 597071 376078 597080
rect 375932 556844 375984 556850
rect 375932 556786 375984 556792
rect 375840 554736 375892 554742
rect 375840 554678 375892 554684
rect 376036 554402 376064 597071
rect 376114 595504 376170 595513
rect 376114 595439 376170 595448
rect 376024 554396 376076 554402
rect 376024 554338 376076 554344
rect 376128 554334 376156 595439
rect 376116 554328 376168 554334
rect 376116 554270 376168 554276
rect 375748 554056 375800 554062
rect 375748 553998 375800 554004
rect 376024 537192 376076 537198
rect 376024 537134 376076 537140
rect 375654 532400 375710 532409
rect 375654 532335 375710 532344
rect 375564 522096 375616 522102
rect 375564 522038 375616 522044
rect 376036 520146 376064 537134
rect 376220 532098 376248 619103
rect 376298 615904 376354 615913
rect 376298 615839 376354 615848
rect 376312 532710 376340 615839
rect 376772 600409 376800 634442
rect 376864 620809 376892 639066
rect 377220 622464 377272 622470
rect 377218 622432 377220 622441
rect 377272 622432 377274 622441
rect 377218 622367 377274 622376
rect 376850 620800 376906 620809
rect 376850 620735 376906 620744
rect 378598 619984 378654 619993
rect 378598 619919 378654 619928
rect 378322 616720 378378 616729
rect 378322 616655 378378 616664
rect 378046 606112 378102 606121
rect 378046 606047 378102 606056
rect 378060 605834 378088 606047
rect 378060 605806 378272 605834
rect 377034 605296 377090 605305
rect 377034 605231 377090 605240
rect 377048 604586 377076 605231
rect 377036 604580 377088 604586
rect 377036 604522 377088 604528
rect 378048 604512 378100 604518
rect 378046 604480 378048 604489
rect 378100 604480 378102 604489
rect 378046 604415 378102 604424
rect 376758 600400 376814 600409
rect 376758 600335 376814 600344
rect 376850 598768 376906 598777
rect 376850 598703 376906 598712
rect 376758 597952 376814 597961
rect 376758 597887 376814 597896
rect 376772 554470 376800 597887
rect 376864 554538 376892 598703
rect 377954 594688 378010 594697
rect 377954 594623 378010 594632
rect 377968 593434 377996 594623
rect 378046 593872 378102 593881
rect 378046 593807 378102 593816
rect 378060 593502 378088 593807
rect 378048 593496 378100 593502
rect 378048 593438 378100 593444
rect 377956 593428 378008 593434
rect 377956 593370 378008 593376
rect 378046 593056 378102 593065
rect 378046 592991 378102 593000
rect 378060 592346 378088 592991
rect 378048 592340 378100 592346
rect 378048 592282 378100 592288
rect 378046 592240 378102 592249
rect 378046 592175 378102 592184
rect 378060 592142 378088 592175
rect 378048 592136 378100 592142
rect 378048 592078 378100 592084
rect 378046 591424 378102 591433
rect 378046 591359 378102 591368
rect 378060 590714 378088 591359
rect 378048 590708 378100 590714
rect 378048 590650 378100 590656
rect 378046 590608 378102 590617
rect 378046 590543 378102 590552
rect 378060 589966 378088 590543
rect 378048 589960 378100 589966
rect 378048 589902 378100 589908
rect 378046 589792 378102 589801
rect 378046 589727 378102 589736
rect 378060 589354 378088 589727
rect 378048 589348 378100 589354
rect 378048 589290 378100 589296
rect 376942 588976 376998 588985
rect 376942 588911 376998 588920
rect 376956 587926 376984 588911
rect 378046 588160 378102 588169
rect 378046 588095 378102 588104
rect 378060 587994 378088 588095
rect 378048 587988 378100 587994
rect 378048 587930 378100 587936
rect 376944 587920 376996 587926
rect 376944 587862 376996 587868
rect 377770 587344 377826 587353
rect 377770 587279 377826 587288
rect 377784 586974 377812 587279
rect 377772 586968 377824 586974
rect 377772 586910 377824 586916
rect 378048 586628 378100 586634
rect 378048 586570 378100 586576
rect 378060 586537 378088 586570
rect 378046 586528 378102 586537
rect 378046 586463 378102 586472
rect 378046 585712 378102 585721
rect 378046 585647 378102 585656
rect 378060 585206 378088 585647
rect 378048 585200 378100 585206
rect 378048 585142 378100 585148
rect 378046 584896 378102 584905
rect 378046 584831 378102 584840
rect 378060 584186 378088 584831
rect 378048 584180 378100 584186
rect 378048 584122 378100 584128
rect 378046 584080 378102 584089
rect 378046 584015 378102 584024
rect 378060 583778 378088 584015
rect 378048 583772 378100 583778
rect 378048 583714 378100 583720
rect 378046 583264 378102 583273
rect 378046 583199 378102 583208
rect 378060 582554 378088 583199
rect 378048 582548 378100 582554
rect 378048 582490 378100 582496
rect 378046 582448 378102 582457
rect 378046 582383 378048 582392
rect 378100 582383 378102 582392
rect 378048 582354 378100 582360
rect 377862 581632 377918 581641
rect 377862 581567 377918 581576
rect 377876 581058 377904 581567
rect 377864 581052 377916 581058
rect 377864 580994 377916 581000
rect 377126 580816 377182 580825
rect 377126 580751 377182 580760
rect 377140 579698 377168 580751
rect 377586 580000 377642 580009
rect 377586 579935 377642 579944
rect 377600 579766 377628 579935
rect 377588 579760 377640 579766
rect 377588 579702 377640 579708
rect 377128 579692 377180 579698
rect 377128 579634 377180 579640
rect 377034 579184 377090 579193
rect 377034 579119 377090 579128
rect 377048 578270 377076 579119
rect 377862 578368 377918 578377
rect 377862 578303 377864 578312
rect 377916 578303 377918 578312
rect 377864 578274 377916 578280
rect 377036 578264 377088 578270
rect 377036 578206 377088 578212
rect 377126 575920 377182 575929
rect 377126 575855 377182 575864
rect 377140 575550 377168 575855
rect 377128 575544 377180 575550
rect 377128 575486 377180 575492
rect 376942 575104 376998 575113
rect 376942 575039 376998 575048
rect 376956 556034 376984 575039
rect 378046 573472 378102 573481
rect 378046 573407 378102 573416
rect 378060 572762 378088 573407
rect 378048 572756 378100 572762
rect 378048 572698 378100 572704
rect 378046 572656 378102 572665
rect 378046 572591 378102 572600
rect 378060 571946 378088 572591
rect 378048 571940 378100 571946
rect 378048 571882 378100 571888
rect 378046 571840 378102 571849
rect 378046 571775 378102 571784
rect 378060 571402 378088 571775
rect 378048 571396 378100 571402
rect 378048 571338 378100 571344
rect 378046 570344 378102 570353
rect 378102 570302 378180 570330
rect 378046 570279 378102 570288
rect 377034 569392 377090 569401
rect 377034 569327 377090 569336
rect 377048 568614 377076 569327
rect 377036 568608 377088 568614
rect 377036 568550 377088 568556
rect 377770 568576 377826 568585
rect 377770 568511 377826 568520
rect 377784 567866 377812 568511
rect 377772 567860 377824 567866
rect 377772 567802 377824 567808
rect 376944 556028 376996 556034
rect 376944 555970 376996 555976
rect 376852 554532 376904 554538
rect 376852 554474 376904 554480
rect 376760 554464 376812 554470
rect 376760 554406 376812 554412
rect 378152 553246 378180 570302
rect 378140 553240 378192 553246
rect 378140 553182 378192 553188
rect 377036 534404 377088 534410
rect 377036 534346 377088 534352
rect 376300 532704 376352 532710
rect 376300 532646 376352 532652
rect 376208 532092 376260 532098
rect 376208 532034 376260 532040
rect 376666 522744 376722 522753
rect 376666 522679 376722 522688
rect 376680 521830 376708 522679
rect 376668 521824 376720 521830
rect 376668 521766 376720 521772
rect 377048 520146 377076 534346
rect 378244 522986 378272 605806
rect 378336 532030 378364 616655
rect 378414 611824 378470 611833
rect 378414 611759 378470 611768
rect 378428 532137 378456 611759
rect 378506 610192 378562 610201
rect 378506 610127 378562 610136
rect 378520 532273 378548 610127
rect 378612 549982 378640 619919
rect 378874 609376 378930 609385
rect 378874 609311 378930 609320
rect 378690 601216 378746 601225
rect 378690 601151 378746 601160
rect 378704 554606 378732 601151
rect 378782 596320 378838 596329
rect 378782 596255 378838 596264
rect 378796 556986 378824 596255
rect 378784 556980 378836 556986
rect 378784 556922 378836 556928
rect 378692 554600 378744 554606
rect 378692 554542 378744 554548
rect 378600 549976 378652 549982
rect 378600 549918 378652 549924
rect 378506 532264 378562 532273
rect 378506 532199 378562 532208
rect 378414 532128 378470 532137
rect 378414 532063 378470 532072
rect 378324 532024 378376 532030
rect 378324 531966 378376 531972
rect 378888 524414 378916 609311
rect 378876 524408 378928 524414
rect 378876 524350 378928 524356
rect 378232 522980 378284 522986
rect 378232 522922 378284 522928
rect 377954 522880 378010 522889
rect 377954 522815 378010 522824
rect 377968 521762 377996 522815
rect 378048 522300 378100 522306
rect 378048 522242 378100 522248
rect 377956 521756 378008 521762
rect 377956 521698 378008 521704
rect 378060 520146 378088 522242
rect 378782 522200 378838 522209
rect 378782 522135 378838 522144
rect 378796 521694 378824 522135
rect 378784 521688 378836 521694
rect 378784 521630 378836 521636
rect 379072 520146 379100 640455
rect 379796 604580 379848 604586
rect 379796 604522 379848 604528
rect 379612 587920 379664 587926
rect 379612 587862 379664 587868
rect 379520 568608 379572 568614
rect 379520 568550 379572 568556
rect 379532 550458 379560 568550
rect 379520 550452 379572 550458
rect 379520 550394 379572 550400
rect 379624 525570 379652 587862
rect 379704 578264 379756 578270
rect 379704 578206 379756 578212
rect 379612 525564 379664 525570
rect 379612 525506 379664 525512
rect 379716 525502 379744 578206
rect 379808 553382 379836 604522
rect 379888 579692 379940 579698
rect 379888 579634 379940 579640
rect 379796 553376 379848 553382
rect 379796 553318 379848 553324
rect 379900 529650 379928 579634
rect 379980 575544 380032 575550
rect 379980 575486 380032 575492
rect 379992 556102 380020 575486
rect 379980 556096 380032 556102
rect 379980 556038 380032 556044
rect 379888 529644 379940 529650
rect 379888 529586 379940 529592
rect 379704 525496 379756 525502
rect 379704 525438 379756 525444
rect 380084 520146 380112 642767
rect 380544 641034 380572 643282
rect 382096 642388 382148 642394
rect 382096 642330 382148 642336
rect 381082 641880 381138 641889
rect 381082 641815 381138 641824
rect 380532 641028 380584 641034
rect 380532 640970 380584 640976
rect 380164 622464 380216 622470
rect 380164 622406 380216 622412
rect 380176 549234 380204 622406
rect 380900 579760 380952 579766
rect 380900 579702 380952 579708
rect 380164 549228 380216 549234
rect 380164 549170 380216 549176
rect 380912 523138 380940 579702
rect 380990 576736 381046 576745
rect 380990 576671 381046 576680
rect 381004 523705 381032 576671
rect 380990 523696 381046 523705
rect 380990 523631 381046 523640
rect 380912 523110 381032 523138
rect 380898 523016 380954 523025
rect 380898 522951 380954 522960
rect 380912 522306 380940 522951
rect 380900 522300 380952 522306
rect 380900 522242 380952 522248
rect 381004 521422 381032 523110
rect 380992 521416 381044 521422
rect 380992 521358 381044 521364
rect 381096 520146 381124 641815
rect 381268 586968 381320 586974
rect 381268 586910 381320 586916
rect 381176 567860 381228 567866
rect 381176 567802 381228 567808
rect 381188 522238 381216 567802
rect 381280 551886 381308 586910
rect 381452 581052 381504 581058
rect 381452 580994 381504 581000
rect 381360 578332 381412 578338
rect 381360 578274 381412 578280
rect 381268 551880 381320 551886
rect 381268 551822 381320 551828
rect 381372 549098 381400 578274
rect 381464 555966 381492 580994
rect 381452 555960 381504 555966
rect 381452 555902 381504 555908
rect 381360 549092 381412 549098
rect 381360 549034 381412 549040
rect 381176 522232 381228 522238
rect 381176 522174 381228 522180
rect 382108 520146 382136 642330
rect 382832 592340 382884 592346
rect 382832 592282 382884 592288
rect 382464 589348 382516 589354
rect 382464 589290 382516 589296
rect 382280 587988 382332 587994
rect 382280 587930 382332 587936
rect 382292 521626 382320 587930
rect 382372 585200 382424 585206
rect 382372 585142 382424 585148
rect 382280 521620 382332 521626
rect 382280 521562 382332 521568
rect 382384 521558 382412 585142
rect 382476 525706 382504 589290
rect 382740 583772 382792 583778
rect 382740 583714 382792 583720
rect 382648 582548 382700 582554
rect 382648 582490 382700 582496
rect 382556 582412 382608 582418
rect 382556 582354 382608 582360
rect 382464 525700 382516 525706
rect 382464 525642 382516 525648
rect 382568 522714 382596 582354
rect 382660 524142 382688 582490
rect 382752 529854 382780 583714
rect 382844 543250 382872 592282
rect 382832 543244 382884 543250
rect 382832 543186 382884 543192
rect 382740 529848 382792 529854
rect 382740 529790 382792 529796
rect 382648 524136 382700 524142
rect 382648 524078 382700 524084
rect 382556 522708 382608 522714
rect 382556 522650 382608 522656
rect 382372 521552 382424 521558
rect 382372 521494 382424 521500
rect 383120 520146 383148 645215
rect 384120 644564 384172 644570
rect 384120 644506 384172 644512
rect 383752 586628 383804 586634
rect 383752 586570 383804 586576
rect 383660 584180 383712 584186
rect 383660 584122 383712 584128
rect 383672 524278 383700 584122
rect 383764 526862 383792 586570
rect 383844 571940 383896 571946
rect 383844 571882 383896 571888
rect 383856 542298 383884 571882
rect 383936 571396 383988 571402
rect 383936 571338 383988 571344
rect 383948 547806 383976 571338
rect 383936 547800 383988 547806
rect 383936 547742 383988 547748
rect 383844 542292 383896 542298
rect 383844 542234 383896 542240
rect 383752 526856 383804 526862
rect 383752 526798 383804 526804
rect 383660 524272 383712 524278
rect 383660 524214 383712 524220
rect 384132 520146 384160 644506
rect 385132 639328 385184 639334
rect 385132 639270 385184 639276
rect 385040 593496 385092 593502
rect 385040 593438 385092 593444
rect 385052 522850 385080 593438
rect 385040 522844 385092 522850
rect 385040 522786 385092 522792
rect 385144 520146 385172 639270
rect 386144 635248 386196 635254
rect 386144 635190 386196 635196
rect 385316 592136 385368 592142
rect 385316 592078 385368 592084
rect 385224 590708 385276 590714
rect 385224 590650 385276 590656
rect 385236 524346 385264 590650
rect 385328 526930 385356 592078
rect 385408 589960 385460 589966
rect 385408 589902 385460 589908
rect 385420 528562 385448 589902
rect 385408 528556 385460 528562
rect 385408 528498 385460 528504
rect 385316 526924 385368 526930
rect 385316 526866 385368 526872
rect 385224 524340 385276 524346
rect 385224 524282 385276 524288
rect 386156 520146 386184 635190
rect 386420 604512 386472 604518
rect 386420 604454 386472 604460
rect 386432 525774 386460 604454
rect 386510 599584 386566 599593
rect 386510 599519 386566 599528
rect 386524 532001 386552 599519
rect 386604 593428 386656 593434
rect 386604 593370 386656 593376
rect 386616 539306 386644 593370
rect 386696 572756 386748 572762
rect 386696 572698 386748 572704
rect 386604 539300 386656 539306
rect 386604 539242 386656 539248
rect 386510 531992 386566 532001
rect 386510 531927 386566 531936
rect 386420 525768 386472 525774
rect 386420 525710 386472 525716
rect 386708 522782 386736 572698
rect 386696 522776 386748 522782
rect 386696 522718 386748 522724
rect 387168 520146 387196 646847
rect 392214 646368 392270 646377
rect 392214 646303 392270 646312
rect 391202 646232 391258 646241
rect 391202 646167 391258 646176
rect 388166 646096 388222 646105
rect 388166 646031 388222 646040
rect 387800 641028 387852 641034
rect 387800 640970 387852 640976
rect 387812 636206 387840 640970
rect 387800 636200 387852 636206
rect 387800 636142 387852 636148
rect 387708 634432 387760 634438
rect 387708 634374 387760 634380
rect 387720 627230 387748 634374
rect 387708 627224 387760 627230
rect 387708 627166 387760 627172
rect 388180 520146 388208 646031
rect 390192 644632 390244 644638
rect 390192 644574 390244 644580
rect 389180 643544 389232 643550
rect 389180 643486 389232 643492
rect 389192 520146 389220 643486
rect 390204 520146 390232 644574
rect 391216 520146 391244 646167
rect 391388 636200 391440 636206
rect 391388 636142 391440 636148
rect 391296 635316 391348 635322
rect 391296 635258 391348 635264
rect 391308 522714 391336 635258
rect 391400 621722 391428 636142
rect 391388 621716 391440 621722
rect 391388 621658 391440 621664
rect 391296 522708 391348 522714
rect 391296 522650 391348 522656
rect 392228 520146 392256 646303
rect 393228 644836 393280 644842
rect 393228 644778 393280 644784
rect 392582 634536 392638 634545
rect 392582 634471 392638 634480
rect 392596 613329 392624 634471
rect 392582 613320 392638 613329
rect 392582 613255 392638 613264
rect 393240 520146 393268 644778
rect 395250 644736 395306 644745
rect 395250 644671 395306 644680
rect 394238 644600 394294 644609
rect 394238 644535 394294 644544
rect 393962 635216 394018 635225
rect 393962 635151 394018 635160
rect 393976 522481 394004 635151
rect 393962 522472 394018 522481
rect 393962 522407 394018 522416
rect 394252 520146 394280 644535
rect 395264 520146 395292 644671
rect 397276 637968 397328 637974
rect 397276 637910 397328 637916
rect 395344 637628 395396 637634
rect 395344 637570 395396 637576
rect 395356 522986 395384 637570
rect 395344 522980 395396 522986
rect 395344 522922 395396 522928
rect 396172 522980 396224 522986
rect 396172 522922 396224 522928
rect 396184 520146 396212 522922
rect 397288 520146 397316 637910
rect 397472 599729 397500 703520
rect 407394 645144 407450 645153
rect 407394 645079 407450 645088
rect 401322 645008 401378 645017
rect 401322 644943 401378 644952
rect 398286 644872 398342 644881
rect 398286 644807 398342 644816
rect 398104 621716 398156 621722
rect 398104 621658 398156 621664
rect 397550 613320 397606 613329
rect 397550 613255 397606 613264
rect 397564 607209 397592 613255
rect 398116 612066 398144 621658
rect 398104 612060 398156 612066
rect 398104 612002 398156 612008
rect 397550 607200 397606 607209
rect 397550 607135 397606 607144
rect 397458 599720 397514 599729
rect 397458 599655 397514 599664
rect 398300 520146 398328 644807
rect 400864 638036 400916 638042
rect 400864 637978 400916 637984
rect 399300 637764 399352 637770
rect 399300 637706 399352 637712
rect 399312 520146 399340 637706
rect 400312 637696 400364 637702
rect 400312 637638 400364 637644
rect 400324 520146 400352 637638
rect 400772 627224 400824 627230
rect 400772 627166 400824 627172
rect 400784 621722 400812 627166
rect 400772 621716 400824 621722
rect 400772 621658 400824 621664
rect 400876 522986 400904 637978
rect 400954 607200 401010 607209
rect 400954 607135 401010 607144
rect 400968 596873 400996 607135
rect 400954 596864 401010 596873
rect 400954 596799 401010 596808
rect 400864 522980 400916 522986
rect 400864 522922 400916 522928
rect 401336 520146 401364 644943
rect 403348 639260 403400 639266
rect 403348 639202 403400 639208
rect 402336 522980 402388 522986
rect 402336 522922 402388 522928
rect 402348 520146 402376 522922
rect 403360 520146 403388 639202
rect 405372 639192 405424 639198
rect 405372 639134 405424 639140
rect 403624 639056 403676 639062
rect 403624 638998 403676 639004
rect 403636 522986 403664 638998
rect 403624 522980 403676 522986
rect 403624 522922 403676 522928
rect 404268 522980 404320 522986
rect 404268 522922 404320 522928
rect 404280 521778 404308 522922
rect 404280 521750 404400 521778
rect 404372 520146 404400 521750
rect 405384 520146 405412 639134
rect 406384 638988 406436 638994
rect 406384 638930 406436 638936
rect 406396 520146 406424 638930
rect 406476 621716 406528 621722
rect 406476 621658 406528 621664
rect 406488 610638 406516 621658
rect 406476 610632 406528 610638
rect 406476 610574 406528 610580
rect 407408 520146 407436 645079
rect 412456 635180 412508 635186
rect 412456 635122 412508 635128
rect 410524 635112 410576 635118
rect 410524 635054 410576 635060
rect 409420 635044 409472 635050
rect 409420 634986 409472 634992
rect 407764 634976 407816 634982
rect 407764 634918 407816 634924
rect 407776 522986 407804 634918
rect 407764 522980 407816 522986
rect 407764 522922 407816 522928
rect 408408 522708 408460 522714
rect 408408 522650 408460 522656
rect 408420 520146 408448 522650
rect 409432 520146 409460 634986
rect 410536 522986 410564 635054
rect 411444 634840 411496 634846
rect 411444 634782 411496 634788
rect 410616 612060 410668 612066
rect 410616 612002 410668 612008
rect 410628 604518 410656 612002
rect 410616 604512 410668 604518
rect 410616 604454 410668 604460
rect 410432 522980 410484 522986
rect 410432 522922 410484 522928
rect 410524 522980 410576 522986
rect 410524 522922 410576 522928
rect 410444 520146 410472 522922
rect 411456 520146 411484 634782
rect 412468 520146 412496 635122
rect 413284 604512 413336 604518
rect 413284 604454 413336 604460
rect 413296 587858 413324 604454
rect 413664 599622 413692 703520
rect 429856 657801 429884 703520
rect 429842 657792 429898 657801
rect 429842 657727 429898 657736
rect 461582 652216 461638 652225
rect 461582 652151 461638 652160
rect 425610 646776 425666 646785
rect 425610 646711 425666 646720
rect 424598 646640 424654 646649
rect 424598 646575 424654 646584
rect 423586 646504 423642 646513
rect 423586 646439 423642 646448
rect 419540 643408 419592 643414
rect 419540 643350 419592 643356
rect 418526 639160 418582 639169
rect 418526 639095 418582 639104
rect 417514 639024 417570 639033
rect 417514 638959 417570 638968
rect 414664 638240 414716 638246
rect 414664 638182 414716 638188
rect 414480 634908 414532 634914
rect 414480 634850 414532 634856
rect 413652 599616 413704 599622
rect 413652 599558 413704 599564
rect 413284 587852 413336 587858
rect 413284 587794 413336 587800
rect 413376 522980 413428 522986
rect 413376 522922 413428 522928
rect 413388 520146 413416 522922
rect 414492 520146 414520 634850
rect 414676 522986 414704 638182
rect 416502 635080 416558 635089
rect 416502 635015 416558 635024
rect 416042 596864 416098 596873
rect 416042 596799 416098 596808
rect 416056 536761 416084 596799
rect 416136 587852 416188 587858
rect 416136 587794 416188 587800
rect 416148 575550 416176 587794
rect 416136 575544 416188 575550
rect 416136 575486 416188 575492
rect 416042 536752 416098 536761
rect 416042 536687 416098 536696
rect 414664 522980 414716 522986
rect 414664 522922 414716 522928
rect 415492 522980 415544 522986
rect 415492 522922 415544 522928
rect 415504 520146 415532 522922
rect 416516 520146 416544 635015
rect 417528 520146 417556 638959
rect 418540 520146 418568 639095
rect 418804 550180 418856 550186
rect 418804 550122 418856 550128
rect 418816 522714 418844 550122
rect 418804 522708 418856 522714
rect 418804 522650 418856 522656
rect 419552 520146 419580 643350
rect 421564 639396 421616 639402
rect 421564 639338 421616 639344
rect 420184 610632 420236 610638
rect 420184 610574 420236 610580
rect 420196 589966 420224 610574
rect 420184 589960 420236 589966
rect 420184 589902 420236 589908
rect 419632 575544 419684 575550
rect 419632 575486 419684 575492
rect 419644 570654 419672 575486
rect 419632 570648 419684 570654
rect 419632 570590 419684 570596
rect 420458 522472 420514 522481
rect 420514 522430 420592 522458
rect 420458 522407 420514 522416
rect 420564 520146 420592 522430
rect 421576 520146 421604 639338
rect 422574 638616 422630 638625
rect 422574 638551 422630 638560
rect 422588 520146 422616 638551
rect 423600 520146 423628 646439
rect 424612 520146 424640 646575
rect 425624 520146 425652 646711
rect 458824 642048 458876 642054
rect 458824 641990 458876 641996
rect 456156 636744 456208 636750
rect 456156 636686 456208 636692
rect 456064 636608 456116 636614
rect 456064 636550 456116 636556
rect 453304 636404 453356 636410
rect 453304 636346 453356 636352
rect 428464 589960 428516 589966
rect 428464 589902 428516 589908
rect 428476 571334 428504 589902
rect 428464 571328 428516 571334
rect 428464 571270 428516 571276
rect 433984 571328 434036 571334
rect 433984 571270 434036 571276
rect 429200 570648 429252 570654
rect 429200 570590 429252 570596
rect 429212 567254 429240 570590
rect 429200 567248 429252 567254
rect 429200 567190 429252 567196
rect 432052 567248 432104 567254
rect 432052 567190 432104 567196
rect 432064 562358 432092 567190
rect 432052 562352 432104 562358
rect 432052 562294 432104 562300
rect 427634 559600 427690 559609
rect 427634 559535 427690 559544
rect 426622 548856 426678 548865
rect 426622 548791 426678 548800
rect 426636 520146 426664 548791
rect 427648 520146 427676 559535
rect 432694 555656 432750 555665
rect 432694 555591 432750 555600
rect 428646 540560 428702 540569
rect 428646 540495 428702 540504
rect 428660 520146 428688 540495
rect 429658 533488 429714 533497
rect 429658 533423 429714 533432
rect 429672 520146 429700 533423
rect 430580 528148 430632 528154
rect 430580 528090 430632 528096
rect 430592 520146 430620 528090
rect 431682 522336 431738 522345
rect 431682 522271 431738 522280
rect 431696 520146 431724 522271
rect 432708 520146 432736 555591
rect 433706 555384 433762 555393
rect 433706 555319 433762 555328
rect 433720 520146 433748 555319
rect 433996 552022 434024 571270
rect 444288 562352 444340 562358
rect 444288 562294 444340 562300
rect 444300 559638 444328 562294
rect 444288 559632 444340 559638
rect 444288 559574 444340 559580
rect 445850 557016 445906 557025
rect 445850 556951 445906 556960
rect 434720 555212 434772 555218
rect 434720 555154 434772 555160
rect 433984 552016 434036 552022
rect 433984 551958 434036 551964
rect 434732 520146 434760 555154
rect 436100 552016 436152 552022
rect 436100 551958 436152 551964
rect 436112 548418 436140 551958
rect 443826 551440 443882 551449
rect 443826 551375 443882 551384
rect 436100 548412 436152 548418
rect 436100 548354 436152 548360
rect 441620 548412 441672 548418
rect 441620 548354 441672 548360
rect 441632 545222 441660 548354
rect 441620 545216 441672 545222
rect 441620 545158 441672 545164
rect 439778 541784 439834 541793
rect 439778 541719 439834 541728
rect 436374 536752 436430 536761
rect 436374 536687 436430 536696
rect 436388 532545 436416 536687
rect 436374 532536 436430 532545
rect 436374 532471 436430 532480
rect 436742 531312 436798 531321
rect 436742 531247 436798 531256
rect 436008 529236 436060 529242
rect 436008 529178 436060 529184
rect 436020 522782 436048 529178
rect 436008 522776 436060 522782
rect 436008 522718 436060 522724
rect 435732 522436 435784 522442
rect 435732 522378 435784 522384
rect 435744 520146 435772 522378
rect 436756 520146 436784 531247
rect 437754 531176 437810 531185
rect 437754 531111 437810 531120
rect 437768 520146 437796 531111
rect 438766 531040 438822 531049
rect 438766 530975 438822 530984
rect 438780 520146 438808 530975
rect 439792 520146 439820 541719
rect 440882 532536 440938 532545
rect 440882 532471 440938 532480
rect 440790 530904 440846 530913
rect 440790 530839 440846 530848
rect 440804 520146 440832 530839
rect 440896 528465 440924 532471
rect 440882 528456 440938 528465
rect 440882 528391 440938 528400
rect 442724 527944 442776 527950
rect 442724 527886 442776 527892
rect 441710 526552 441766 526561
rect 441766 526510 441844 526538
rect 441710 526487 441766 526496
rect 441816 520146 441844 526510
rect 442736 520146 442764 527886
rect 443840 520146 443868 551375
rect 444380 545216 444432 545222
rect 444380 545158 444432 545164
rect 444392 540938 444420 545158
rect 444380 540932 444432 540938
rect 444380 540874 444432 540880
rect 444838 536072 444894 536081
rect 444838 536007 444894 536016
rect 444286 528456 444342 528465
rect 444286 528391 444342 528400
rect 444300 526561 444328 528391
rect 444286 526552 444342 526561
rect 444286 526487 444342 526496
rect 444852 520146 444880 536007
rect 445864 520146 445892 556951
rect 446862 556880 446918 556889
rect 446862 556815 446918 556824
rect 446876 520146 446904 556815
rect 447874 556744 447930 556753
rect 447874 556679 447930 556688
rect 447232 540932 447284 540938
rect 447232 540874 447284 540880
rect 447244 536382 447272 540874
rect 447232 536376 447284 536382
rect 447232 536318 447284 536324
rect 447888 520146 447916 556679
rect 448888 556640 448940 556646
rect 448888 556582 448940 556588
rect 448900 520146 448928 556582
rect 449900 556572 449952 556578
rect 449900 556514 449952 556520
rect 449912 520146 449940 556514
rect 450912 556504 450964 556510
rect 450912 556446 450964 556452
rect 450924 520146 450952 556446
rect 452936 556436 452988 556442
rect 452936 556378 452988 556384
rect 451924 522164 451976 522170
rect 451924 522106 451976 522112
rect 451936 520146 451964 522106
rect 452948 520146 452976 556378
rect 453316 525094 453344 636346
rect 453948 556368 454000 556374
rect 453948 556310 454000 556316
rect 453304 525088 453356 525094
rect 453304 525030 453356 525036
rect 453960 520146 453988 556310
rect 454960 556300 455012 556306
rect 454960 556242 455012 556248
rect 454972 520146 455000 556242
rect 455970 544640 456026 544649
rect 455970 544575 456026 544584
rect 455984 520146 456012 544575
rect 456076 523734 456104 636550
rect 456168 536314 456196 636686
rect 456800 536376 456852 536382
rect 456800 536318 456852 536324
rect 456156 536308 456208 536314
rect 456156 536250 456208 536256
rect 456812 529582 456840 536318
rect 457996 536240 458048 536246
rect 457996 536182 458048 536188
rect 456800 529576 456852 529582
rect 456800 529518 456852 529524
rect 456064 523728 456116 523734
rect 456064 523670 456116 523676
rect 456984 522368 457036 522374
rect 456984 522310 457036 522316
rect 456996 520146 457024 522310
rect 458008 520146 458036 536182
rect 458836 529514 458864 641990
rect 458916 640552 458968 640558
rect 458916 640494 458968 640500
rect 458824 529508 458876 529514
rect 458824 529450 458876 529456
rect 458928 529242 458956 640494
rect 459008 636676 459060 636682
rect 459008 636618 459060 636624
rect 459020 536246 459048 636618
rect 459100 559632 459152 559638
rect 459100 559574 459152 559580
rect 459112 548826 459140 559574
rect 460020 555144 460072 555150
rect 460020 555086 460072 555092
rect 459100 548820 459152 548826
rect 459100 548762 459152 548768
rect 459008 536240 459060 536246
rect 459008 536182 459060 536188
rect 459006 530632 459062 530641
rect 459006 530567 459062 530576
rect 458916 529236 458968 529242
rect 458916 529178 458968 529184
rect 459020 520146 459048 530567
rect 460032 520146 460060 555086
rect 461030 554160 461086 554169
rect 461030 554095 461086 554104
rect 461044 520146 461072 554095
rect 461596 523705 461624 652151
rect 461766 650856 461822 650865
rect 461766 650791 461822 650800
rect 461674 648136 461730 648145
rect 461674 648071 461730 648080
rect 461582 523696 461638 523705
rect 461582 523631 461638 523640
rect 461688 521529 461716 648071
rect 461780 530777 461808 650791
rect 462332 600030 462360 703520
rect 478524 699718 478552 703520
rect 478512 699712 478564 699718
rect 478512 699654 478564 699660
rect 479524 699712 479576 699718
rect 479524 699654 479576 699660
rect 475382 654936 475438 654945
rect 475382 654871 475438 654880
rect 463146 653576 463202 653585
rect 463146 653511 463202 653520
rect 462964 646128 463016 646134
rect 462964 646070 463016 646076
rect 462320 600024 462372 600030
rect 462320 599966 462372 599972
rect 462044 548140 462096 548146
rect 462044 548082 462096 548088
rect 461766 530768 461822 530777
rect 461766 530703 461822 530712
rect 461674 521520 461730 521529
rect 461674 521455 461730 521464
rect 462056 520146 462084 548082
rect 462976 526522 463004 646070
rect 463056 552832 463108 552838
rect 463056 552774 463108 552780
rect 462964 526516 463016 526522
rect 462964 526458 463016 526464
rect 463068 520146 463096 552774
rect 463160 533497 463188 653511
rect 465722 653440 465778 653449
rect 465722 653375 465778 653384
rect 464344 651500 464396 651506
rect 464344 651442 464396 651448
rect 463240 637900 463292 637906
rect 463240 637842 463292 637848
rect 463146 533488 463202 533497
rect 463146 533423 463202 533432
rect 463252 527950 463280 637842
rect 464066 534712 464122 534721
rect 464066 534647 464122 534656
rect 463240 527944 463292 527950
rect 463240 527886 463292 527892
rect 464080 520146 464108 534647
rect 464356 530806 464384 651442
rect 464436 644768 464488 644774
rect 464436 644710 464488 644716
rect 464344 530800 464396 530806
rect 464344 530742 464396 530748
rect 464448 530602 464476 644710
rect 464528 643272 464580 643278
rect 464528 643214 464580 643220
rect 464540 530874 464568 643214
rect 464620 642184 464672 642190
rect 464620 642126 464672 642132
rect 464528 530868 464580 530874
rect 464528 530810 464580 530816
rect 464632 530670 464660 642126
rect 465080 544604 465132 544610
rect 465080 544546 465132 544552
rect 464620 530664 464672 530670
rect 464620 530606 464672 530612
rect 464436 530596 464488 530602
rect 464436 530538 464488 530544
rect 465092 520146 465120 544546
rect 465736 533633 465764 653375
rect 471334 653304 471390 653313
rect 471334 653239 471390 653248
rect 469862 651944 469918 651953
rect 469862 651879 469918 651888
rect 468482 651808 468538 651817
rect 468482 651743 468538 651752
rect 467378 650720 467434 650729
rect 467378 650655 467434 650664
rect 467194 650448 467250 650457
rect 467194 650383 467250 650392
rect 467104 648848 467156 648854
rect 467104 648790 467156 648796
rect 465816 640756 465868 640762
rect 465816 640698 465868 640704
rect 465722 533624 465778 533633
rect 465722 533559 465778 533568
rect 465828 530738 465856 640698
rect 465906 636984 465962 636993
rect 465906 636919 465962 636928
rect 465920 536081 465948 636919
rect 466920 548820 466972 548826
rect 466920 548762 466972 548768
rect 466932 542978 466960 548762
rect 467012 547324 467064 547330
rect 467012 547266 467064 547272
rect 466920 542972 466972 542978
rect 466920 542914 466972 542920
rect 466092 539844 466144 539850
rect 466092 539786 466144 539792
rect 465906 536072 465962 536081
rect 465906 536007 465962 536016
rect 465816 530732 465868 530738
rect 465816 530674 465868 530680
rect 466104 520146 466132 539786
rect 467024 520146 467052 547266
rect 467116 525162 467144 648790
rect 467208 527921 467236 650383
rect 467286 649496 467342 649505
rect 467286 649431 467342 649440
rect 467300 530641 467328 649431
rect 467286 530632 467342 530641
rect 467286 530567 467342 530576
rect 467194 527912 467250 527921
rect 467194 527847 467250 527856
rect 467392 527785 467420 650655
rect 468116 541816 468168 541822
rect 468116 541758 468168 541764
rect 467378 527776 467434 527785
rect 467378 527711 467434 527720
rect 467104 525156 467156 525162
rect 467104 525098 467156 525104
rect 468128 520146 468156 541758
rect 468496 528193 468524 651743
rect 468574 636576 468630 636585
rect 468574 636511 468630 636520
rect 468482 528184 468538 528193
rect 468482 528119 468538 528128
rect 468588 521665 468616 636511
rect 469128 530392 469180 530398
rect 469128 530334 469180 530340
rect 468574 521656 468630 521665
rect 468574 521591 468630 521600
rect 469140 520146 469168 530334
rect 469876 523569 469904 651879
rect 469956 648712 470008 648718
rect 469956 648654 470008 648660
rect 469968 525230 469996 648654
rect 471244 647420 471296 647426
rect 471244 647362 471296 647368
rect 470046 636440 470102 636449
rect 470046 636375 470102 636384
rect 469956 525224 470008 525230
rect 469956 525166 470008 525172
rect 470060 523938 470088 636375
rect 470140 542972 470192 542978
rect 470140 542914 470192 542920
rect 470152 534954 470180 542914
rect 470140 534948 470192 534954
rect 470140 534890 470192 534896
rect 470140 530256 470192 530262
rect 470140 530198 470192 530204
rect 470048 523932 470100 523938
rect 470048 523874 470100 523880
rect 469862 523560 469918 523569
rect 469862 523495 469918 523504
rect 470152 520146 470180 530198
rect 471060 522096 471112 522102
rect 471060 522038 471112 522044
rect 471072 520146 471100 522038
rect 471256 521150 471284 647362
rect 471348 533905 471376 653239
rect 472624 648644 472676 648650
rect 472624 648586 472676 648592
rect 471520 639464 471572 639470
rect 471520 639406 471572 639412
rect 471428 635452 471480 635458
rect 471428 635394 471480 635400
rect 471334 533896 471390 533905
rect 471334 533831 471390 533840
rect 471244 521144 471296 521150
rect 471244 521086 471296 521092
rect 471440 521082 471468 635394
rect 471532 530942 471560 639406
rect 471520 530936 471572 530942
rect 471520 530878 471572 530884
rect 472164 530188 472216 530194
rect 472164 530130 472216 530136
rect 471428 521076 471480 521082
rect 471428 521018 471480 521024
rect 472176 520146 472204 530130
rect 472636 522374 472664 648586
rect 472900 647488 472952 647494
rect 472900 647430 472952 647436
rect 472716 643136 472768 643142
rect 472716 643078 472768 643084
rect 472728 525298 472756 643078
rect 472808 640688 472860 640694
rect 472808 640630 472860 640636
rect 472716 525292 472768 525298
rect 472716 525234 472768 525240
rect 472820 522442 472848 640630
rect 472912 531010 472940 647430
rect 472992 636336 473044 636342
rect 472992 636278 473044 636284
rect 473004 536382 473032 636278
rect 473176 555076 473228 555082
rect 473176 555018 473228 555024
rect 472992 536376 473044 536382
rect 472992 536318 473044 536324
rect 472900 531004 472952 531010
rect 472900 530946 472952 530952
rect 472808 522436 472860 522442
rect 472808 522378 472860 522384
rect 472624 522368 472676 522374
rect 472624 522310 472676 522316
rect 473188 520146 473216 555018
rect 475200 555008 475252 555014
rect 475200 554950 475252 554956
rect 474096 522572 474148 522578
rect 474096 522514 474148 522520
rect 474108 520146 474136 522514
rect 475212 520146 475240 554950
rect 475396 533089 475424 654871
rect 478234 651400 478290 651409
rect 478234 651335 478290 651344
rect 478144 647352 478196 647358
rect 478144 647294 478196 647300
rect 476764 644700 476816 644706
rect 476764 644642 476816 644648
rect 475566 642288 475622 642297
rect 475566 642223 475622 642232
rect 475476 641912 475528 641918
rect 475476 641854 475528 641860
rect 475382 533080 475438 533089
rect 475382 533015 475438 533024
rect 475488 522578 475516 641854
rect 475476 522572 475528 522578
rect 475476 522514 475528 522520
rect 475580 522481 475608 642223
rect 475750 642152 475806 642161
rect 475750 642087 475806 642096
rect 475660 638172 475712 638178
rect 475660 638114 475712 638120
rect 475672 522850 475700 638114
rect 475660 522844 475712 522850
rect 475660 522786 475712 522792
rect 475566 522472 475622 522481
rect 475566 522407 475622 522416
rect 475764 522345 475792 642087
rect 475844 534948 475896 534954
rect 475844 534890 475896 534896
rect 475856 528426 475884 534890
rect 476776 531078 476804 644642
rect 477224 554192 477276 554198
rect 477224 554134 477276 554140
rect 476764 531072 476816 531078
rect 476764 531014 476816 531020
rect 475844 528420 475896 528426
rect 475844 528362 475896 528368
rect 476120 522640 476172 522646
rect 476120 522582 476172 522588
rect 475750 522336 475806 522345
rect 475750 522271 475806 522280
rect 476132 520146 476160 522582
rect 477236 520146 477264 554134
rect 478156 525434 478184 647294
rect 478248 534041 478276 651335
rect 479248 538892 479300 538898
rect 479248 538834 479300 538840
rect 478328 537600 478380 537606
rect 478328 537542 478380 537548
rect 478234 534032 478290 534041
rect 478234 533967 478290 533976
rect 478144 525428 478196 525434
rect 478144 525370 478196 525376
rect 478340 520146 478368 537542
rect 314304 520118 314348 520146
rect 315316 520118 315360 520146
rect 316328 520118 316372 520146
rect 317340 520118 317384 520146
rect 318352 520118 318396 520146
rect 319364 520118 319408 520146
rect 320376 520118 320420 520146
rect 321388 520118 321432 520146
rect 322400 520118 322444 520146
rect 323412 520118 323456 520146
rect 324424 520118 324468 520146
rect 325436 520118 325480 520146
rect 326448 520118 326492 520146
rect 327460 520118 327504 520146
rect 328472 520118 328516 520146
rect 329484 520118 329528 520146
rect 330496 520118 330540 520146
rect 331508 520118 331552 520146
rect 332520 520118 332564 520146
rect 333532 520118 333576 520146
rect 334544 520118 334588 520146
rect 335556 520118 335600 520146
rect 336568 520118 336612 520146
rect 337488 520118 337624 520146
rect 338592 520118 338636 520146
rect 339604 520118 339648 520146
rect 340616 520118 340660 520146
rect 341628 520118 341672 520146
rect 342640 520118 342684 520146
rect 343652 520118 343696 520146
rect 344664 520118 344708 520146
rect 345676 520118 345720 520146
rect 346688 520118 346732 520146
rect 347700 520118 347744 520146
rect 348712 520118 348756 520146
rect 349724 520118 349768 520146
rect 350736 520118 350780 520146
rect 351748 520118 351792 520146
rect 352760 520118 352804 520146
rect 353772 520118 353816 520146
rect 354784 520118 354828 520146
rect 355796 520118 355840 520146
rect 356808 520118 356852 520146
rect 357820 520118 357864 520146
rect 358832 520118 358876 520146
rect 359844 520118 359888 520146
rect 360856 520118 360900 520146
rect 361868 520118 361912 520146
rect 362880 520118 362924 520146
rect 363892 520118 363936 520146
rect 364904 520118 364948 520146
rect 365916 520118 365960 520146
rect 366928 520118 366972 520146
rect 367940 520118 367984 520146
rect 368952 520118 368996 520146
rect 369964 520118 370008 520146
rect 370976 520118 371020 520146
rect 371988 520118 372032 520146
rect 373000 520118 373044 520146
rect 374012 520118 374056 520146
rect 375024 520118 375068 520146
rect 376036 520118 376080 520146
rect 377048 520118 377092 520146
rect 378060 520118 378104 520146
rect 379072 520118 379116 520146
rect 380084 520118 380128 520146
rect 381096 520118 381140 520146
rect 382108 520118 382152 520146
rect 383120 520118 383164 520146
rect 384132 520118 384176 520146
rect 385144 520118 385188 520146
rect 386156 520118 386200 520146
rect 387168 520118 387212 520146
rect 388180 520118 388224 520146
rect 389192 520118 389236 520146
rect 390204 520118 390248 520146
rect 391216 520118 391260 520146
rect 392228 520118 392272 520146
rect 393240 520118 393284 520146
rect 394252 520118 394296 520146
rect 395264 520118 395308 520146
rect 396184 520118 396320 520146
rect 397288 520118 397332 520146
rect 398300 520118 398344 520146
rect 399312 520118 399356 520146
rect 400324 520118 400368 520146
rect 401336 520118 401380 520146
rect 402348 520118 402392 520146
rect 403360 520118 403404 520146
rect 404372 520118 404416 520146
rect 405384 520118 405428 520146
rect 406396 520118 406440 520146
rect 407408 520118 407452 520146
rect 408420 520118 408464 520146
rect 409432 520118 409476 520146
rect 410444 520118 410488 520146
rect 411456 520118 411500 520146
rect 412468 520118 412512 520146
rect 413388 520118 413524 520146
rect 414492 520118 414536 520146
rect 415504 520118 415548 520146
rect 416516 520118 416560 520146
rect 417528 520118 417572 520146
rect 418540 520118 418584 520146
rect 419552 520118 419596 520146
rect 420564 520118 420608 520146
rect 421576 520118 421620 520146
rect 422588 520118 422632 520146
rect 423600 520118 423644 520146
rect 424612 520118 424656 520146
rect 425624 520118 425668 520146
rect 426636 520118 426680 520146
rect 427648 520118 427692 520146
rect 428660 520118 428704 520146
rect 429672 520118 429716 520146
rect 430592 520118 430728 520146
rect 431696 520118 431740 520146
rect 432708 520118 432752 520146
rect 433720 520118 433764 520146
rect 434732 520118 434776 520146
rect 435744 520118 435788 520146
rect 436756 520118 436800 520146
rect 437768 520118 437812 520146
rect 438780 520118 438824 520146
rect 439792 520118 439836 520146
rect 440804 520118 440848 520146
rect 441816 520118 441860 520146
rect 442736 520118 442872 520146
rect 443840 520118 443884 520146
rect 444852 520118 444896 520146
rect 445864 520118 445908 520146
rect 446876 520118 446920 520146
rect 447888 520118 447932 520146
rect 448900 520118 448944 520146
rect 449912 520118 449956 520146
rect 450924 520118 450968 520146
rect 451936 520118 451980 520146
rect 452948 520118 452992 520146
rect 453960 520118 454004 520146
rect 454972 520118 455016 520146
rect 455984 520118 456028 520146
rect 456996 520118 457040 520146
rect 458008 520118 458052 520146
rect 459020 520118 459064 520146
rect 460032 520118 460076 520146
rect 461044 520118 461088 520146
rect 462056 520118 462100 520146
rect 463068 520118 463112 520146
rect 464080 520118 464124 520146
rect 465092 520118 465136 520146
rect 466104 520118 466148 520146
rect 467024 520118 467160 520146
rect 468128 520118 468172 520146
rect 469140 520118 469184 520146
rect 470152 520118 470196 520146
rect 471072 520118 471208 520146
rect 472176 520118 472220 520146
rect 473188 520118 473232 520146
rect 474108 520118 474244 520146
rect 475212 520118 475256 520146
rect 476132 520118 476268 520146
rect 477236 520118 477280 520146
rect 313308 519860 313336 520118
rect 314320 519860 314348 520118
rect 315332 519860 315360 520118
rect 316344 519860 316372 520118
rect 317356 519860 317384 520118
rect 318368 519860 318396 520118
rect 319380 519860 319408 520118
rect 320392 519860 320420 520118
rect 321404 519860 321432 520118
rect 322416 519860 322444 520118
rect 323428 519860 323456 520118
rect 324440 519860 324468 520118
rect 325452 519860 325480 520118
rect 326464 519860 326492 520118
rect 327476 519860 327504 520118
rect 328488 519860 328516 520118
rect 329500 519860 329528 520118
rect 330512 519860 330540 520118
rect 331524 519860 331552 520118
rect 332536 519860 332564 520118
rect 333548 519860 333576 520118
rect 334560 519860 334588 520118
rect 335572 519860 335600 520118
rect 336584 519860 336612 520118
rect 337596 519860 337624 520118
rect 338608 519860 338636 520118
rect 339620 519860 339648 520118
rect 340632 519860 340660 520118
rect 341644 519860 341672 520118
rect 342656 519860 342684 520118
rect 343668 519860 343696 520118
rect 344680 519860 344708 520118
rect 345692 519860 345720 520118
rect 346704 519860 346732 520118
rect 347716 519860 347744 520118
rect 348728 519860 348756 520118
rect 349740 519860 349768 520118
rect 350752 519860 350780 520118
rect 351764 519860 351792 520118
rect 352776 519860 352804 520118
rect 353788 519860 353816 520118
rect 354800 519860 354828 520118
rect 355812 519860 355840 520118
rect 356824 519860 356852 520118
rect 357836 519860 357864 520118
rect 358848 519860 358876 520118
rect 359860 519860 359888 520118
rect 360872 519860 360900 520118
rect 361884 519860 361912 520118
rect 362896 519860 362924 520118
rect 363908 519860 363936 520118
rect 364920 519860 364948 520118
rect 365932 519860 365960 520118
rect 366944 519860 366972 520118
rect 367956 519860 367984 520118
rect 368968 519860 368996 520118
rect 369980 519860 370008 520118
rect 370992 519860 371020 520118
rect 372004 519860 372032 520118
rect 373016 519860 373044 520118
rect 374028 519860 374056 520118
rect 375040 519860 375068 520118
rect 376052 519860 376080 520118
rect 377064 519860 377092 520118
rect 378076 519860 378104 520118
rect 379088 519860 379116 520118
rect 380100 519860 380128 520118
rect 381112 519860 381140 520118
rect 382124 519860 382152 520118
rect 383136 519860 383164 520118
rect 384148 519860 384176 520118
rect 385160 519860 385188 520118
rect 386172 519860 386200 520118
rect 387184 519860 387212 520118
rect 388196 519860 388224 520118
rect 389208 519860 389236 520118
rect 390220 519860 390248 520118
rect 391232 519860 391260 520118
rect 392244 519860 392272 520118
rect 393256 519860 393284 520118
rect 394268 519860 394296 520118
rect 395280 519860 395308 520118
rect 396292 519860 396320 520118
rect 397304 519860 397332 520118
rect 398316 519860 398344 520118
rect 399328 519860 399356 520118
rect 400340 519860 400368 520118
rect 401352 519860 401380 520118
rect 402364 519860 402392 520118
rect 403376 519860 403404 520118
rect 404388 519860 404416 520118
rect 405400 519860 405428 520118
rect 406412 519860 406440 520118
rect 407424 519860 407452 520118
rect 408436 519860 408464 520118
rect 409448 519860 409476 520118
rect 410460 519860 410488 520118
rect 411472 519860 411500 520118
rect 412484 519860 412512 520118
rect 413496 519860 413524 520118
rect 414508 519860 414536 520118
rect 415520 519860 415548 520118
rect 416532 519860 416560 520118
rect 417544 519860 417572 520118
rect 418556 519860 418584 520118
rect 419568 519860 419596 520118
rect 420580 519860 420608 520118
rect 421592 519860 421620 520118
rect 422604 519860 422632 520118
rect 423616 519860 423644 520118
rect 424628 519860 424656 520118
rect 425640 519860 425668 520118
rect 426652 519860 426680 520118
rect 427664 519860 427692 520118
rect 428676 519860 428704 520118
rect 429688 519860 429716 520118
rect 430700 519860 430728 520118
rect 431712 519860 431740 520118
rect 432724 519860 432752 520118
rect 433736 519860 433764 520118
rect 434748 519860 434776 520118
rect 435760 519860 435788 520118
rect 436772 519860 436800 520118
rect 437784 519860 437812 520118
rect 438796 519860 438824 520118
rect 439808 519860 439836 520118
rect 440820 519860 440848 520118
rect 441832 519860 441860 520118
rect 442844 519860 442872 520118
rect 443856 519860 443884 520118
rect 444868 519860 444896 520118
rect 445880 519860 445908 520118
rect 446892 519860 446920 520118
rect 447904 519860 447932 520118
rect 448916 519860 448944 520118
rect 449928 519860 449956 520118
rect 450940 519860 450968 520118
rect 451952 519860 451980 520118
rect 452964 519860 452992 520118
rect 453976 519860 454004 520118
rect 454988 519860 455016 520118
rect 456000 519860 456028 520118
rect 457012 519860 457040 520118
rect 458024 519860 458052 520118
rect 459036 519860 459064 520118
rect 460048 519860 460076 520118
rect 461060 519860 461088 520118
rect 462072 519860 462100 520118
rect 463084 519860 463112 520118
rect 464096 519860 464124 520118
rect 465108 519860 465136 520118
rect 466120 519860 466148 520118
rect 467132 519860 467160 520118
rect 468144 519860 468172 520118
rect 469156 519860 469184 520118
rect 470168 519860 470196 520118
rect 471180 519860 471208 520118
rect 472192 519860 472220 520118
rect 473204 519860 473232 520118
rect 474216 519860 474244 520118
rect 475228 519860 475256 520118
rect 476240 519860 476268 520118
rect 477252 519860 477280 520118
rect 478264 520118 478368 520146
rect 479260 520146 479288 538834
rect 479536 521626 479564 699654
rect 494808 663794 494836 703520
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 509148 700324 509200 700330
rect 509148 700266 509200 700272
rect 507766 670712 507822 670721
rect 507766 670647 507822 670656
rect 494716 663766 494836 663794
rect 489736 658028 489788 658034
rect 489736 657970 489788 657976
rect 486976 657892 487028 657898
rect 486976 657834 487028 657840
rect 485688 657076 485740 657082
rect 485688 657018 485740 657024
rect 482466 654800 482522 654809
rect 482466 654735 482522 654744
rect 479614 652080 479670 652089
rect 479614 652015 479670 652024
rect 479628 527105 479656 652015
rect 480994 650176 481050 650185
rect 480994 650111 481050 650120
rect 479708 645924 479760 645930
rect 479708 645866 479760 645872
rect 479720 536450 479748 645866
rect 480902 632632 480958 632641
rect 480902 632567 480958 632576
rect 480916 613329 480944 632567
rect 480902 613320 480958 613329
rect 480902 613255 480958 613264
rect 479708 536444 479760 536450
rect 479708 536386 479760 536392
rect 479614 527096 479670 527105
rect 479614 527031 479670 527040
rect 481008 523870 481036 650111
rect 482376 645992 482428 645998
rect 482376 645934 482428 645940
rect 482284 554124 482336 554130
rect 482284 554066 482336 554072
rect 481272 529372 481324 529378
rect 481272 529314 481324 529320
rect 480996 523864 481048 523870
rect 480996 523806 481048 523812
rect 480260 522504 480312 522510
rect 480260 522446 480312 522452
rect 479524 521620 479576 521626
rect 479524 521562 479576 521568
rect 480272 520146 480300 522446
rect 481284 520146 481312 529314
rect 481546 524376 481602 524385
rect 481546 524311 481602 524320
rect 481560 523462 481588 524311
rect 481548 523456 481600 523462
rect 481548 523398 481600 523404
rect 482296 520146 482324 554066
rect 482388 522510 482416 645934
rect 482480 530913 482508 654735
rect 485596 654424 485648 654430
rect 485596 654366 485648 654372
rect 483664 651432 483716 651438
rect 483664 651374 483716 651380
rect 482560 642116 482612 642122
rect 482560 642058 482612 642064
rect 482466 530904 482522 530913
rect 482466 530839 482522 530848
rect 482572 525366 482600 642058
rect 483296 545964 483348 545970
rect 483296 545906 483348 545912
rect 482560 525360 482612 525366
rect 482560 525302 482612 525308
rect 482376 522504 482428 522510
rect 482376 522446 482428 522452
rect 483308 520146 483336 545906
rect 483676 528154 483704 651374
rect 485042 650584 485098 650593
rect 485042 650519 485098 650528
rect 483756 646060 483808 646066
rect 483756 646002 483808 646008
rect 483768 528358 483796 646002
rect 483848 643204 483900 643210
rect 483848 643146 483900 643152
rect 483756 528352 483808 528358
rect 483756 528294 483808 528300
rect 483664 528148 483716 528154
rect 483664 528090 483716 528096
rect 483860 526658 483888 643146
rect 484308 533520 484360 533526
rect 484308 533462 484360 533468
rect 483848 526652 483900 526658
rect 483848 526594 483900 526600
rect 484320 520146 484348 533462
rect 485056 533225 485084 650519
rect 485136 636268 485188 636274
rect 485136 636210 485188 636216
rect 485042 533216 485098 533225
rect 485042 533151 485098 533160
rect 485044 533112 485096 533118
rect 485042 533080 485044 533089
rect 485096 533080 485098 533089
rect 485042 533015 485098 533024
rect 485148 526590 485176 636210
rect 485608 599826 485636 654366
rect 485700 599962 485728 657018
rect 486884 654628 486936 654634
rect 486884 654570 486936 654576
rect 486424 648780 486476 648786
rect 486424 648722 486476 648728
rect 485688 599956 485740 599962
rect 485688 599898 485740 599904
rect 485596 599820 485648 599826
rect 485596 599762 485648 599768
rect 486332 551404 486384 551410
rect 486332 551346 486384 551352
rect 485320 543108 485372 543114
rect 485320 543050 485372 543056
rect 485136 526584 485188 526590
rect 485136 526526 485188 526532
rect 485332 520146 485360 543050
rect 486344 520146 486372 551346
rect 486436 528222 486464 648722
rect 486516 636540 486568 636546
rect 486516 636482 486568 636488
rect 486528 529378 486556 636482
rect 486896 599758 486924 654570
rect 486988 599894 487016 657834
rect 488448 657416 488500 657422
rect 488448 657358 488500 657364
rect 488264 657280 488316 657286
rect 488264 657222 488316 657228
rect 488170 654528 488226 654537
rect 488170 654463 488226 654472
rect 487986 651672 488042 651681
rect 487986 651607 488042 651616
rect 487802 651536 487858 651545
rect 487802 651471 487858 651480
rect 487066 613320 487122 613329
rect 487066 613255 487122 613264
rect 486976 599888 487028 599894
rect 486976 599830 487028 599836
rect 486884 599752 486936 599758
rect 486884 599694 486936 599700
rect 487080 599593 487108 613255
rect 487066 599584 487122 599593
rect 487066 599519 487122 599528
rect 487344 532160 487396 532166
rect 487344 532102 487396 532108
rect 486516 529372 486568 529378
rect 486516 529314 486568 529320
rect 486424 528216 486476 528222
rect 486424 528158 486476 528164
rect 487356 520146 487384 532102
rect 487816 525745 487844 651471
rect 488000 528329 488028 651607
rect 488078 641200 488134 641209
rect 488078 641135 488134 641144
rect 488092 600137 488120 641135
rect 488078 600128 488134 600137
rect 488078 600063 488134 600072
rect 488184 599865 488212 654463
rect 488276 600234 488304 657222
rect 488460 654378 488488 657358
rect 489644 654492 489696 654498
rect 489644 654434 489696 654440
rect 488460 654350 488580 654378
rect 488448 654288 488500 654294
rect 488368 654236 488448 654242
rect 488368 654230 488500 654236
rect 488368 654214 488488 654230
rect 488368 600302 488396 654214
rect 488552 654134 488580 654350
rect 488460 654106 488580 654134
rect 488356 600296 488408 600302
rect 488356 600238 488408 600244
rect 488264 600228 488316 600234
rect 488264 600170 488316 600176
rect 488460 600166 488488 654106
rect 489368 640416 489420 640422
rect 489368 640358 489420 640364
rect 489184 640348 489236 640354
rect 489184 640290 489236 640296
rect 488448 600160 488500 600166
rect 488448 600102 488500 600108
rect 488170 599856 488226 599865
rect 488170 599791 488226 599800
rect 488356 537532 488408 537538
rect 488356 537474 488408 537480
rect 487986 528320 488042 528329
rect 487986 528255 488042 528264
rect 487802 525736 487858 525745
rect 487802 525671 487858 525680
rect 488368 520146 488396 537474
rect 488540 528420 488592 528426
rect 488540 528362 488592 528368
rect 488552 522918 488580 528362
rect 489196 523802 489224 640290
rect 489274 633720 489330 633729
rect 489274 633655 489330 633664
rect 489288 528554 489316 633655
rect 489380 533526 489408 640358
rect 489460 636472 489512 636478
rect 489460 636414 489512 636420
rect 489368 533520 489420 533526
rect 489368 533462 489420 533468
rect 489472 531146 489500 636414
rect 489656 600098 489684 654434
rect 489644 600092 489696 600098
rect 489644 600034 489696 600040
rect 489748 599690 489776 657970
rect 494716 657937 494744 663766
rect 501788 658028 501840 658034
rect 501788 657970 501840 657976
rect 489826 657928 489882 657937
rect 489826 657863 489882 657872
rect 494702 657928 494758 657937
rect 494702 657863 494758 657872
rect 496268 657892 496320 657898
rect 489840 600001 489868 657863
rect 491024 657824 491076 657830
rect 491024 657766 491076 657772
rect 491114 657792 491170 657801
rect 490472 657756 490524 657762
rect 490472 657698 490524 657704
rect 490380 657008 490432 657014
rect 490380 656950 490432 656956
rect 490392 654378 490420 656950
rect 490300 654350 490420 654378
rect 490300 654134 490328 654350
rect 490300 654106 490420 654134
rect 489826 599992 489882 600001
rect 489826 599927 489882 599936
rect 489736 599684 489788 599690
rect 489736 599626 489788 599632
rect 490392 581670 490420 654106
rect 490380 581664 490432 581670
rect 490380 581606 490432 581612
rect 490484 552022 490512 657698
rect 490564 657212 490616 657218
rect 490564 657154 490616 657160
rect 490472 552016 490524 552022
rect 490472 551958 490524 551964
rect 490380 536172 490432 536178
rect 490380 536114 490432 536120
rect 489460 531140 489512 531146
rect 489460 531082 489512 531088
rect 489288 528526 489592 528554
rect 489184 523796 489236 523802
rect 489184 523738 489236 523744
rect 488540 522912 488592 522918
rect 488540 522854 488592 522860
rect 489276 522708 489328 522714
rect 489276 522650 489328 522656
rect 489288 520146 489316 522650
rect 489564 520577 489592 528526
rect 489550 520568 489606 520577
rect 489550 520503 489606 520512
rect 490392 520146 490420 536114
rect 490576 522209 490604 657154
rect 491036 657014 491064 657766
rect 494716 657762 494744 657863
rect 496268 657834 496320 657840
rect 491114 657727 491170 657736
rect 491208 657756 491260 657762
rect 491128 657218 491156 657727
rect 491208 657698 491260 657704
rect 494704 657756 494756 657762
rect 494704 657698 494756 657704
rect 491116 657212 491168 657218
rect 491116 657154 491168 657160
rect 491220 657150 491248 657698
rect 493508 657416 493560 657422
rect 493508 657358 493560 657364
rect 491208 657144 491260 657150
rect 491208 657086 491260 657092
rect 491024 657008 491076 657014
rect 491024 656950 491076 656956
rect 493520 654908 493548 657358
rect 494888 657076 494940 657082
rect 494888 657018 494940 657024
rect 494900 654908 494928 657018
rect 496280 654908 496308 657834
rect 501800 654908 501828 657970
rect 507780 657393 507808 670647
rect 509160 657422 509188 700266
rect 543476 699825 543504 703520
rect 543924 700392 543976 700398
rect 543924 700334 543976 700340
rect 543462 699816 543518 699825
rect 543462 699751 543518 699760
rect 510068 657756 510120 657762
rect 510068 657698 510120 657704
rect 509148 657416 509200 657422
rect 507766 657384 507822 657393
rect 507688 657342 507766 657370
rect 503168 657280 503220 657286
rect 503168 657222 503220 657228
rect 503180 654908 503208 657222
rect 505928 655648 505980 655654
rect 505928 655590 505980 655596
rect 504548 655580 504600 655586
rect 504548 655522 504600 655528
rect 504560 654908 504588 655522
rect 505940 654908 505968 655590
rect 507688 654922 507716 657342
rect 509148 657358 509200 657364
rect 507766 657319 507822 657328
rect 509160 654922 509188 657358
rect 507334 654894 507716 654922
rect 508714 654894 509188 654922
rect 510080 654908 510108 657698
rect 516140 657688 516192 657694
rect 515586 657656 515642 657665
rect 516140 657630 516192 657636
rect 515586 657591 515642 657600
rect 511448 657212 511500 657218
rect 511448 657154 511500 657160
rect 511460 654908 511488 657154
rect 514208 657144 514260 657150
rect 515600 657121 515628 657591
rect 514208 657086 514260 657092
rect 515586 657112 515642 657121
rect 512828 657076 512880 657082
rect 512828 657018 512880 657024
rect 512840 654908 512868 657018
rect 514220 654908 514248 657086
rect 515586 657047 515642 657056
rect 515600 654908 515628 657047
rect 516152 656946 516180 657630
rect 518348 657620 518400 657626
rect 518348 657562 518400 657568
rect 516140 656940 516192 656946
rect 516140 656882 516192 656888
rect 516968 656940 517020 656946
rect 516968 656882 517020 656888
rect 516980 654908 517008 656882
rect 518360 654908 518388 657562
rect 519728 657552 519780 657558
rect 519728 657494 519780 657500
rect 521106 657520 521162 657529
rect 519740 654908 519768 657494
rect 521106 657455 521162 657464
rect 525248 657484 525300 657490
rect 521120 654908 521148 657455
rect 525248 657426 525300 657432
rect 532148 657484 532200 657490
rect 532148 657426 532200 657432
rect 522488 657348 522540 657354
rect 522488 657290 522540 657296
rect 522500 654908 522528 657290
rect 525260 654908 525288 657426
rect 526628 657348 526680 657354
rect 526628 657290 526680 657296
rect 526640 654908 526668 657290
rect 530768 657280 530820 657286
rect 530768 657222 530820 657228
rect 528008 657212 528060 657218
rect 528008 657154 528060 657160
rect 528020 654908 528048 657154
rect 529388 657144 529440 657150
rect 529388 657086 529440 657092
rect 529400 654908 529428 657086
rect 530780 654908 530808 657222
rect 532160 654908 532188 657426
rect 540980 657416 541032 657422
rect 540980 657358 541032 657364
rect 541070 657384 541126 657393
rect 537666 657248 537722 657257
rect 537666 657183 537722 657192
rect 535458 657112 535514 657121
rect 534908 657076 534960 657082
rect 535458 657047 535514 657056
rect 536286 657112 536342 657121
rect 536286 657047 536342 657056
rect 534908 657018 534960 657024
rect 533528 657008 533580 657014
rect 533528 656950 533580 656956
rect 533540 654908 533568 656950
rect 534920 654908 534948 657018
rect 535472 655625 535500 657047
rect 535458 655616 535514 655625
rect 535458 655551 535514 655560
rect 536300 654908 536328 657047
rect 537680 654908 537708 657183
rect 539046 656976 539102 656985
rect 539046 656911 539102 656920
rect 540336 656940 540388 656946
rect 539060 654908 539088 656911
rect 540336 656882 540388 656888
rect 540242 655480 540298 655489
rect 540242 655415 540298 655424
rect 498672 654634 499054 654650
rect 498660 654628 499054 654634
rect 498712 654622 499054 654628
rect 498660 654570 498712 654576
rect 523500 654560 523552 654566
rect 500406 654528 500462 654537
rect 491864 654498 492154 654514
rect 497384 654498 497674 654514
rect 491852 654492 492154 654498
rect 491904 654486 492154 654492
rect 497372 654492 497674 654498
rect 491852 654434 491904 654440
rect 497424 654486 497674 654492
rect 523552 654508 523894 654514
rect 523500 654502 523894 654508
rect 523512 654486 523894 654502
rect 500406 654463 500462 654472
rect 497372 654434 497424 654440
rect 490656 654288 490708 654294
rect 490708 654236 490774 654242
rect 490656 654230 490774 654236
rect 490668 654214 490774 654230
rect 539598 640520 539654 640529
rect 539598 640455 539654 640464
rect 539414 608696 539470 608705
rect 539414 608631 539470 608640
rect 539428 601769 539456 608631
rect 539414 601760 539470 601769
rect 539414 601695 539470 601704
rect 539506 601080 539562 601089
rect 539232 601044 539284 601050
rect 539506 601015 539562 601024
rect 539232 600986 539284 600992
rect 537298 600536 537354 600545
rect 537298 600471 537354 600480
rect 498844 600296 498896 600302
rect 498844 600238 498896 600244
rect 490760 598233 490788 600100
rect 490746 598224 490802 598233
rect 492140 598194 492168 600100
rect 493520 598262 493548 600100
rect 494900 598505 494928 600100
rect 494886 598496 494942 598505
rect 494886 598431 494942 598440
rect 493508 598256 493560 598262
rect 493508 598198 493560 598204
rect 490746 598159 490802 598168
rect 492128 598188 492180 598194
rect 492128 598130 492180 598136
rect 496280 598126 496308 600100
rect 497660 598369 497688 600100
rect 497646 598360 497702 598369
rect 497646 598295 497702 598304
rect 498752 598188 498804 598194
rect 498752 598130 498804 598136
rect 496268 598120 496320 598126
rect 496268 598062 496320 598068
rect 493324 581664 493376 581670
rect 493324 581606 493376 581612
rect 493336 568546 493364 581606
rect 493324 568540 493376 568546
rect 493324 568482 493376 568488
rect 496084 568540 496136 568546
rect 496084 568482 496136 568488
rect 496096 553586 496124 568482
rect 496084 553580 496136 553586
rect 496084 553522 496136 553528
rect 497464 553580 497516 553586
rect 497464 553522 497516 553528
rect 493324 552016 493376 552022
rect 493324 551958 493376 551964
rect 492404 548548 492456 548554
rect 492404 548490 492456 548496
rect 491300 522776 491352 522782
rect 491300 522718 491352 522724
rect 490562 522200 490618 522209
rect 490562 522135 490618 522144
rect 491312 520146 491340 522718
rect 492416 520146 492444 548490
rect 493336 545222 493364 551958
rect 496084 546780 496136 546786
rect 496084 546722 496136 546728
rect 493324 545216 493376 545222
rect 493324 545158 493376 545164
rect 496096 522714 496124 546722
rect 496176 545216 496228 545222
rect 496176 545158 496228 545164
rect 496084 522708 496136 522714
rect 496084 522650 496136 522656
rect 496188 520606 496216 545158
rect 496268 538416 496320 538422
rect 496268 538358 496320 538364
rect 496280 522646 496308 538358
rect 496728 523184 496780 523190
rect 496728 523126 496780 523132
rect 496268 522640 496320 522646
rect 496268 522582 496320 522588
rect 496740 520946 496768 523126
rect 497372 522912 497424 522918
rect 497372 522854 497424 522860
rect 496728 520940 496780 520946
rect 496728 520882 496780 520888
rect 496176 520600 496228 520606
rect 496176 520542 496228 520548
rect 497384 520169 497412 522854
rect 497476 521898 497504 553522
rect 497556 534336 497608 534342
rect 497556 534278 497608 534284
rect 497464 521892 497516 521898
rect 497464 521834 497516 521840
rect 497568 521558 497596 534278
rect 498764 528554 498792 598130
rect 498580 528526 498792 528554
rect 498200 526040 498252 526046
rect 498200 525982 498252 525988
rect 498106 521656 498162 521665
rect 498106 521591 498162 521600
rect 497556 521552 497608 521558
rect 497556 521494 497608 521500
rect 498120 520742 498148 521591
rect 498108 520736 498160 520742
rect 498108 520678 498160 520684
rect 498106 520568 498162 520577
rect 498106 520503 498162 520512
rect 498120 520470 498148 520503
rect 498016 520464 498068 520470
rect 498016 520406 498068 520412
rect 498108 520464 498160 520470
rect 498108 520406 498160 520412
rect 497370 520160 497426 520169
rect 479260 520118 479304 520146
rect 480272 520118 480316 520146
rect 481284 520118 481328 520146
rect 482296 520118 482340 520146
rect 483308 520118 483352 520146
rect 484320 520118 484364 520146
rect 485332 520118 485376 520146
rect 486344 520118 486388 520146
rect 487356 520118 487400 520146
rect 488368 520118 488412 520146
rect 489288 520118 489424 520146
rect 490392 520118 490436 520146
rect 491312 520118 491448 520146
rect 492416 520118 492460 520146
rect 478264 519860 478292 520118
rect 479276 519860 479304 520118
rect 480288 519860 480316 520118
rect 481300 519860 481328 520118
rect 482312 519860 482340 520118
rect 483324 519860 483352 520118
rect 484336 519860 484364 520118
rect 485348 519860 485376 520118
rect 486360 519860 486388 520118
rect 487372 519860 487400 520118
rect 488384 519860 488412 520118
rect 489396 519860 489424 520118
rect 490408 519860 490436 520118
rect 491420 519860 491448 520118
rect 492432 519860 492460 520118
rect 498028 520130 498056 520406
rect 498212 520266 498240 525982
rect 498580 521778 498608 528526
rect 498660 525496 498712 525502
rect 498660 525438 498712 525444
rect 498672 524634 498700 525438
rect 498672 524606 498792 524634
rect 498764 522322 498792 524606
rect 498856 524414 498884 600238
rect 510344 600228 510396 600234
rect 510344 600170 510396 600176
rect 504822 600128 504878 600137
rect 499040 598777 499068 600100
rect 499396 600024 499448 600030
rect 499396 599966 499448 599972
rect 499304 599616 499356 599622
rect 499304 599558 499356 599564
rect 499026 598768 499082 598777
rect 499026 598703 499082 598712
rect 498936 598256 498988 598262
rect 498936 598198 498988 598204
rect 498948 524906 498976 598198
rect 499120 598120 499172 598126
rect 499120 598062 499172 598068
rect 499026 550216 499082 550225
rect 499026 550151 499082 550160
rect 499040 525042 499068 550151
rect 499132 525502 499160 598062
rect 499120 525496 499172 525502
rect 499120 525438 499172 525444
rect 499040 525014 499252 525042
rect 498948 524878 499160 524906
rect 499132 524414 499160 524878
rect 498856 524386 498976 524414
rect 498764 522294 498884 522322
rect 498580 521750 498792 521778
rect 498764 521354 498792 521750
rect 498752 521348 498804 521354
rect 498752 521290 498804 521296
rect 498856 520878 498884 522294
rect 498948 521218 498976 524386
rect 499040 524386 499160 524414
rect 499040 521286 499068 524386
rect 499028 521280 499080 521286
rect 499028 521222 499080 521228
rect 498936 521212 498988 521218
rect 498936 521154 498988 521160
rect 499224 520946 499252 525014
rect 499212 520940 499264 520946
rect 499212 520882 499264 520888
rect 498844 520872 498896 520878
rect 498844 520814 498896 520820
rect 498200 520260 498252 520266
rect 498200 520202 498252 520208
rect 499316 520198 499344 599558
rect 499408 538214 499436 599966
rect 500420 598641 500448 600100
rect 500406 598632 500462 598641
rect 500406 598567 500462 598576
rect 501418 559736 501474 559745
rect 501418 559671 501474 559680
rect 500224 559360 500276 559366
rect 500224 559302 500276 559308
rect 500038 555792 500094 555801
rect 500038 555727 500094 555736
rect 499762 549944 499818 549953
rect 499762 549879 499818 549888
rect 499670 547360 499726 547369
rect 499670 547295 499726 547304
rect 499408 538186 499528 538214
rect 499304 520192 499356 520198
rect 499304 520134 499356 520140
rect 499500 520146 499528 538186
rect 499580 534200 499632 534206
rect 499578 534168 499580 534177
rect 499632 534168 499634 534177
rect 499578 534103 499634 534112
rect 499580 531480 499632 531486
rect 499578 531448 499580 531457
rect 499632 531448 499634 531457
rect 499578 531383 499634 531392
rect 499578 520160 499634 520169
rect 497370 520095 497426 520104
rect 498016 520124 498068 520130
rect 499500 520118 499578 520146
rect 499578 520095 499634 520104
rect 498016 520066 498068 520072
rect 499578 519616 499634 519625
rect 499578 519551 499634 519560
rect 60648 519046 60700 519052
rect 60556 353116 60608 353122
rect 60556 353058 60608 353064
rect 60660 347274 60688 519046
rect 60936 519042 61608 519058
rect 60924 519036 61608 519042
rect 60976 519030 61608 519036
rect 60924 518978 60976 518984
rect 499592 402974 499620 519551
rect 499684 442354 499712 547295
rect 499776 444394 499804 549879
rect 499854 543280 499910 543289
rect 499854 543215 499910 543224
rect 499868 447250 499896 543215
rect 500052 531314 500080 555727
rect 500052 531286 500172 531314
rect 499948 526176 500000 526182
rect 499948 526118 500000 526124
rect 499960 460934 499988 526118
rect 500040 523388 500092 523394
rect 500040 523330 500092 523336
rect 500052 521937 500080 523330
rect 500038 521928 500094 521937
rect 500038 521863 500094 521872
rect 500144 521812 500172 531286
rect 500236 522986 500264 559302
rect 500316 548072 500368 548078
rect 500316 548014 500368 548020
rect 500328 523666 500356 548014
rect 501142 541648 501198 541657
rect 501142 541583 501198 541592
rect 500408 539708 500460 539714
rect 500408 539650 500460 539656
rect 500316 523660 500368 523666
rect 500316 523602 500368 523608
rect 500316 523524 500368 523530
rect 500316 523466 500368 523472
rect 500224 522980 500276 522986
rect 500224 522922 500276 522928
rect 500052 521784 500172 521812
rect 500052 486130 500080 521784
rect 500132 521620 500184 521626
rect 500132 521562 500184 521568
rect 500144 521121 500172 521562
rect 500130 521112 500186 521121
rect 500130 521047 500186 521056
rect 500328 520962 500356 523466
rect 500420 523394 500448 539650
rect 500958 539472 501014 539481
rect 500958 539407 501014 539416
rect 500972 533769 501000 539407
rect 501052 538484 501104 538490
rect 501052 538426 501104 538432
rect 500958 533760 501014 533769
rect 500958 533695 501014 533704
rect 500960 529916 501012 529922
rect 500960 529858 501012 529864
rect 500972 529281 501000 529858
rect 500958 529272 501014 529281
rect 500958 529207 501014 529216
rect 500960 528624 501012 528630
rect 500958 528592 500960 528601
rect 501012 528592 501014 528601
rect 500958 528527 501014 528536
rect 500868 524680 500920 524686
rect 500868 524622 500920 524628
rect 500880 524414 500908 524622
rect 500512 524386 500908 524414
rect 500408 523388 500460 523394
rect 500408 523330 500460 523336
rect 500408 522980 500460 522986
rect 500408 522922 500460 522928
rect 500144 520934 500356 520962
rect 500040 486124 500092 486130
rect 500040 486066 500092 486072
rect 499960 460906 500080 460934
rect 499868 447222 499988 447250
rect 499856 444508 499908 444514
rect 499856 444450 499908 444456
rect 499868 444394 499896 444450
rect 499776 444366 499896 444394
rect 499960 443714 499988 447222
rect 500052 446706 500080 460906
rect 500144 451353 500172 520934
rect 500420 520724 500448 522922
rect 500236 520696 500448 520724
rect 500236 487257 500264 520696
rect 500408 520600 500460 520606
rect 500314 520568 500370 520577
rect 500408 520542 500460 520548
rect 500314 520503 500370 520512
rect 500328 520169 500356 520503
rect 500314 520160 500370 520169
rect 500314 520095 500370 520104
rect 500420 520033 500448 520542
rect 500406 520024 500462 520033
rect 500406 519959 500462 519968
rect 500316 513324 500368 513330
rect 500316 513266 500368 513272
rect 500222 487248 500278 487257
rect 500222 487183 500278 487192
rect 500222 482896 500278 482905
rect 500222 482831 500278 482840
rect 500236 474609 500264 482831
rect 500222 474600 500278 474609
rect 500222 474535 500278 474544
rect 500130 451344 500186 451353
rect 500130 451279 500186 451288
rect 500052 446678 500264 446706
rect 500130 444544 500186 444553
rect 500130 444479 500132 444488
rect 500184 444479 500186 444488
rect 500132 444450 500184 444456
rect 499960 443686 500172 443714
rect 500144 443465 500172 443686
rect 500130 443456 500186 443465
rect 500130 443391 500186 443400
rect 500130 442368 500186 442377
rect 499684 442326 500130 442354
rect 500130 442303 500186 442312
rect 500236 442105 500264 446678
rect 500222 442096 500278 442105
rect 500222 442031 500278 442040
rect 500224 441992 500276 441998
rect 500224 441934 500276 441940
rect 499592 402946 499712 402974
rect 499578 391912 499634 391921
rect 499578 391847 499634 391856
rect 62028 391672 62080 391678
rect 62028 391614 62080 391620
rect 60922 390688 60978 390697
rect 60922 390623 60978 390632
rect 60936 389065 60964 390623
rect 62040 390046 62068 391614
rect 498290 390688 498346 390697
rect 498200 390652 498252 390658
rect 499592 390674 499620 391847
rect 498290 390623 498346 390632
rect 499500 390646 499620 390674
rect 498200 390594 498252 390600
rect 323582 390416 323638 390425
rect 323582 390351 323638 390360
rect 316590 390280 316646 390289
rect 96528 390244 96580 390250
rect 96528 390186 96580 390192
rect 306288 390244 306340 390250
rect 316590 390215 316646 390224
rect 306288 390186 306340 390192
rect 62028 390040 62080 390046
rect 62028 389982 62080 389988
rect 60922 389056 60978 389065
rect 60922 388991 60978 389000
rect 66902 389056 66958 389065
rect 66902 388991 66958 389000
rect 66916 384985 66944 388991
rect 66902 384976 66958 384985
rect 66902 384911 66958 384920
rect 68388 348265 68416 390116
rect 68926 384976 68982 384985
rect 68926 384911 68982 384920
rect 68940 383654 68968 384911
rect 68940 383626 69244 383654
rect 69216 381993 69244 383626
rect 69202 381984 69258 381993
rect 69202 381919 69258 381928
rect 70136 380497 70164 390116
rect 71778 381984 71834 381993
rect 71778 381919 71834 381928
rect 70122 380488 70178 380497
rect 70122 380423 70178 380432
rect 71792 380225 71820 381919
rect 71778 380216 71834 380225
rect 71778 380151 71834 380160
rect 71884 355609 71912 390116
rect 73632 380361 73660 390116
rect 73618 380352 73674 380361
rect 73618 380287 73674 380296
rect 71870 355600 71926 355609
rect 71870 355535 71926 355544
rect 75380 351801 75408 390116
rect 77128 359689 77156 390116
rect 77574 380216 77630 380225
rect 77574 380151 77630 380160
rect 77588 377097 77616 380151
rect 77574 377088 77630 377097
rect 77574 377023 77630 377032
rect 78876 373561 78904 390116
rect 80624 384985 80652 390116
rect 80610 384976 80666 384985
rect 80610 384911 80666 384920
rect 80702 377088 80758 377097
rect 80702 377023 80758 377032
rect 78862 373552 78918 373561
rect 78862 373487 78918 373496
rect 80716 369730 80744 377023
rect 80716 369702 81480 369730
rect 81452 367713 81480 369702
rect 81438 367704 81494 367713
rect 81438 367639 81494 367648
rect 77114 359680 77170 359689
rect 77114 359615 77170 359624
rect 82372 359145 82400 390116
rect 82358 359136 82414 359145
rect 82358 359071 82414 359080
rect 75366 351792 75422 351801
rect 75366 351727 75422 351736
rect 68374 348256 68430 348265
rect 68374 348191 68430 348200
rect 71686 347848 71742 347857
rect 71686 347783 71742 347792
rect 60648 347268 60700 347274
rect 60648 347210 60700 347216
rect 62026 345128 62082 345137
rect 62026 345063 62082 345072
rect 61936 343664 61988 343670
rect 61936 343606 61988 343612
rect 60004 342916 60056 342922
rect 60004 342858 60056 342864
rect 50342 340096 50398 340105
rect 50342 340031 50398 340040
rect 49330 303240 49386 303249
rect 49330 303175 49386 303184
rect 48042 302968 48098 302977
rect 48042 302903 48098 302912
rect 46848 302388 46900 302394
rect 46848 302330 46900 302336
rect 45376 302320 45428 302326
rect 45376 302262 45428 302268
rect 38568 186992 38620 186998
rect 38568 186934 38620 186940
rect 41878 184784 41934 184793
rect 41878 184719 41934 184728
rect 37186 117872 37242 117881
rect 37186 117807 37242 117816
rect 35990 101416 36046 101425
rect 35990 101351 36046 101360
rect 35162 8936 35218 8945
rect 35162 8871 35218 8880
rect 36004 480 36032 101351
rect 37200 480 37228 117807
rect 40682 117600 40738 117609
rect 40682 117535 40738 117544
rect 38382 91896 38438 91905
rect 38382 91831 38438 91840
rect 38396 480 38424 91831
rect 39578 90400 39634 90409
rect 39578 90335 39634 90344
rect 39592 480 39620 90335
rect 40696 480 40724 117535
rect 41892 480 41920 184719
rect 44270 118008 44326 118017
rect 44270 117943 44326 117952
rect 43074 106856 43130 106865
rect 43074 106791 43130 106800
rect 43088 480 43116 106791
rect 44284 480 44312 117943
rect 45388 117298 45416 302262
rect 46756 300960 46808 300966
rect 46756 300902 46808 300908
rect 45466 185872 45522 185881
rect 45466 185807 45522 185816
rect 45376 117292 45428 117298
rect 45376 117234 45428 117240
rect 45480 480 45508 185807
rect 46768 117230 46796 300902
rect 46756 117224 46808 117230
rect 46756 117166 46808 117172
rect 46860 117065 46888 302330
rect 47950 301064 48006 301073
rect 47950 300999 48006 301008
rect 47860 300892 47912 300898
rect 47860 300834 47912 300840
rect 47584 299600 47636 299606
rect 47584 299542 47636 299548
rect 47596 267714 47624 299542
rect 47584 267708 47636 267714
rect 47584 267650 47636 267656
rect 47872 120057 47900 300834
rect 47858 120048 47914 120057
rect 47858 119983 47914 119992
rect 47964 118386 47992 300999
rect 48056 118522 48084 302903
rect 48134 302424 48190 302433
rect 48134 302359 48190 302368
rect 48044 118516 48096 118522
rect 48044 118458 48096 118464
rect 47952 118380 48004 118386
rect 47952 118322 48004 118328
rect 48148 118318 48176 302359
rect 48226 255096 48282 255105
rect 48226 255031 48282 255040
rect 48240 185065 48268 255031
rect 49344 237425 49372 303175
rect 49606 303104 49662 303113
rect 49606 303039 49662 303048
rect 49514 301200 49570 301209
rect 49514 301135 49570 301144
rect 49422 300928 49478 300937
rect 49422 300863 49478 300872
rect 49330 237416 49386 237425
rect 49330 237351 49386 237360
rect 48226 185056 48282 185065
rect 48226 184991 48282 185000
rect 48240 173233 48268 184991
rect 48226 173224 48282 173233
rect 48226 173159 48282 173168
rect 49436 120465 49464 300863
rect 49422 120456 49478 120465
rect 49422 120391 49478 120400
rect 49528 118658 49556 301135
rect 49516 118652 49568 118658
rect 49516 118594 49568 118600
rect 49620 118454 49648 303039
rect 50252 299532 50304 299538
rect 50252 299474 50304 299480
rect 50264 120086 50292 299474
rect 50356 244254 50384 340031
rect 61948 306374 61976 343606
rect 61304 306346 61976 306374
rect 50526 302832 50582 302841
rect 50526 302767 50582 302776
rect 50434 302288 50490 302297
rect 50434 302223 50490 302232
rect 50344 244248 50396 244254
rect 50344 244190 50396 244196
rect 50448 120601 50476 302223
rect 50434 120592 50490 120601
rect 50434 120527 50490 120536
rect 50252 120080 50304 120086
rect 50252 120022 50304 120028
rect 50540 118590 50568 302767
rect 57152 302388 57204 302394
rect 57152 302330 57204 302336
rect 55588 302320 55640 302326
rect 55588 302262 55640 302268
rect 53932 300960 53984 300966
rect 53932 300902 53984 300908
rect 53944 299962 53972 300902
rect 55600 299962 55628 302262
rect 57164 299962 57192 302330
rect 61304 301209 61332 306346
rect 62040 303249 62068 345063
rect 68928 341148 68980 341154
rect 68928 341090 68980 341096
rect 66076 341080 66128 341086
rect 66076 341022 66128 341028
rect 62026 303240 62082 303249
rect 62026 303175 62082 303184
rect 62040 302954 62068 303175
rect 62040 302926 62160 302954
rect 61290 301200 61346 301209
rect 61290 301135 61346 301144
rect 58900 300892 58952 300898
rect 58900 300834 58952 300840
rect 58912 299962 58940 300834
rect 61304 299962 61332 301135
rect 53944 299934 54280 299962
rect 55600 299934 55936 299962
rect 57164 299934 57592 299962
rect 58912 299934 59248 299962
rect 60904 299934 61332 299962
rect 62132 299962 62160 302926
rect 63500 302932 63552 302938
rect 63500 302874 63552 302880
rect 64328 302932 64380 302938
rect 64328 302874 64380 302880
rect 63512 302433 63540 302874
rect 63498 302424 63554 302433
rect 63498 302359 63554 302368
rect 62132 299934 62560 299962
rect 64340 299690 64368 302874
rect 66088 301073 66116 341022
rect 66168 341012 66220 341018
rect 66168 340954 66220 340960
rect 66180 303113 66208 340954
rect 66166 303104 66222 303113
rect 66166 303039 66222 303048
rect 66180 302870 66208 303039
rect 68940 302977 68968 341090
rect 71596 340944 71648 340950
rect 71596 340886 71648 340892
rect 68926 302968 68982 302977
rect 68926 302903 68982 302912
rect 66168 302864 66220 302870
rect 66168 302806 66220 302812
rect 67180 302864 67232 302870
rect 67180 302806 67232 302812
rect 68940 302818 68968 302903
rect 71608 302870 71636 340886
rect 71596 302864 71648 302870
rect 71594 302832 71596 302841
rect 71648 302832 71650 302841
rect 66074 301064 66130 301073
rect 66074 300999 66130 301008
rect 66088 299962 66116 300999
rect 65872 299934 66116 299962
rect 67192 299962 67220 302806
rect 68940 302790 69060 302818
rect 69032 299962 69060 302790
rect 71594 302767 71650 302776
rect 71700 301730 71728 347783
rect 84120 346361 84148 390116
rect 85580 387388 85632 387394
rect 85580 387330 85632 387336
rect 85592 387190 85620 387330
rect 85580 387184 85632 387190
rect 85580 387126 85632 387132
rect 85868 347721 85896 390116
rect 86868 387388 86920 387394
rect 86868 387330 86920 387336
rect 85854 347712 85910 347721
rect 85854 347647 85910 347656
rect 84106 346352 84162 346361
rect 84106 346287 84162 346296
rect 86222 321600 86278 321609
rect 86222 321535 86278 321544
rect 79416 303136 79468 303142
rect 79416 303078 79468 303084
rect 77852 303000 77904 303006
rect 75826 302968 75882 302977
rect 77852 302942 77904 302948
rect 75826 302903 75882 302912
rect 72148 302864 72200 302870
rect 72148 302806 72200 302812
rect 71240 301702 71728 301730
rect 71240 300937 71268 301702
rect 71226 300928 71282 300937
rect 71226 300863 71282 300872
rect 71240 299962 71268 300863
rect 67192 299934 67528 299962
rect 69032 299934 69184 299962
rect 70840 299934 71268 299962
rect 72160 299962 72188 302806
rect 74262 302288 74318 302297
rect 74262 302223 74318 302232
rect 72160 299934 72496 299962
rect 74276 299690 74304 302223
rect 75840 300098 75868 302903
rect 75794 300070 75868 300098
rect 75794 299948 75822 300070
rect 77864 299962 77892 302942
rect 79428 299962 79456 303078
rect 83924 303068 83976 303074
rect 83924 303010 83976 303016
rect 82728 302320 82780 302326
rect 81070 302288 81126 302297
rect 82728 302262 82780 302268
rect 81070 302223 81126 302232
rect 81084 299962 81112 302223
rect 82740 299962 82768 302262
rect 77464 299934 77892 299962
rect 79120 299934 79456 299962
rect 80776 299934 81112 299962
rect 82432 299934 82768 299962
rect 64216 299662 64368 299690
rect 74152 299662 74304 299690
rect 83936 299690 83964 303010
rect 86236 302977 86264 321535
rect 86222 302968 86278 302977
rect 86222 302903 86278 302912
rect 86880 300898 86908 387330
rect 86960 387320 87012 387326
rect 86960 387262 87012 387268
rect 86972 387122 87000 387262
rect 86960 387116 87012 387122
rect 86960 387058 87012 387064
rect 87616 346225 87644 390116
rect 88248 387320 88300 387326
rect 88248 387262 88300 387268
rect 88154 367704 88210 367713
rect 88154 367639 88210 367648
rect 88168 365809 88196 367639
rect 88154 365800 88210 365809
rect 88154 365735 88210 365744
rect 87602 346216 87658 346225
rect 87602 346151 87658 346160
rect 88260 302258 88288 387262
rect 89364 345001 89392 390116
rect 89720 387592 89772 387598
rect 89720 387534 89772 387540
rect 89628 387252 89680 387258
rect 89628 387194 89680 387200
rect 89350 344992 89406 345001
rect 89350 344927 89406 344936
rect 88984 317484 89036 317490
rect 88984 317426 89036 317432
rect 88996 303006 89024 317426
rect 88984 303000 89036 303006
rect 88984 302942 89036 302948
rect 89640 302462 89668 387194
rect 89732 387190 89760 387534
rect 89720 387184 89772 387190
rect 89720 387126 89772 387132
rect 91008 387184 91060 387190
rect 91008 387126 91060 387132
rect 90364 320884 90416 320890
rect 90364 320826 90416 320832
rect 90376 303142 90404 320826
rect 90364 303136 90416 303142
rect 90364 303078 90416 303084
rect 89628 302456 89680 302462
rect 89628 302398 89680 302404
rect 88248 302252 88300 302258
rect 88248 302194 88300 302200
rect 86132 300892 86184 300898
rect 86132 300834 86184 300840
rect 86868 300892 86920 300898
rect 86868 300834 86920 300840
rect 86144 299962 86172 300834
rect 88260 299962 88288 302194
rect 89640 299962 89668 302398
rect 91020 300966 91048 387126
rect 91112 341601 91140 390116
rect 91192 387524 91244 387530
rect 91192 387466 91244 387472
rect 91204 387122 91232 387466
rect 91192 387116 91244 387122
rect 91192 387058 91244 387064
rect 92388 387116 92440 387122
rect 92388 387058 92440 387064
rect 91098 341592 91154 341601
rect 91098 341527 91154 341536
rect 92400 302394 92428 387058
rect 92860 343641 92888 390116
rect 94502 365800 94558 365809
rect 94502 365735 94558 365744
rect 94516 350577 94544 365735
rect 94502 350568 94558 350577
rect 94502 350503 94558 350512
rect 94608 348945 94636 390116
rect 95148 388476 95200 388482
rect 95148 388418 95200 388424
rect 95160 387734 95188 388418
rect 95148 387728 95200 387734
rect 95148 387670 95200 387676
rect 94594 348936 94650 348945
rect 94594 348871 94650 348880
rect 92846 343632 92902 343641
rect 92846 343567 92902 343576
rect 95160 302802 95188 387670
rect 96356 385801 96384 390116
rect 96540 387802 96568 390186
rect 144184 390176 144236 390182
rect 306300 390130 306328 390186
rect 144184 390118 144236 390124
rect 96528 387796 96580 387802
rect 96528 387738 96580 387744
rect 96342 385792 96398 385801
rect 96342 385727 96398 385736
rect 95882 350568 95938 350577
rect 95882 350503 95938 350512
rect 95896 339425 95924 350503
rect 95882 339416 95938 339425
rect 95882 339351 95938 339360
rect 94320 302796 94372 302802
rect 94320 302738 94372 302744
rect 95148 302796 95200 302802
rect 95148 302738 95200 302744
rect 92388 302388 92440 302394
rect 92388 302330 92440 302336
rect 91008 300960 91060 300966
rect 91008 300902 91060 300908
rect 91020 299962 91048 300902
rect 92400 300234 92428 302330
rect 85744 299934 86172 299962
rect 87400 299934 88288 299962
rect 89056 299934 89668 299962
rect 90712 299934 91048 299962
rect 92354 300206 92428 300234
rect 92354 299948 92382 300206
rect 94332 299962 94360 302738
rect 95148 302320 95200 302326
rect 96540 302297 96568 387738
rect 97908 371884 97960 371890
rect 97908 371826 97960 371832
rect 97920 371278 97948 371826
rect 97908 371272 97960 371278
rect 97908 371214 97960 371220
rect 97262 339416 97318 339425
rect 97262 339351 97318 339360
rect 95148 302262 95200 302268
rect 96526 302288 96582 302297
rect 95160 301510 95188 302262
rect 96526 302223 96582 302232
rect 95148 301504 95200 301510
rect 95148 301446 95200 301452
rect 96540 299962 96568 302223
rect 97276 300121 97304 339351
rect 97920 306374 97948 371214
rect 98104 347585 98132 390116
rect 99852 349761 99880 390116
rect 99838 349752 99894 349761
rect 99838 349687 99894 349696
rect 98090 347576 98146 347585
rect 98090 347511 98146 347520
rect 101600 346089 101628 390116
rect 101586 346080 101642 346089
rect 101586 346015 101642 346024
rect 103348 343505 103376 390116
rect 105096 352753 105124 390116
rect 106188 387456 106240 387462
rect 106188 387398 106240 387404
rect 105082 352744 105138 352753
rect 105082 352679 105138 352688
rect 103334 343496 103390 343505
rect 103334 343431 103390 343440
rect 103428 340196 103480 340202
rect 103428 340138 103480 340144
rect 98642 339552 98698 339561
rect 98642 339487 98698 339496
rect 98656 319462 98684 339487
rect 98644 319456 98696 319462
rect 98644 319398 98696 319404
rect 97736 306346 97948 306374
rect 97736 300937 97764 306346
rect 98656 301034 98684 319398
rect 103440 302598 103468 340138
rect 104806 339824 104862 339833
rect 104806 339759 104862 339768
rect 102600 302592 102652 302598
rect 102600 302534 102652 302540
rect 103428 302592 103480 302598
rect 103428 302534 103480 302540
rect 100484 301096 100536 301102
rect 100484 301038 100536 301044
rect 98644 301028 98696 301034
rect 98644 300970 98696 300976
rect 97722 300928 97778 300937
rect 97722 300863 97778 300872
rect 97262 300112 97318 300121
rect 97262 300047 97318 300056
rect 97736 299962 97764 300863
rect 94024 299934 94360 299962
rect 95680 299934 96568 299962
rect 97336 299934 97764 299962
rect 98656 299962 98684 300970
rect 98656 299934 98992 299962
rect 83936 299662 84088 299690
rect 100496 299554 100524 301038
rect 102612 299962 102640 302534
rect 104820 302530 104848 339759
rect 106200 303686 106228 387398
rect 106844 365265 106872 390116
rect 106830 365256 106886 365265
rect 106830 365191 106886 365200
rect 108592 344865 108620 390116
rect 108578 344856 108634 344865
rect 108578 344791 108634 344800
rect 110340 341465 110368 390116
rect 112088 351665 112116 390116
rect 112074 351656 112130 351665
rect 112074 351591 112130 351600
rect 113836 348809 113864 390116
rect 113822 348800 113878 348809
rect 113822 348735 113878 348744
rect 110326 341456 110382 341465
rect 110326 341391 110382 341400
rect 115584 340785 115612 390116
rect 117332 343369 117360 390116
rect 119080 367713 119108 390116
rect 119066 367704 119122 367713
rect 119066 367639 119122 367648
rect 120828 366353 120856 390116
rect 122576 379273 122604 390116
rect 122562 379264 122618 379273
rect 122562 379199 122618 379208
rect 120814 366344 120870 366353
rect 120814 366279 120870 366288
rect 124324 347449 124352 390116
rect 126072 349897 126100 390116
rect 127820 370841 127848 390116
rect 129568 377641 129596 390116
rect 129554 377632 129610 377641
rect 129554 377567 129610 377576
rect 127806 370832 127862 370841
rect 127806 370767 127862 370776
rect 126058 349888 126114 349897
rect 126058 349823 126114 349832
rect 124310 347440 124366 347449
rect 124310 347375 124366 347384
rect 131316 344321 131344 390116
rect 133064 381857 133092 390116
rect 134812 386073 134840 390116
rect 134798 386064 134854 386073
rect 134798 385999 134854 386008
rect 136560 383081 136588 390116
rect 136546 383072 136602 383081
rect 136546 383007 136602 383016
rect 133050 381848 133106 381857
rect 133050 381783 133106 381792
rect 138308 345817 138336 390116
rect 140056 373833 140084 390116
rect 141804 376553 141832 390116
rect 143552 384577 143580 390116
rect 143538 384568 143594 384577
rect 143538 384503 143594 384512
rect 144196 378826 144224 390118
rect 144184 378820 144236 378826
rect 144184 378762 144236 378768
rect 141790 376544 141846 376553
rect 141790 376479 141846 376488
rect 140042 373824 140098 373833
rect 140042 373759 140098 373768
rect 138294 345808 138350 345817
rect 138294 345743 138350 345752
rect 145300 344593 145328 390116
rect 146944 378820 146996 378826
rect 146944 378762 146996 378768
rect 146956 364410 146984 378762
rect 146944 364404 146996 364410
rect 146944 364346 146996 364352
rect 145286 344584 145342 344593
rect 145286 344519 145342 344528
rect 131302 344312 131358 344321
rect 131302 344247 131358 344256
rect 125508 343732 125560 343738
rect 125508 343674 125560 343680
rect 117318 343360 117374 343369
rect 117318 343295 117374 343304
rect 115570 340776 115626 340785
rect 115570 340711 115626 340720
rect 113822 321464 113878 321473
rect 113822 321399 113878 321408
rect 106188 303680 106240 303686
rect 106188 303622 106240 303628
rect 106200 303074 106228 303622
rect 106188 303068 106240 303074
rect 106188 303010 106240 303016
rect 111800 302592 111852 302598
rect 111800 302534 111852 302540
rect 104808 302524 104860 302530
rect 104808 302466 104860 302472
rect 104820 299962 104848 302466
rect 105910 301064 105966 301073
rect 105910 300999 105966 301008
rect 105924 299962 105952 300999
rect 110326 300112 110382 300121
rect 110326 300047 110382 300056
rect 102304 299934 102640 299962
rect 103960 299934 104848 299962
rect 105616 299934 105952 299962
rect 107244 299704 107300 299713
rect 107244 299639 107300 299648
rect 52472 299538 52624 299554
rect 100312 299538 100524 299554
rect 52460 299532 52624 299538
rect 52512 299526 52624 299532
rect 100300 299532 100524 299538
rect 52460 299474 52512 299480
rect 100352 299526 100524 299532
rect 100300 299474 100352 299480
rect 100496 299418 100524 299526
rect 108900 299568 108956 299577
rect 108900 299503 108956 299512
rect 110340 299418 110368 300047
rect 100496 299390 100648 299418
rect 110340 299390 110460 299418
rect 50632 299254 50968 299282
rect 50632 120018 50660 299254
rect 110432 291825 110460 299390
rect 110418 291816 110474 291825
rect 110418 291751 110474 291760
rect 50712 244248 50764 244254
rect 50712 244190 50764 244196
rect 50724 240666 50752 244190
rect 50724 240638 50968 240666
rect 77436 240136 77492 240145
rect 52624 240094 52960 240122
rect 54280 240094 54616 240122
rect 55936 240094 56272 240122
rect 57592 240094 57836 240122
rect 52932 238105 52960 240094
rect 52918 238096 52974 238105
rect 52918 238031 52974 238040
rect 53102 237416 53158 237425
rect 53102 237351 53158 237360
rect 50620 120012 50672 120018
rect 50620 119954 50672 119960
rect 53116 119921 53144 237351
rect 54588 234569 54616 240094
rect 56244 238377 56272 240094
rect 56230 238368 56286 238377
rect 56230 238303 56286 238312
rect 57808 237969 57836 240094
rect 59234 239850 59262 240108
rect 60904 240094 61240 240122
rect 62560 240094 62896 240122
rect 64216 240094 64552 240122
rect 65872 240094 66208 240122
rect 59234 239822 59308 239850
rect 59280 238241 59308 239822
rect 59266 238232 59322 238241
rect 59266 238167 59322 238176
rect 57794 237960 57850 237969
rect 57794 237895 57850 237904
rect 61212 237425 61240 240094
rect 61198 237416 61254 237425
rect 61198 237351 61254 237360
rect 62868 237017 62896 240094
rect 62854 237008 62910 237017
rect 62854 236943 62910 236952
rect 64524 235793 64552 240094
rect 66180 238513 66208 240094
rect 67514 239850 67542 240108
rect 69184 240094 69520 240122
rect 70840 240094 71176 240122
rect 72496 240094 72832 240122
rect 74152 240094 74488 240122
rect 67514 239822 67588 239850
rect 66166 238504 66222 238513
rect 66166 238439 66222 238448
rect 64510 235784 64566 235793
rect 64510 235719 64566 235728
rect 56506 235376 56562 235385
rect 56506 235311 56562 235320
rect 54574 234560 54630 234569
rect 54574 234495 54630 234504
rect 55126 187368 55182 187377
rect 55126 187303 55182 187312
rect 54484 184952 54536 184958
rect 54484 184894 54536 184900
rect 54496 164218 54524 184894
rect 54484 164212 54536 164218
rect 54484 164154 54536 164160
rect 55140 120329 55168 187303
rect 56520 124681 56548 235311
rect 59266 232656 59322 232665
rect 59266 232591 59322 232600
rect 58622 230480 58678 230489
rect 58622 230415 58678 230424
rect 57518 202192 57574 202201
rect 57518 202127 57574 202136
rect 57426 199336 57482 199345
rect 57426 199271 57482 199280
rect 57334 185328 57390 185337
rect 57334 185263 57390 185272
rect 57150 184920 57206 184929
rect 57150 184855 57206 184864
rect 57164 144809 57192 184855
rect 57242 173224 57298 173233
rect 57242 173159 57298 173168
rect 57150 144800 57206 144809
rect 57150 144735 57206 144744
rect 56506 124672 56562 124681
rect 56506 124607 56562 124616
rect 57256 122777 57284 173159
rect 57348 128489 57376 185263
rect 57440 175273 57468 199271
rect 57532 176497 57560 202127
rect 57702 198112 57758 198121
rect 57702 198047 57758 198056
rect 57610 185464 57666 185473
rect 57610 185399 57666 185408
rect 57518 176488 57574 176497
rect 57518 176423 57574 176432
rect 57426 175264 57482 175273
rect 57426 175199 57482 175208
rect 57624 154465 57652 185399
rect 57716 158817 57744 198047
rect 57886 191176 57942 191185
rect 57886 191111 57942 191120
rect 57794 187232 57850 187241
rect 57794 187167 57850 187176
rect 57808 177993 57836 187167
rect 57900 179489 57928 191111
rect 57886 179480 57942 179489
rect 57886 179415 57942 179424
rect 57794 177984 57850 177993
rect 57794 177919 57850 177928
rect 58636 175001 58664 230415
rect 58990 196616 59046 196625
rect 58990 196551 59046 196560
rect 58898 194032 58954 194041
rect 58898 193967 58954 193976
rect 58806 185736 58862 185745
rect 58806 185671 58862 185680
rect 57886 174992 57942 175001
rect 57886 174927 57942 174936
rect 58622 174992 58678 175001
rect 58622 174927 58678 174936
rect 57900 172417 57928 174927
rect 57886 172408 57942 172417
rect 57886 172343 57942 172352
rect 57702 158808 57758 158817
rect 57702 158743 57758 158752
rect 58820 156641 58848 185671
rect 58912 162761 58940 193967
rect 58898 162752 58954 162761
rect 58898 162687 58954 162696
rect 59004 160177 59032 196551
rect 59082 192672 59138 192681
rect 59082 192607 59138 192616
rect 58990 160168 59046 160177
rect 58990 160103 59046 160112
rect 58806 156632 58862 156641
rect 58806 156567 58862 156576
rect 59096 155961 59124 192607
rect 59174 187776 59230 187785
rect 59174 187711 59230 187720
rect 59082 155952 59138 155961
rect 59082 155887 59138 155896
rect 57610 154456 57666 154465
rect 57610 154391 57666 154400
rect 57794 143440 57850 143449
rect 57794 143375 57850 143384
rect 57808 134201 57836 143375
rect 57794 134192 57850 134201
rect 57794 134127 57850 134136
rect 57334 128480 57390 128489
rect 57334 128415 57390 128424
rect 59188 126585 59216 187711
rect 59280 167113 59308 232591
rect 61382 223952 61438 223961
rect 61382 223887 61438 223896
rect 60278 221776 60334 221785
rect 60278 221711 60334 221720
rect 59910 220688 59966 220697
rect 59910 220623 59966 220632
rect 59924 182073 59952 220623
rect 60002 220144 60058 220153
rect 60002 220079 60058 220088
rect 59910 182064 59966 182073
rect 59910 181999 59966 182008
rect 59266 167104 59322 167113
rect 59266 167039 59322 167048
rect 60016 143449 60044 220079
rect 60094 217288 60150 217297
rect 60094 217223 60150 217232
rect 60002 143440 60058 143449
rect 60002 143375 60058 143384
rect 60108 132569 60136 217223
rect 60186 197976 60242 197985
rect 60186 197911 60242 197920
rect 60094 132560 60150 132569
rect 60094 132495 60150 132504
rect 60200 130937 60228 197911
rect 60292 168745 60320 221711
rect 61396 184929 61424 223887
rect 61474 222864 61530 222873
rect 61474 222799 61530 222808
rect 61488 185473 61516 222799
rect 67560 219337 67588 239822
rect 69492 237289 69520 240094
rect 69478 237280 69534 237289
rect 69478 237215 69534 237224
rect 71148 237153 71176 240094
rect 71134 237144 71190 237153
rect 71134 237079 71190 237088
rect 72804 236881 72832 240094
rect 74460 237833 74488 240094
rect 75794 239850 75822 240108
rect 88706 240136 88762 240145
rect 79120 240094 79456 240122
rect 80776 240094 81112 240122
rect 82432 240094 82768 240122
rect 77436 240071 77492 240080
rect 79428 240009 79456 240094
rect 79414 240000 79470 240009
rect 79414 239935 79470 239944
rect 75794 239822 75868 239850
rect 74446 237824 74502 237833
rect 74446 237759 74502 237768
rect 72790 236872 72846 236881
rect 72790 236807 72846 236816
rect 75840 235657 75868 239822
rect 81084 236745 81112 240094
rect 81440 238740 81492 238746
rect 81440 238682 81492 238688
rect 81452 238105 81480 238682
rect 82740 238105 82768 240094
rect 84074 239850 84102 240108
rect 85744 240094 86080 240122
rect 87400 240094 87736 240122
rect 84074 239822 84148 239850
rect 81438 238096 81494 238105
rect 81438 238031 81494 238040
rect 82726 238096 82782 238105
rect 82726 238031 82782 238040
rect 81070 236736 81126 236745
rect 81070 236671 81126 236680
rect 84120 236609 84148 239822
rect 86052 237697 86080 240094
rect 86868 238536 86920 238542
rect 86868 238478 86920 238484
rect 86880 237969 86908 238478
rect 87708 237969 87736 240094
rect 90684 240136 90740 240145
rect 89056 240094 89392 240122
rect 88706 240071 88762 240080
rect 88720 239601 88748 240071
rect 88706 239592 88762 239601
rect 88706 239527 88762 239536
rect 88984 238672 89036 238678
rect 88984 238614 89036 238620
rect 88248 238468 88300 238474
rect 88248 238410 88300 238416
rect 88260 238377 88288 238410
rect 88246 238368 88302 238377
rect 88246 238303 88302 238312
rect 88996 238241 89024 238614
rect 88982 238232 89038 238241
rect 88982 238167 89038 238176
rect 86866 237960 86922 237969
rect 86866 237895 86922 237904
rect 87694 237960 87750 237969
rect 87694 237895 87750 237904
rect 86038 237688 86094 237697
rect 86038 237623 86094 237632
rect 89364 237561 89392 240094
rect 93306 240136 93362 240145
rect 90684 240071 90740 240080
rect 92354 239873 92382 240108
rect 93306 240071 93362 240080
rect 93490 240136 93546 240145
rect 94024 240094 94360 240122
rect 95680 240094 96016 240122
rect 97336 240094 97672 240122
rect 98992 240094 99236 240122
rect 93490 240071 93546 240080
rect 93320 239873 93348 240071
rect 92340 239864 92396 239873
rect 92340 239799 92396 239808
rect 93306 239864 93362 239873
rect 93306 239799 93362 239808
rect 93504 239601 93532 240071
rect 93490 239592 93546 239601
rect 93490 239527 93546 239536
rect 94332 239465 94360 240094
rect 95988 239601 96016 240094
rect 95974 239592 96030 239601
rect 95974 239527 96030 239536
rect 94318 239456 94374 239465
rect 94318 239391 94374 239400
rect 97644 238649 97672 240094
rect 97630 238640 97686 238649
rect 97630 238575 97686 238584
rect 97908 238604 97960 238610
rect 97908 238546 97960 238552
rect 89350 237552 89406 237561
rect 89350 237487 89406 237496
rect 97920 237425 97948 238546
rect 98642 238504 98698 238513
rect 98642 238439 98698 238448
rect 98656 238134 98684 238439
rect 99208 238377 99236 240094
rect 100634 239850 100662 240108
rect 102304 240094 102640 240122
rect 103960 240094 104296 240122
rect 105616 240094 105952 240122
rect 107272 240094 107608 240122
rect 100634 239822 100708 239850
rect 100680 238513 100708 239822
rect 100666 238504 100722 238513
rect 100666 238439 100722 238448
rect 102140 238400 102192 238406
rect 99194 238368 99250 238377
rect 102140 238342 102192 238348
rect 99194 238303 99250 238312
rect 99380 238264 99432 238270
rect 99380 238206 99432 238212
rect 98644 238128 98696 238134
rect 98644 238070 98696 238076
rect 99392 237833 99420 238206
rect 102152 238105 102180 238342
rect 102612 238241 102640 240094
rect 102598 238232 102654 238241
rect 102598 238167 102654 238176
rect 104268 238105 104296 240094
rect 104808 238332 104860 238338
rect 104808 238274 104860 238280
rect 102138 238096 102194 238105
rect 102138 238031 102194 238040
rect 104254 238096 104310 238105
rect 104254 238031 104310 238040
rect 104820 237969 104848 238274
rect 105924 237969 105952 240094
rect 107580 239329 107608 240094
rect 108914 239850 108942 240108
rect 108868 239822 108942 239850
rect 107566 239320 107622 239329
rect 107566 239255 107622 239264
rect 108394 238504 108450 238513
rect 108132 238462 108394 238490
rect 108132 238377 108160 238462
rect 108394 238439 108450 238448
rect 108118 238368 108174 238377
rect 108118 238303 108174 238312
rect 106188 238196 106240 238202
rect 106188 238138 106240 238144
rect 104806 237960 104862 237969
rect 104806 237895 104862 237904
rect 105910 237960 105966 237969
rect 105910 237895 105966 237904
rect 99378 237824 99434 237833
rect 99378 237759 99434 237768
rect 106200 237697 106228 238138
rect 108304 238060 108356 238066
rect 108304 238002 108356 238008
rect 106186 237688 106242 237697
rect 106186 237623 106242 237632
rect 108316 237561 108344 238002
rect 108868 237833 108896 239822
rect 108854 237824 108910 237833
rect 108854 237759 108910 237768
rect 108302 237552 108358 237561
rect 108302 237487 108358 237496
rect 97906 237416 97962 237425
rect 97906 237351 97962 237360
rect 84106 236600 84162 236609
rect 84106 236535 84162 236544
rect 75826 235648 75882 235657
rect 75826 235583 75882 235592
rect 67546 219328 67602 219337
rect 67546 219263 67602 219272
rect 64142 215384 64198 215393
rect 64142 215319 64198 215328
rect 61474 185464 61530 185473
rect 61474 185399 61530 185408
rect 64156 185337 64184 215319
rect 102784 213988 102836 213994
rect 102784 213930 102836 213936
rect 102796 209098 102824 213930
rect 111812 209774 111840 302534
rect 112442 291816 112498 291825
rect 112442 291751 112498 291760
rect 112456 275369 112484 291751
rect 112442 275360 112498 275369
rect 112442 275295 112498 275304
rect 111720 209746 111840 209774
rect 111720 209098 111748 209746
rect 102784 209092 102836 209098
rect 102784 209034 102836 209040
rect 111708 209092 111760 209098
rect 111708 209034 111760 209040
rect 92386 187096 92442 187105
rect 92386 187031 92442 187040
rect 64142 185328 64198 185337
rect 64142 185263 64198 185272
rect 61382 184920 61438 184929
rect 92400 184892 92428 187031
rect 111720 185638 111748 209034
rect 113836 187377 113864 321399
rect 125520 320906 125548 343674
rect 147048 341873 147076 390116
rect 148796 353025 148824 390116
rect 148782 353016 148838 353025
rect 148782 352951 148838 352960
rect 150544 348673 150572 390116
rect 152292 384713 152320 390116
rect 152278 384704 152334 384713
rect 152278 384639 152334 384648
rect 154040 365401 154068 390116
rect 154026 365392 154082 365401
rect 154026 365327 154082 365336
rect 153844 364404 153896 364410
rect 153844 364346 153896 364352
rect 153856 349790 153884 364346
rect 153844 349784 153896 349790
rect 153844 349726 153896 349732
rect 150530 348664 150586 348673
rect 150530 348599 150586 348608
rect 147034 341864 147090 341873
rect 147034 341799 147090 341808
rect 155788 340649 155816 390116
rect 157536 361457 157564 390116
rect 159284 364177 159312 390116
rect 159270 364168 159326 364177
rect 159270 364103 159326 364112
rect 161032 362545 161060 390116
rect 161018 362536 161074 362545
rect 161018 362471 161074 362480
rect 157522 361448 157578 361457
rect 157522 361383 157578 361392
rect 158720 349784 158772 349790
rect 158720 349726 158772 349732
rect 158732 345370 158760 349726
rect 158720 345364 158772 345370
rect 158720 345306 158772 345312
rect 161572 345364 161624 345370
rect 161572 345306 161624 345312
rect 161584 342990 161612 345306
rect 162780 343233 162808 390116
rect 162766 343224 162822 343233
rect 162766 343159 162822 343168
rect 161572 342984 161624 342990
rect 161572 342926 161624 342932
rect 164528 341737 164556 390116
rect 166276 367985 166304 390116
rect 166262 367976 166318 367985
rect 166262 367911 166318 367920
rect 168024 366625 168052 390116
rect 169772 379409 169800 390116
rect 169758 379400 169814 379409
rect 169758 379335 169814 379344
rect 171520 375193 171548 390116
rect 171506 375184 171562 375193
rect 171506 375119 171562 375128
rect 168010 366616 168066 366625
rect 168010 366551 168066 366560
rect 173268 347041 173296 390116
rect 175016 350033 175044 390116
rect 176764 370977 176792 390116
rect 178512 375057 178540 390116
rect 180260 381993 180288 390116
rect 180246 381984 180302 381993
rect 180246 381919 180302 381928
rect 182008 378049 182036 390116
rect 183756 383353 183784 390116
rect 183742 383344 183798 383353
rect 183742 383279 183798 383288
rect 181994 378040 182050 378049
rect 181994 377975 182050 377984
rect 178498 375048 178554 375057
rect 178498 374983 178554 374992
rect 185504 372065 185532 390116
rect 185490 372056 185546 372065
rect 185490 371991 185546 372000
rect 176750 370968 176806 370977
rect 176750 370903 176806 370912
rect 175002 350024 175058 350033
rect 175002 349959 175058 349968
rect 187252 348537 187280 390116
rect 187238 348528 187294 348537
rect 187238 348463 187294 348472
rect 173254 347032 173310 347041
rect 173254 346967 173310 346976
rect 189000 345545 189028 390116
rect 188986 345536 189042 345545
rect 188986 345471 189042 345480
rect 176660 342984 176712 342990
rect 176660 342926 176712 342932
rect 164514 341728 164570 341737
rect 164514 341663 164570 341672
rect 155774 340640 155830 340649
rect 155774 340575 155830 340584
rect 176672 339454 176700 342926
rect 190748 340513 190776 390116
rect 192496 380905 192524 390116
rect 192482 380896 192538 380905
rect 192482 380831 192538 380840
rect 194244 369345 194272 390116
rect 195992 375873 196020 390116
rect 195978 375864 196034 375873
rect 195978 375799 196034 375808
rect 194230 369336 194286 369345
rect 194230 369271 194286 369280
rect 197740 344457 197768 390116
rect 199488 353161 199516 390116
rect 199474 353152 199530 353161
rect 199474 353087 199530 353096
rect 201236 351257 201264 390116
rect 202984 365673 203012 390116
rect 204732 368257 204760 390116
rect 204718 368248 204774 368257
rect 204718 368183 204774 368192
rect 202970 365664 203026 365673
rect 202970 365599 203026 365608
rect 201222 351248 201278 351257
rect 201222 351183 201278 351192
rect 197726 344448 197782 344457
rect 197726 344383 197782 344392
rect 206480 342145 206508 390116
rect 208228 361593 208256 390116
rect 209976 362953 210004 390116
rect 211724 372337 211752 390116
rect 211710 372328 211766 372337
rect 211710 372263 211766 372272
rect 213472 366761 213500 390116
rect 213458 366752 213514 366761
rect 213458 366687 213514 366696
rect 209962 362944 210018 362953
rect 209962 362879 210018 362888
rect 208214 361584 208270 361593
rect 208214 361519 208270 361528
rect 215220 354674 215248 390116
rect 216968 386209 216996 390116
rect 216954 386200 217010 386209
rect 216954 386135 217010 386144
rect 215128 354646 215248 354674
rect 211802 350704 211858 350713
rect 211802 350639 211858 350648
rect 209042 350568 209098 350577
rect 209042 350503 209098 350512
rect 206466 342136 206522 342145
rect 206466 342071 206522 342080
rect 190734 340504 190790 340513
rect 190734 340439 190790 340448
rect 176660 339448 176712 339454
rect 176660 339390 176712 339396
rect 181444 339448 181496 339454
rect 181444 339390 181496 339396
rect 125520 320890 125640 320906
rect 125520 320884 125652 320890
rect 125520 320878 125600 320884
rect 125600 320826 125652 320832
rect 124864 317416 124916 317422
rect 124864 317358 124916 317364
rect 124220 302524 124272 302530
rect 124220 302466 124272 302472
rect 113914 275360 113970 275369
rect 113914 275295 113970 275304
rect 113928 265033 113956 275295
rect 113914 265024 113970 265033
rect 113914 264959 113970 264968
rect 115202 265024 115258 265033
rect 115202 264959 115258 264968
rect 115216 242865 115244 264959
rect 115202 242856 115258 242865
rect 115202 242791 115258 242800
rect 116582 242856 116638 242865
rect 116582 242791 116638 242800
rect 116596 225049 116624 242791
rect 116582 225040 116638 225049
rect 116582 224975 116638 224984
rect 118054 225040 118110 225049
rect 118054 224975 118110 224984
rect 118068 222329 118096 224975
rect 118054 222320 118110 222329
rect 118054 222255 118110 222264
rect 122102 222184 122158 222193
rect 122102 222119 122158 222128
rect 122116 208049 122144 222119
rect 122102 208040 122158 208049
rect 122102 207975 122158 207984
rect 124126 208040 124182 208049
rect 124126 207975 124182 207984
rect 124140 204105 124168 207975
rect 124126 204096 124182 204105
rect 124126 204031 124182 204040
rect 113822 187368 113878 187377
rect 113822 187303 113878 187312
rect 111708 185632 111760 185638
rect 111708 185574 111760 185580
rect 124232 184958 124260 302466
rect 124312 302456 124364 302462
rect 124312 302398 124364 302404
rect 124220 184952 124272 184958
rect 124220 184894 124272 184900
rect 61382 184855 61438 184864
rect 60278 168736 60334 168745
rect 60278 168671 60334 168680
rect 60186 130928 60242 130937
rect 60186 130863 60242 130872
rect 59174 126576 59230 126585
rect 59174 126511 59230 126520
rect 124324 122834 124352 302398
rect 124404 184952 124456 184958
rect 124404 184894 124456 184900
rect 124232 122806 124352 122834
rect 57242 122768 57298 122777
rect 57242 122703 57298 122712
rect 57256 121553 57284 122703
rect 57242 121544 57298 121553
rect 57242 121479 57298 121488
rect 86314 120592 86370 120601
rect 86314 120527 86370 120536
rect 82818 120456 82874 120465
rect 82818 120391 82874 120400
rect 55126 120320 55182 120329
rect 55126 120255 55182 120264
rect 88062 120320 88118 120329
rect 88062 120255 88118 120264
rect 63500 120080 63552 120086
rect 61488 120020 61870 120034
rect 70398 120048 70454 120057
rect 63552 120028 63618 120034
rect 63500 120022 63618 120028
rect 63512 120020 63618 120022
rect 61488 120018 61884 120020
rect 61476 120012 61884 120018
rect 61528 120006 61884 120012
rect 63512 120006 63632 120020
rect 61476 119954 61528 119960
rect 53102 119912 53158 119921
rect 53102 119847 53158 119856
rect 50528 118584 50580 118590
rect 50528 118526 50580 118532
rect 49608 118448 49660 118454
rect 49608 118390 49660 118396
rect 48136 118312 48188 118318
rect 48136 118254 48188 118260
rect 61856 117978 61884 120006
rect 61844 117972 61896 117978
rect 61844 117914 61896 117920
rect 46846 117056 46902 117065
rect 46846 116991 46902 117000
rect 63604 115297 63632 120006
rect 65352 117230 65380 120020
rect 67114 120006 67588 120034
rect 67560 117298 67588 120006
rect 67548 117292 67600 117298
rect 67548 117234 67600 117240
rect 65340 117224 65392 117230
rect 65340 117166 65392 117172
rect 66168 117224 66220 117230
rect 66168 117166 66220 117172
rect 66180 115938 66208 117166
rect 66168 115932 66220 115938
rect 66168 115874 66220 115880
rect 67560 115870 67588 117234
rect 68848 116929 68876 120020
rect 70454 120006 70610 120034
rect 70398 119983 70454 119992
rect 72344 118658 72372 120020
rect 74092 119921 74120 120020
rect 74078 119912 74134 119921
rect 74078 119847 74134 119856
rect 72332 118652 72384 118658
rect 72332 118594 72384 118600
rect 75840 118318 75868 120020
rect 77588 118386 77616 120020
rect 79336 118454 79364 120020
rect 81084 118522 81112 120020
rect 84580 118590 84608 120020
rect 84568 118584 84620 118590
rect 84568 118526 84620 118532
rect 81072 118516 81124 118522
rect 81072 118458 81124 118464
rect 79324 118448 79376 118454
rect 79324 118390 79376 118396
rect 77576 118380 77628 118386
rect 77576 118322 77628 118328
rect 75828 118312 75880 118318
rect 75828 118254 75880 118260
rect 89824 117910 89852 120020
rect 89812 117904 89864 117910
rect 89812 117846 89864 117852
rect 91572 117842 91600 120020
rect 93320 119921 93348 120020
rect 93306 119912 93362 119921
rect 93306 119847 93362 119856
rect 95068 119785 95096 120020
rect 95054 119776 95110 119785
rect 95054 119711 95110 119720
rect 96816 119649 96844 120020
rect 96802 119640 96858 119649
rect 96802 119575 96858 119584
rect 91560 117836 91612 117842
rect 91560 117778 91612 117784
rect 98564 117065 98592 120020
rect 100312 117201 100340 120020
rect 102060 118454 102088 120020
rect 102048 118448 102100 118454
rect 102048 118390 102100 118396
rect 103808 118386 103836 120020
rect 103796 118380 103848 118386
rect 103796 118322 103848 118328
rect 105556 118250 105584 120020
rect 107304 118318 107332 120020
rect 109052 118658 109080 120020
rect 109040 118652 109092 118658
rect 109040 118594 109092 118600
rect 107292 118312 107344 118318
rect 107292 118254 107344 118260
rect 105544 118244 105596 118250
rect 105544 118186 105596 118192
rect 110800 118182 110828 120020
rect 110788 118176 110840 118182
rect 110788 118118 110840 118124
rect 112548 118114 112576 120020
rect 114296 118590 114324 120020
rect 114284 118584 114336 118590
rect 114284 118526 114336 118532
rect 116044 118522 116072 120020
rect 116032 118516 116084 118522
rect 116032 118458 116084 118464
rect 117792 118454 117820 120020
rect 117688 118448 117740 118454
rect 117688 118390 117740 118396
rect 117780 118448 117832 118454
rect 117780 118390 117832 118396
rect 112536 118108 112588 118114
rect 112536 118050 112588 118056
rect 117700 118046 117728 118390
rect 117688 118040 117740 118046
rect 117688 117982 117740 117988
rect 107568 117224 107620 117230
rect 100298 117192 100354 117201
rect 100298 117127 100354 117136
rect 106186 117192 106242 117201
rect 107568 117166 107620 117172
rect 106186 117127 106188 117136
rect 106240 117127 106242 117136
rect 106188 117098 106240 117104
rect 107580 117065 107608 117166
rect 98550 117056 98606 117065
rect 98550 116991 98606 117000
rect 107566 117056 107622 117065
rect 107566 116991 107622 117000
rect 68834 116920 68890 116929
rect 68834 116855 68890 116864
rect 106922 116512 106978 116521
rect 106922 116447 106978 116456
rect 67548 115864 67600 115870
rect 67548 115806 67600 115812
rect 63590 115288 63646 115297
rect 63590 115223 63646 115232
rect 85670 112568 85726 112577
rect 85670 112503 85726 112512
rect 46662 102776 46718 102785
rect 46662 102711 46718 102720
rect 46676 480 46704 102711
rect 65614 87952 65670 87961
rect 65536 87910 65614 87938
rect 54666 87816 54722 87825
rect 54588 87774 54666 87802
rect 52918 87000 52974 87009
rect 52918 86935 52974 86944
rect 50986 85912 51042 85921
rect 50908 85870 50986 85898
rect 50908 84810 50936 85870
rect 50986 85847 51042 85856
rect 52932 84946 52960 86935
rect 54588 84946 54616 87774
rect 54666 87751 54722 87760
rect 63866 87680 63922 87689
rect 63866 87615 63922 87624
rect 62026 87544 62082 87553
rect 62026 87479 62082 87488
rect 59266 87408 59322 87417
rect 59266 87343 59322 87352
rect 57610 87272 57666 87281
rect 57610 87207 57666 87216
rect 56230 87136 56286 87145
rect 56152 87094 56230 87122
rect 56152 84946 56180 87094
rect 56230 87071 56286 87080
rect 57624 84946 57652 87207
rect 59280 84946 59308 87343
rect 60738 87000 60794 87009
rect 60738 86935 60794 86944
rect 60752 86193 60780 86935
rect 60738 86184 60794 86193
rect 60738 86119 60794 86128
rect 60646 85776 60702 85785
rect 60646 85711 60702 85720
rect 60660 84946 60688 85711
rect 62040 85082 62068 87479
rect 52624 84918 52960 84946
rect 54188 84918 54616 84946
rect 55752 84918 56180 84946
rect 57316 84918 57652 84946
rect 58880 84918 59308 84946
rect 60444 84918 60688 84946
rect 61994 85054 62068 85082
rect 61994 84932 62022 85054
rect 63880 84946 63908 87615
rect 65536 84946 65564 87910
rect 65614 87887 65670 87896
rect 84842 87680 84898 87689
rect 84842 87615 84898 87624
rect 73068 87304 73120 87310
rect 73068 87246 73120 87252
rect 68650 86048 68706 86057
rect 68650 85983 68706 85992
rect 66994 85640 67050 85649
rect 66994 85575 67050 85584
rect 67008 84946 67036 85575
rect 68664 84946 68692 85983
rect 73080 84946 73108 87246
rect 74448 87236 74500 87242
rect 74448 87178 74500 87184
rect 74460 85762 74488 87178
rect 76472 87168 76524 87174
rect 76472 87110 76524 87116
rect 63572 84918 63908 84946
rect 65136 84918 65564 84946
rect 66700 84918 67036 84946
rect 68264 84918 68692 84946
rect 72956 84918 73108 84946
rect 74368 85734 74488 85762
rect 69800 84824 69856 84833
rect 50908 84782 51060 84810
rect 74368 84810 74396 85734
rect 76484 84946 76512 87110
rect 84016 87100 84068 87106
rect 84016 87042 84068 87048
rect 80748 85096 80804 85105
rect 80748 85031 80804 85040
rect 76084 84918 76512 84946
rect 77620 84960 77676 84969
rect 80762 84932 80790 85031
rect 84028 84946 84056 87042
rect 83904 84918 84056 84946
rect 77620 84895 77676 84904
rect 74368 84782 74520 84810
rect 69800 84759 69856 84768
rect 71364 84688 71420 84697
rect 71364 84623 71420 84632
rect 79184 84552 79240 84561
rect 79184 84487 79240 84496
rect 82312 84280 82368 84289
rect 82312 84215 82368 84224
rect 48134 81696 48190 81705
rect 48134 81631 48190 81640
rect 47674 65376 47730 65385
rect 47674 65311 47730 65320
rect 47582 62656 47638 62665
rect 47582 62591 47638 62600
rect 47490 55856 47546 55865
rect 47490 55791 47546 55800
rect 47504 18601 47532 55791
rect 47596 21321 47624 62591
rect 47688 43625 47716 65311
rect 47950 64016 48006 64025
rect 47950 63951 48006 63960
rect 47858 59936 47914 59945
rect 47858 59871 47914 59880
rect 47766 58576 47822 58585
rect 47766 58511 47822 58520
rect 47674 43616 47730 43625
rect 47674 43551 47730 43560
rect 47780 25537 47808 58511
rect 47766 25528 47822 25537
rect 47766 25463 47822 25472
rect 47872 24177 47900 59871
rect 47964 48929 47992 63951
rect 48042 61296 48098 61305
rect 48042 61231 48098 61240
rect 47950 48920 48006 48929
rect 47950 48855 48006 48864
rect 47858 24168 47914 24177
rect 47858 24103 47914 24112
rect 48056 22681 48084 61231
rect 48148 42265 48176 81631
rect 48226 80336 48282 80345
rect 48226 80271 48282 80280
rect 48240 49337 48268 80271
rect 84856 79393 84884 87615
rect 85026 87408 85082 87417
rect 85026 87343 85082 87352
rect 85040 80753 85068 87343
rect 85210 87136 85266 87145
rect 85210 87071 85266 87080
rect 85224 82113 85252 87071
rect 85210 82104 85266 82113
rect 85210 82039 85266 82048
rect 85026 80744 85082 80753
rect 85026 80679 85082 80688
rect 84842 79384 84898 79393
rect 84842 79319 84898 79328
rect 49330 78976 49386 78985
rect 49330 78911 49386 78920
rect 49238 68096 49294 68105
rect 49238 68031 49294 68040
rect 49054 66736 49110 66745
rect 49054 66671 49110 66680
rect 48226 49328 48282 49337
rect 48226 49263 48282 49272
rect 49068 49065 49096 66671
rect 49146 54496 49202 54505
rect 49146 54431 49202 54440
rect 49054 49056 49110 49065
rect 49054 48991 49110 49000
rect 48134 42256 48190 42265
rect 48134 42191 48190 42200
rect 49160 28257 49188 54431
rect 49252 39273 49280 68031
rect 49344 44849 49372 78911
rect 50250 77344 50306 77353
rect 50250 77279 50306 77288
rect 49606 76256 49662 76265
rect 49606 76191 49662 76200
rect 49514 73536 49570 73545
rect 49514 73471 49570 73480
rect 49422 70816 49478 70825
rect 49422 70751 49478 70760
rect 49330 44840 49386 44849
rect 49330 44775 49386 44784
rect 49238 39264 49294 39273
rect 49238 39199 49294 39208
rect 49436 36553 49464 70751
rect 49422 36544 49478 36553
rect 49422 36479 49478 36488
rect 49528 35193 49556 73471
rect 49514 35184 49570 35193
rect 49514 35119 49570 35128
rect 49620 30977 49648 76191
rect 50158 71904 50214 71913
rect 50158 71839 50214 71848
rect 49606 30968 49662 30977
rect 49606 30903 49662 30912
rect 49146 28248 49202 28257
rect 49146 28183 49202 28192
rect 48042 22672 48098 22681
rect 48042 22607 48098 22616
rect 47582 21312 47638 21321
rect 47582 21247 47638 21256
rect 47490 18592 47546 18601
rect 47490 18527 47546 18536
rect 50172 17241 50200 71839
rect 50264 29617 50292 77279
rect 50342 74624 50398 74633
rect 50342 74559 50398 74568
rect 50356 33833 50384 74559
rect 50434 69048 50490 69057
rect 50434 68983 50490 68992
rect 50448 37913 50476 68983
rect 50526 56672 50582 56681
rect 50526 56607 50582 56616
rect 50434 37904 50490 37913
rect 50434 37839 50490 37848
rect 50342 33824 50398 33833
rect 50342 33759 50398 33768
rect 50434 29744 50490 29753
rect 50434 29679 50490 29688
rect 50250 29608 50306 29617
rect 50250 29543 50306 29552
rect 50158 17232 50214 17241
rect 50158 17167 50214 17176
rect 48962 5128 49018 5137
rect 48962 5063 49018 5072
rect 47858 3496 47914 3505
rect 47858 3431 47914 3440
rect 47872 480 47900 3431
rect 48976 480 49004 5063
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 354 50242 480
rect 50448 354 50476 29679
rect 50540 26897 50568 56607
rect 85578 53272 85634 53281
rect 85578 53207 85634 53216
rect 50618 52592 50674 52601
rect 50618 52527 50674 52536
rect 50632 32609 50660 52527
rect 84474 51504 84530 51513
rect 84474 51439 84530 51448
rect 82082 50280 82138 50289
rect 82082 50215 82138 50224
rect 50876 50102 51028 50130
rect 52256 50102 52408 50130
rect 53636 50102 53788 50130
rect 51000 47841 51028 50102
rect 50986 47832 51042 47841
rect 50986 47767 51042 47776
rect 52380 47705 52408 50102
rect 52366 47696 52422 47705
rect 52366 47631 52422 47640
rect 53760 47569 53788 50102
rect 55002 49858 55030 50116
rect 56396 50102 56548 50130
rect 55002 49830 55076 49858
rect 53746 47560 53802 47569
rect 53746 47495 53802 47504
rect 53746 44976 53802 44985
rect 53746 44911 53802 44920
rect 51354 36680 51410 36689
rect 51354 36615 51410 36624
rect 50618 32600 50674 32609
rect 50618 32535 50674 32544
rect 50526 26888 50582 26897
rect 50526 26823 50582 26832
rect 51368 480 51396 36615
rect 51722 22944 51778 22953
rect 51722 22879 51778 22888
rect 51736 3505 51764 22879
rect 52550 10432 52606 10441
rect 52550 10367 52606 10376
rect 51722 3496 51778 3505
rect 51722 3431 51778 3440
rect 52564 480 52592 10367
rect 53760 480 53788 44911
rect 55048 19961 55076 49830
rect 56520 46345 56548 50102
rect 57762 49858 57790 50116
rect 59142 49858 59170 50116
rect 60536 50102 60688 50130
rect 57762 49830 57836 49858
rect 59142 49830 59216 49858
rect 56506 46336 56562 46345
rect 56506 46271 56562 46280
rect 55862 35320 55918 35329
rect 55862 35255 55918 35264
rect 55034 19952 55090 19961
rect 55034 19887 55090 19896
rect 55876 4049 55904 35255
rect 56046 32736 56102 32745
rect 56046 32671 56102 32680
rect 54942 4040 54998 4049
rect 54942 3975 54998 3984
rect 55862 4040 55918 4049
rect 55862 3975 55918 3984
rect 54956 480 54984 3975
rect 56060 480 56088 32671
rect 57808 8945 57836 49830
rect 58438 24304 58494 24313
rect 58438 24239 58494 24248
rect 57794 8936 57850 8945
rect 57794 8871 57850 8880
rect 57242 3224 57298 3233
rect 57242 3159 57298 3168
rect 57256 480 57284 3159
rect 58452 480 58480 24239
rect 59188 10305 59216 49830
rect 60660 47977 60688 50102
rect 61902 49858 61930 50116
rect 63282 49858 63310 50116
rect 64676 50102 64828 50130
rect 61902 49830 61976 49858
rect 63282 49830 63356 49858
rect 60646 47968 60702 47977
rect 60646 47903 60702 47912
rect 61948 13025 61976 49830
rect 62762 47968 62818 47977
rect 62762 47903 62818 47912
rect 61934 13016 61990 13025
rect 61934 12951 61990 12960
rect 62776 11665 62804 47903
rect 63328 43489 63356 49830
rect 64800 47025 64828 50102
rect 66042 49858 66070 50116
rect 67422 49858 67450 50116
rect 68802 49858 68830 50116
rect 70196 50102 70348 50130
rect 71576 50102 71728 50130
rect 66042 49830 66116 49858
rect 67422 49830 67496 49858
rect 68802 49830 68876 49858
rect 64786 47016 64842 47025
rect 64786 46951 64842 46960
rect 65614 47016 65670 47025
rect 65614 46951 65670 46960
rect 63314 43480 63370 43489
rect 63314 43415 63370 43424
rect 62854 33960 62910 33969
rect 62854 33895 62910 33904
rect 62762 11656 62818 11665
rect 62762 11591 62818 11600
rect 59174 10296 59230 10305
rect 59174 10231 59230 10240
rect 59634 7848 59690 7857
rect 59634 7783 59690 7792
rect 59648 480 59676 7783
rect 62868 3505 62896 33895
rect 65522 25664 65578 25673
rect 65522 25599 65578 25608
rect 63222 20088 63278 20097
rect 63222 20023 63278 20032
rect 62026 3496 62082 3505
rect 62026 3431 62082 3440
rect 62854 3496 62910 3505
rect 62854 3431 62910 3440
rect 60830 3360 60886 3369
rect 60830 3295 60886 3304
rect 60844 480 60872 3295
rect 62040 480 62068 3431
rect 63236 480 63264 20023
rect 64326 3632 64382 3641
rect 64326 3567 64382 3576
rect 64340 480 64368 3567
rect 65536 480 65564 25599
rect 65628 14521 65656 46951
rect 66088 42129 66116 49830
rect 66074 42120 66130 42129
rect 66074 42055 66130 42064
rect 67468 15881 67496 49830
rect 67914 49192 67970 49201
rect 67914 49127 67970 49136
rect 67454 15872 67510 15881
rect 67454 15807 67510 15816
rect 65614 14512 65670 14521
rect 65614 14447 65670 14456
rect 66718 9208 66774 9217
rect 66718 9143 66774 9152
rect 66732 480 66760 9143
rect 67928 480 67956 49127
rect 68848 40633 68876 49830
rect 70320 47818 70348 50102
rect 71700 47818 71728 50102
rect 72942 49858 72970 50116
rect 74336 50102 74488 50130
rect 75716 50102 75868 50130
rect 72942 49830 73016 49858
rect 70320 47790 71084 47818
rect 71700 47790 72464 47818
rect 68834 40624 68890 40633
rect 68834 40559 68890 40568
rect 69110 27024 69166 27033
rect 69110 26959 69166 26968
rect 69124 480 69152 26959
rect 70306 17504 70362 17513
rect 70306 17439 70362 17448
rect 70320 480 70348 17439
rect 71056 4865 71084 47790
rect 71502 22808 71558 22817
rect 71502 22743 71558 22752
rect 71042 4856 71098 4865
rect 71042 4791 71098 4800
rect 71516 480 71544 22743
rect 72436 11801 72464 47790
rect 72606 31104 72662 31113
rect 72606 31039 72662 31048
rect 72422 11792 72478 11801
rect 72422 11727 72478 11736
rect 72620 480 72648 31039
rect 72988 14657 73016 49830
rect 74460 47025 74488 50102
rect 75840 47818 75868 50102
rect 77082 49858 77110 50116
rect 78476 50102 78628 50130
rect 79856 50102 80008 50130
rect 77082 49830 77156 49858
rect 75840 47790 76604 47818
rect 74446 47016 74502 47025
rect 74446 46951 74502 46960
rect 75182 47016 75238 47025
rect 75182 46951 75238 46960
rect 74998 46200 75054 46209
rect 74998 46135 75054 46144
rect 72974 14648 73030 14657
rect 72974 14583 73030 14592
rect 73802 11928 73858 11937
rect 73802 11863 73858 11872
rect 73816 480 73844 11863
rect 75012 480 75040 46135
rect 75196 13161 75224 46951
rect 76194 28384 76250 28393
rect 76194 28319 76250 28328
rect 75182 13152 75238 13161
rect 75182 13087 75238 13096
rect 76208 480 76236 28319
rect 76576 16017 76604 47790
rect 77128 40769 77156 49830
rect 78600 47818 78628 50102
rect 79980 47818 80008 50102
rect 81222 49858 81250 50116
rect 81222 49830 81296 49858
rect 78600 47790 79364 47818
rect 79980 47790 80744 47818
rect 77114 40760 77170 40769
rect 77114 40695 77170 40704
rect 79336 18737 79364 47790
rect 80716 21457 80744 47790
rect 81268 39409 81296 49830
rect 81254 39400 81310 39409
rect 81254 39335 81310 39344
rect 80702 21448 80758 21457
rect 80702 21383 80758 21392
rect 79322 18728 79378 18737
rect 79322 18663 79378 18672
rect 76562 16008 76618 16017
rect 76562 15943 76618 15952
rect 80886 14784 80942 14793
rect 80886 14719 80942 14728
rect 77390 13288 77446 13297
rect 77390 13223 77446 13232
rect 77404 480 77432 13223
rect 79690 6488 79746 6497
rect 79690 6423 79746 6432
rect 78586 4992 78642 5001
rect 78586 4927 78642 4936
rect 78600 480 78628 4927
rect 79704 480 79732 6423
rect 80900 480 80928 14719
rect 82096 480 82124 50215
rect 82616 50102 82768 50130
rect 82740 47818 82768 50102
rect 83982 49858 84010 50116
rect 83982 49830 84056 49858
rect 82740 47790 83504 47818
rect 83278 29880 83334 29889
rect 83278 29815 83334 29824
rect 83292 480 83320 29815
rect 83476 17377 83504 47790
rect 84028 38049 84056 49830
rect 84014 38040 84070 38049
rect 84014 37975 84070 37984
rect 83462 17368 83518 17377
rect 83462 17303 83518 17312
rect 84488 480 84516 51439
rect 85592 5273 85620 53207
rect 85578 5264 85634 5273
rect 85578 5199 85634 5208
rect 85684 480 85712 112503
rect 87970 111208 88026 111217
rect 87970 111143 88026 111152
rect 86866 98968 86922 98977
rect 86866 98903 86922 98912
rect 86406 87816 86462 87825
rect 86406 87751 86462 87760
rect 86222 87272 86278 87281
rect 86222 87207 86278 87216
rect 86316 87236 86368 87242
rect 86236 51785 86264 87207
rect 86316 87178 86368 87184
rect 86328 69698 86356 87178
rect 86316 69692 86368 69698
rect 86316 69634 86368 69640
rect 86420 53145 86448 87751
rect 86406 53136 86462 53145
rect 86406 53071 86462 53080
rect 86222 51776 86278 51785
rect 86222 51711 86278 51720
rect 86880 480 86908 98903
rect 87786 87952 87842 87961
rect 87786 87887 87842 87896
rect 87602 87544 87658 87553
rect 87602 87479 87658 87488
rect 87616 7585 87644 87479
rect 87800 9081 87828 87887
rect 87786 9072 87842 9081
rect 87786 9007 87842 9016
rect 87602 7576 87658 7585
rect 87602 7511 87658 7520
rect 87984 480 88012 111143
rect 98642 108488 98698 108497
rect 98642 108423 98698 108432
rect 93950 102912 94006 102921
rect 93950 102847 94006 102856
rect 91558 101552 91614 101561
rect 91558 101487 91614 101496
rect 90362 95840 90418 95849
rect 90362 95775 90418 95784
rect 89166 72448 89222 72457
rect 89166 72383 89222 72392
rect 89180 480 89208 72383
rect 90376 480 90404 95775
rect 90548 87168 90600 87174
rect 90548 87110 90600 87116
rect 90454 62792 90510 62801
rect 90454 62727 90510 62736
rect 90468 3641 90496 62727
rect 90560 50386 90588 87110
rect 90548 50380 90600 50386
rect 90548 50322 90600 50328
rect 90454 3632 90510 3641
rect 90454 3567 90510 3576
rect 91572 480 91600 101487
rect 91744 87304 91796 87310
rect 91744 87246 91796 87252
rect 91756 54534 91784 87246
rect 91744 54528 91796 54534
rect 91744 54470 91796 54476
rect 92754 3632 92810 3641
rect 92754 3567 92810 3576
rect 92768 480 92796 3567
rect 93964 480 93992 102847
rect 97446 97336 97502 97345
rect 97446 97271 97502 97280
rect 95146 94616 95202 94625
rect 95146 94551 95202 94560
rect 95160 480 95188 94551
rect 97262 87544 97318 87553
rect 97262 87479 97318 87488
rect 96250 64152 96306 64161
rect 96250 64087 96306 64096
rect 96264 480 96292 64087
rect 97276 3641 97304 87479
rect 97262 3632 97318 3641
rect 97262 3567 97318 3576
rect 97460 480 97488 97271
rect 98656 480 98684 108423
rect 104530 105632 104586 105641
rect 104530 105567 104586 105576
rect 99838 105496 99894 105505
rect 99838 105431 99894 105440
rect 98736 87100 98788 87106
rect 98736 87042 98788 87048
rect 98748 10334 98776 87042
rect 98736 10328 98788 10334
rect 98736 10270 98788 10276
rect 99852 480 99880 105431
rect 101034 104272 101090 104281
rect 101034 104207 101090 104216
rect 101048 480 101076 104207
rect 102782 100192 102838 100201
rect 102782 100127 102838 100136
rect 102230 3632 102286 3641
rect 102230 3567 102286 3576
rect 102244 480 102272 3567
rect 102796 3505 102824 100127
rect 102782 3496 102838 3505
rect 102782 3431 102838 3440
rect 103334 3496 103390 3505
rect 103334 3431 103390 3440
rect 103348 480 103376 3431
rect 104544 480 104572 105567
rect 105542 78976 105598 78985
rect 105542 78911 105598 78920
rect 105556 55865 105584 78911
rect 105542 55856 105598 55865
rect 105542 55791 105598 55800
rect 105726 3768 105782 3777
rect 105726 3703 105782 3712
rect 105740 480 105768 3703
rect 106936 480 106964 116447
rect 119540 115569 119568 120020
rect 121288 115705 121316 120020
rect 123050 120006 123616 120034
rect 121458 118144 121514 118153
rect 121458 118079 121514 118088
rect 122286 118144 122342 118153
rect 122286 118079 122342 118088
rect 121472 117774 121500 118079
rect 121460 117768 121512 117774
rect 121460 117710 121512 117716
rect 121274 115696 121330 115705
rect 121274 115631 121330 115640
rect 119526 115560 119582 115569
rect 119526 115495 119582 115504
rect 112810 114200 112866 114209
rect 112810 114135 112866 114144
rect 110510 113792 110566 113801
rect 110510 113727 110566 113736
rect 108118 89176 108174 89185
rect 108118 89111 108174 89120
rect 108132 480 108160 89111
rect 109314 3904 109370 3913
rect 109314 3839 109370 3848
rect 109328 480 109356 3839
rect 110524 480 110552 113727
rect 111614 90536 111670 90545
rect 111614 90471 111670 90480
rect 111628 480 111656 90471
rect 112824 480 112852 114135
rect 114006 111072 114062 111081
rect 114006 111007 114062 111016
rect 114020 480 114048 111007
rect 119540 110673 119568 115495
rect 119526 110664 119582 110673
rect 119526 110599 119582 110608
rect 119894 109984 119950 109993
rect 119894 109919 119950 109928
rect 116398 103048 116454 103057
rect 116398 102983 116454 102992
rect 115202 91760 115258 91769
rect 115202 91695 115258 91704
rect 115216 480 115244 91695
rect 116412 480 116440 102983
rect 118790 93120 118846 93129
rect 118790 93055 118846 93064
rect 117594 58712 117650 58721
rect 117594 58647 117650 58656
rect 117608 480 117636 58647
rect 118804 480 118832 93055
rect 119908 480 119936 109919
rect 121090 60072 121146 60081
rect 121090 60007 121146 60016
rect 121104 480 121132 60007
rect 122300 480 122328 118079
rect 123588 115433 123616 120006
rect 124232 118046 124260 122806
rect 124416 118454 124444 184894
rect 124404 118448 124456 118454
rect 124404 118390 124456 118396
rect 124220 118040 124272 118046
rect 124220 117982 124272 117988
rect 124876 117910 124904 317358
rect 125232 118448 125284 118454
rect 125232 118390 125284 118396
rect 124864 117904 124916 117910
rect 124864 117846 124916 117852
rect 125244 115841 125272 118390
rect 125508 118040 125560 118046
rect 125508 117982 125560 117988
rect 125520 116385 125548 117982
rect 125612 117842 125640 320826
rect 178682 312488 178738 312497
rect 178682 312423 178738 312432
rect 129924 303680 129976 303686
rect 129924 303622 129976 303628
rect 126796 303000 126848 303006
rect 126796 302942 126848 302948
rect 125690 302288 125746 302297
rect 125690 302223 125746 302232
rect 125704 118658 125732 302223
rect 126808 301102 126836 302942
rect 129832 302388 129884 302394
rect 129832 302330 129884 302336
rect 126886 301608 126942 301617
rect 126886 301543 126942 301552
rect 125784 301096 125836 301102
rect 125784 301038 125836 301044
rect 126796 301096 126848 301102
rect 126796 301038 126848 301044
rect 125692 118652 125744 118658
rect 125692 118594 125744 118600
rect 125796 118590 125824 301038
rect 126900 300801 126928 301543
rect 128452 301504 128504 301510
rect 128452 301446 128504 301452
rect 128360 300960 128412 300966
rect 128360 300902 128412 300908
rect 126334 300792 126390 300801
rect 126334 300727 126390 300736
rect 126886 300792 126942 300801
rect 126886 300727 126942 300736
rect 126242 204368 126298 204377
rect 126242 204303 126298 204312
rect 125784 118584 125836 118590
rect 125784 118526 125836 118532
rect 125600 117836 125652 117842
rect 125600 117778 125652 117784
rect 125506 116376 125562 116385
rect 125506 116311 125562 116320
rect 125230 115832 125286 115841
rect 125230 115767 125286 115776
rect 123574 115424 123630 115433
rect 123574 115359 123630 115368
rect 123482 57352 123538 57361
rect 123482 57287 123538 57296
rect 123496 480 123524 57287
rect 123588 32473 123616 115359
rect 124678 61432 124734 61441
rect 124678 61367 124734 61376
rect 123574 32464 123630 32473
rect 123574 32399 123630 32408
rect 124692 480 124720 61367
rect 126256 3777 126284 204303
rect 126348 119921 126376 300727
rect 126426 205456 126482 205465
rect 126426 205391 126482 205400
rect 126334 119912 126390 119921
rect 126334 119847 126390 119856
rect 126440 3913 126468 205391
rect 126610 203280 126666 203289
rect 126610 203215 126666 203224
rect 126426 3904 126482 3913
rect 126426 3839 126482 3848
rect 126242 3768 126298 3777
rect 126242 3703 126298 3712
rect 126624 3641 126652 203215
rect 127714 141808 127770 141817
rect 127714 141743 127770 141752
rect 127622 140176 127678 140185
rect 127622 140111 127678 140120
rect 127438 132016 127494 132025
rect 127438 131951 127494 131960
rect 127346 130384 127402 130393
rect 127346 130319 127402 130328
rect 127254 127120 127310 127129
rect 127254 127055 127310 127064
rect 126980 120080 127032 120086
rect 126980 120022 127032 120028
rect 126992 119785 127020 120022
rect 126978 119776 127034 119785
rect 126978 119711 127034 119720
rect 127268 118969 127296 127055
rect 127360 120873 127388 130319
rect 127346 120864 127402 120873
rect 127346 120799 127402 120808
rect 127452 119513 127480 131951
rect 127636 120986 127664 140111
rect 127728 121145 127756 141743
rect 127898 138544 127954 138553
rect 127898 138479 127954 138488
rect 127806 128752 127862 128761
rect 127806 128687 127862 128696
rect 127714 121136 127770 121145
rect 127714 121071 127770 121080
rect 127636 120958 127756 120986
rect 127622 120048 127678 120057
rect 127622 119983 127624 119992
rect 127676 119983 127678 119992
rect 127624 119954 127676 119960
rect 127532 119944 127584 119950
rect 127532 119886 127584 119892
rect 127438 119504 127494 119513
rect 127438 119439 127494 119448
rect 127544 119377 127572 119886
rect 127530 119368 127586 119377
rect 127530 119303 127586 119312
rect 127622 119096 127678 119105
rect 127728 119082 127756 120958
rect 127820 119882 127848 128687
rect 127912 121009 127940 138479
rect 128082 135280 128138 135289
rect 128082 135215 128138 135224
rect 128096 132494 128124 135215
rect 128266 133648 128322 133657
rect 128266 133583 128322 133592
rect 128004 132466 128124 132494
rect 127898 121000 127954 121009
rect 127898 120935 127954 120944
rect 127808 119876 127860 119882
rect 127808 119818 127860 119824
rect 127808 119740 127860 119746
rect 127808 119682 127860 119688
rect 127820 119649 127848 119682
rect 128004 119649 128032 132466
rect 128082 125488 128138 125497
rect 128082 125423 128138 125432
rect 128096 119814 128124 125423
rect 128084 119808 128136 119814
rect 128084 119750 128136 119756
rect 127806 119640 127862 119649
rect 127806 119575 127862 119584
rect 127990 119640 128046 119649
rect 127990 119575 128046 119584
rect 128280 119241 128308 133583
rect 128372 132494 128400 300902
rect 128464 300830 128492 301446
rect 129740 300892 129792 300898
rect 129740 300834 129792 300840
rect 128452 300824 128504 300830
rect 128452 300766 128504 300772
rect 129004 300824 129056 300830
rect 129004 300766 129056 300772
rect 128372 132466 128584 132494
rect 128266 119232 128322 119241
rect 128266 119167 128322 119176
rect 127678 119054 127756 119082
rect 127622 119031 127678 119040
rect 127254 118960 127310 118969
rect 127254 118895 127310 118904
rect 126888 118584 126940 118590
rect 126888 118526 126940 118532
rect 126900 118046 126928 118526
rect 128556 118386 128584 132466
rect 129016 120086 129044 300766
rect 129094 204096 129150 204105
rect 129094 204031 129150 204040
rect 129108 196081 129136 204031
rect 129094 196072 129150 196081
rect 129094 196007 129150 196016
rect 129096 185632 129148 185638
rect 129096 185574 129148 185580
rect 129108 120737 129136 185574
rect 129094 120728 129150 120737
rect 129094 120663 129150 120672
rect 129004 120080 129056 120086
rect 129004 120022 129056 120028
rect 129108 118522 129136 120663
rect 129096 118516 129148 118522
rect 129096 118458 129148 118464
rect 128544 118380 128596 118386
rect 128544 118322 128596 118328
rect 126888 118040 126940 118046
rect 126888 117982 126940 117988
rect 128556 117298 128584 118322
rect 128544 117292 128596 117298
rect 128544 117234 128596 117240
rect 129752 117230 129780 300834
rect 129844 118250 129872 302330
rect 129936 120086 129964 303622
rect 132500 302660 132552 302666
rect 132500 302602 132552 302608
rect 131120 302252 131172 302258
rect 131120 302194 131172 302200
rect 130290 196072 130346 196081
rect 130290 196007 130346 196016
rect 130304 193225 130332 196007
rect 130290 193216 130346 193225
rect 130290 193151 130346 193160
rect 130382 178256 130438 178265
rect 130382 178191 130438 178200
rect 129924 120080 129976 120086
rect 129924 120022 129976 120028
rect 129936 119746 129964 120022
rect 129924 119740 129976 119746
rect 129924 119682 129976 119688
rect 129832 118244 129884 118250
rect 129832 118186 129884 118192
rect 129740 117224 129792 117230
rect 129844 117201 129872 118186
rect 129740 117166 129792 117172
rect 129830 117192 129886 117201
rect 129830 117127 129886 117136
rect 126978 116648 127034 116657
rect 126978 116583 127034 116592
rect 126610 3632 126666 3641
rect 126610 3567 126666 3576
rect 126992 480 127020 116583
rect 130396 109857 130424 178191
rect 131132 117162 131160 302194
rect 131304 301028 131356 301034
rect 131304 300970 131356 300976
rect 131210 299704 131266 299713
rect 131210 299639 131266 299648
rect 131224 118266 131252 299639
rect 131316 132494 131344 300970
rect 131486 193216 131542 193225
rect 131486 193151 131542 193160
rect 131500 184929 131528 193151
rect 131486 184920 131542 184929
rect 131486 184855 131542 184864
rect 131316 132466 131528 132494
rect 131224 118238 131344 118266
rect 131212 118108 131264 118114
rect 131212 118050 131264 118056
rect 131120 117156 131172 117162
rect 131120 117098 131172 117104
rect 131224 117065 131252 118050
rect 131210 117056 131266 117065
rect 131210 116991 131266 117000
rect 131210 115696 131266 115705
rect 131316 115682 131344 118238
rect 131500 118114 131528 132466
rect 132512 118522 132540 302602
rect 133878 301064 133934 301073
rect 133878 300999 133934 301008
rect 132590 300928 132646 300937
rect 132590 300863 132646 300872
rect 132500 118516 132552 118522
rect 132500 118458 132552 118464
rect 132604 118182 132632 300863
rect 133142 184920 133198 184929
rect 133142 184855 133198 184864
rect 133156 176769 133184 184855
rect 133142 176760 133198 176769
rect 133142 176695 133198 176704
rect 132592 118176 132644 118182
rect 132592 118118 132644 118124
rect 131488 118108 131540 118114
rect 131488 118050 131540 118056
rect 131266 115654 131344 115682
rect 131210 115631 131266 115640
rect 133892 115569 133920 300999
rect 135258 299568 135314 299577
rect 135258 299503 135314 299512
rect 134522 176760 134578 176769
rect 134522 176695 134578 176704
rect 134536 167113 134564 176695
rect 134522 167104 134578 167113
rect 134522 167039 134578 167048
rect 133878 115560 133934 115569
rect 133878 115495 133934 115504
rect 135272 115433 135300 299503
rect 175922 244624 175978 244633
rect 175922 244559 175978 244568
rect 159362 208720 159418 208729
rect 159362 208655 159418 208664
rect 155222 206544 155278 206553
rect 155222 206479 155278 206488
rect 146942 190224 146998 190233
rect 146942 190159 146998 190168
rect 140042 188048 140098 188057
rect 140042 187983 140098 187992
rect 137282 183696 137338 183705
rect 137282 183631 137338 183640
rect 136546 167104 136602 167113
rect 136546 167039 136602 167048
rect 136560 164234 136588 167039
rect 136560 164206 136680 164234
rect 136652 160177 136680 164206
rect 136638 160168 136694 160177
rect 136638 160103 136694 160112
rect 135258 115424 135314 115433
rect 135258 115359 135314 115368
rect 130382 109848 130438 109857
rect 130382 109783 130438 109792
rect 137296 91905 137324 183631
rect 138662 174992 138718 175001
rect 138662 174927 138718 174936
rect 137650 113928 137706 113937
rect 137650 113863 137706 113872
rect 137282 91896 137338 91905
rect 137282 91831 137338 91840
rect 130566 77888 130622 77897
rect 130566 77823 130622 77832
rect 130580 480 130608 77823
rect 134154 76528 134210 76537
rect 134154 76463 134210 76472
rect 134168 480 134196 76463
rect 137664 480 137692 113863
rect 138676 53281 138704 174927
rect 138662 53272 138718 53281
rect 138662 53207 138718 53216
rect 140056 10441 140084 187983
rect 141422 179344 141478 179353
rect 141422 179279 141478 179288
rect 141436 93401 141464 179279
rect 142802 176080 142858 176089
rect 142802 176015 142858 176024
rect 141422 93392 141478 93401
rect 141422 93327 141478 93336
rect 141238 93256 141294 93265
rect 141238 93191 141294 93200
rect 140042 10432 140098 10441
rect 140042 10367 140098 10376
rect 141252 480 141280 93191
rect 142816 20233 142844 176015
rect 143446 160168 143502 160177
rect 143446 160103 143502 160112
rect 143460 155961 143488 160103
rect 143446 155952 143502 155961
rect 143446 155887 143502 155896
rect 144734 109848 144790 109857
rect 144734 109783 144790 109792
rect 142802 20224 142858 20233
rect 142802 20159 142858 20168
rect 144748 480 144776 109783
rect 146956 7857 146984 190159
rect 151082 180432 151138 180441
rect 151082 180367 151138 180376
rect 147678 155952 147734 155961
rect 147678 155887 147734 155896
rect 147692 153377 147720 155887
rect 147678 153368 147734 153377
rect 147678 153303 147734 153312
rect 148322 114064 148378 114073
rect 148322 113999 148378 114008
rect 146942 7848 146998 7857
rect 146942 7783 146998 7792
rect 148336 480 148364 113999
rect 151096 16153 151124 180367
rect 155236 114209 155264 206479
rect 155222 114200 155278 114209
rect 155222 114135 155278 114144
rect 159376 109993 159404 208655
rect 175936 187241 175964 244559
rect 175922 187232 175978 187241
rect 175922 187167 175978 187176
rect 178696 157593 178724 312423
rect 181456 303686 181484 339390
rect 181444 303680 181496 303686
rect 181444 303622 181496 303628
rect 186964 303680 187016 303686
rect 186964 303622 187016 303628
rect 186976 259418 187004 303622
rect 186964 259412 187016 259418
rect 186964 259354 187016 259360
rect 189724 259412 189776 259418
rect 189724 259354 189776 259360
rect 189736 234598 189764 259354
rect 209056 239465 209084 350503
rect 209136 345228 209188 345234
rect 209136 345170 209188 345176
rect 209042 239456 209098 239465
rect 209042 239391 209098 239400
rect 209148 238134 209176 345170
rect 209228 342712 209280 342718
rect 209228 342654 209280 342660
rect 209240 238542 209268 342654
rect 209318 338600 209374 338609
rect 209318 338535 209374 338544
rect 209228 238536 209280 238542
rect 209228 238478 209280 238484
rect 209332 238474 209360 338535
rect 209320 238468 209372 238474
rect 209320 238410 209372 238416
rect 209136 238128 209188 238134
rect 209136 238070 209188 238076
rect 211816 236609 211844 350639
rect 212262 349072 212318 349081
rect 212318 349030 212396 349058
rect 212262 349007 212318 349016
rect 212264 348424 212316 348430
rect 212078 348392 212134 348401
rect 212264 348366 212316 348372
rect 212078 348327 212134 348336
rect 211894 347984 211950 347993
rect 211894 347919 211950 347928
rect 211802 236600 211858 236609
rect 211802 236535 211858 236544
rect 211908 235657 211936 347919
rect 211988 347880 212040 347886
rect 211988 347822 212040 347828
rect 212000 238270 212028 347822
rect 212092 240145 212120 348327
rect 212276 347857 212304 348366
rect 212262 347848 212318 347857
rect 212262 347783 212318 347792
rect 212170 345264 212226 345273
rect 212170 345199 212226 345208
rect 212078 240136 212134 240145
rect 212078 240071 212134 240080
rect 211988 238264 212040 238270
rect 211988 238206 212040 238212
rect 212184 237833 212212 345199
rect 212368 345014 212396 349030
rect 212446 348256 212502 348265
rect 212446 348191 212502 348200
rect 212460 348022 212488 348191
rect 212448 348016 212500 348022
rect 212448 347958 212500 347964
rect 212276 344986 212396 345014
rect 214562 344992 214618 345001
rect 212276 240009 212304 344986
rect 214562 344927 214618 344936
rect 213182 344720 213238 344729
rect 213182 344655 213238 344664
rect 212354 344040 212410 344049
rect 212354 343975 212410 343984
rect 212262 240000 212318 240009
rect 212262 239935 212318 239944
rect 212368 237969 212396 343975
rect 212446 343088 212502 343097
rect 212446 343023 212502 343032
rect 212460 239329 212488 343023
rect 212446 239320 212502 239329
rect 212446 239255 212502 239264
rect 212354 237960 212410 237969
rect 212354 237895 212410 237904
rect 212170 237824 212226 237833
rect 212170 237759 212226 237768
rect 213196 237017 213224 344655
rect 214576 343806 214604 344927
rect 214746 344176 214802 344185
rect 214746 344111 214802 344120
rect 214564 343800 214616 343806
rect 214564 343742 214616 343748
rect 214378 343632 214434 343641
rect 214378 343567 214434 343576
rect 214286 342680 214342 342689
rect 214286 342615 214342 342624
rect 214300 238513 214328 342615
rect 214392 342310 214420 343567
rect 214470 343496 214526 343505
rect 214470 343431 214526 343440
rect 214484 342582 214512 343431
rect 214654 343360 214710 343369
rect 214654 343295 214710 343304
rect 214562 343224 214618 343233
rect 214562 343159 214618 343168
rect 214576 342650 214604 343159
rect 214564 342644 214616 342650
rect 214564 342586 214616 342592
rect 214472 342576 214524 342582
rect 214472 342518 214524 342524
rect 214668 342378 214696 343295
rect 214656 342372 214708 342378
rect 214656 342314 214708 342320
rect 214380 342304 214432 342310
rect 214760 342258 214788 344111
rect 215128 343641 215156 354646
rect 217416 350804 217468 350810
rect 217416 350746 217468 350752
rect 217324 350736 217376 350742
rect 217324 350678 217376 350684
rect 216680 345704 216732 345710
rect 216680 345646 216732 345652
rect 216692 345137 216720 345646
rect 216678 345128 216734 345137
rect 216678 345063 216734 345072
rect 216678 344856 216734 344865
rect 216678 344791 216734 344800
rect 216692 344010 216720 344791
rect 216680 344004 216732 344010
rect 216680 343946 216732 343952
rect 215114 343632 215170 343641
rect 215114 343567 215170 343576
rect 214930 342408 214986 342417
rect 214930 342343 214986 342352
rect 214380 342246 214432 342252
rect 214576 342230 214788 342258
rect 214838 342272 214894 342281
rect 214286 238504 214342 238513
rect 214286 238439 214342 238448
rect 214576 238105 214604 342230
rect 214838 342207 214894 342216
rect 214654 341320 214710 341329
rect 214654 341255 214710 341264
rect 214668 239601 214696 341255
rect 214852 335354 214880 342207
rect 214760 335326 214880 335354
rect 214654 239592 214710 239601
rect 214654 239527 214710 239536
rect 214760 238241 214788 335326
rect 214944 238377 214972 342343
rect 216678 341592 216734 341601
rect 216678 341527 216680 341536
rect 216732 341527 216734 341536
rect 216680 341498 216732 341504
rect 216680 340876 216732 340882
rect 216680 340818 216732 340824
rect 216692 339833 216720 340818
rect 216864 340808 216916 340814
rect 216770 340776 216826 340785
rect 216864 340750 216916 340756
rect 216770 340711 216826 340720
rect 216678 339824 216734 339833
rect 216678 339759 216734 339768
rect 216784 339658 216812 340711
rect 216772 339652 216824 339658
rect 216772 339594 216824 339600
rect 216876 339561 216904 340750
rect 216862 339552 216918 339561
rect 216862 339487 216918 339496
rect 215114 339144 215170 339153
rect 215114 339079 215170 339088
rect 215128 238649 215156 339079
rect 215114 238640 215170 238649
rect 215114 238575 215170 238584
rect 214930 238368 214986 238377
rect 214930 238303 214986 238312
rect 214746 238232 214802 238241
rect 214746 238167 214802 238176
rect 214562 238096 214618 238105
rect 217336 238066 217364 350678
rect 217428 238202 217456 350746
rect 218716 347177 218744 390116
rect 218794 350976 218850 350985
rect 218794 350911 218850 350920
rect 218702 347168 218758 347177
rect 218702 347103 218758 347112
rect 218058 344312 218114 344321
rect 218058 344247 218114 344256
rect 218072 344146 218100 344247
rect 218060 344140 218112 344146
rect 218060 344082 218112 344088
rect 217966 341048 218022 341057
rect 217966 340983 218022 340992
rect 217782 339960 217838 339969
rect 217782 339895 217838 339904
rect 217598 339824 217654 339833
rect 217598 339759 217654 339768
rect 217508 338360 217560 338366
rect 217508 338302 217560 338308
rect 217520 238338 217548 338302
rect 217612 239737 217640 339759
rect 217796 239873 217824 339895
rect 217980 298081 218008 340983
rect 217966 298072 218022 298081
rect 217966 298007 218022 298016
rect 217782 239864 217838 239873
rect 217782 239799 217838 239808
rect 217598 239728 217654 239737
rect 217598 239663 217654 239672
rect 217508 238332 217560 238338
rect 217508 238274 217560 238280
rect 217416 238196 217468 238202
rect 217416 238138 217468 238144
rect 214562 238031 214618 238040
rect 217324 238060 217376 238066
rect 217324 238002 217376 238008
rect 213182 237008 213238 237017
rect 213182 236943 213238 236952
rect 218808 235793 218836 350911
rect 218978 350840 219034 350849
rect 218978 350775 219034 350784
rect 218992 248033 219020 350775
rect 220176 349240 220228 349246
rect 220176 349182 220228 349188
rect 220082 348120 220138 348129
rect 220082 348055 220138 348064
rect 218978 248024 219034 248033
rect 218978 247959 219034 247968
rect 220096 236745 220124 348055
rect 220188 238406 220216 349182
rect 220464 347313 220492 390116
rect 220728 390108 220780 390114
rect 220728 390050 220780 390056
rect 220740 386374 220768 390050
rect 221832 387524 221884 387530
rect 221832 387466 221884 387472
rect 220728 386368 220780 386374
rect 220728 386310 220780 386316
rect 221464 350940 221516 350946
rect 221464 350882 221516 350888
rect 220726 348936 220782 348945
rect 220726 348871 220782 348880
rect 220740 347954 220768 348871
rect 220728 347948 220780 347954
rect 220728 347890 220780 347896
rect 220726 347712 220782 347721
rect 220726 347647 220782 347656
rect 220450 347304 220506 347313
rect 220450 347239 220506 347248
rect 220740 346662 220768 347647
rect 220728 346656 220780 346662
rect 220728 346598 220780 346604
rect 220726 346352 220782 346361
rect 220726 346287 220782 346296
rect 221002 346352 221058 346361
rect 221002 346287 221058 346296
rect 220266 345944 220322 345953
rect 220266 345879 220322 345888
rect 220176 238400 220228 238406
rect 220176 238342 220228 238348
rect 220280 236881 220308 345879
rect 220740 345098 220768 346287
rect 221016 345953 221044 346287
rect 221002 345944 221058 345953
rect 221002 345879 221058 345888
rect 220728 345092 220780 345098
rect 220728 345034 220780 345040
rect 220360 342508 220412 342514
rect 220360 342450 220412 342456
rect 220372 302938 220400 342450
rect 220726 341456 220782 341465
rect 220726 341391 220782 341400
rect 220740 341222 220768 341391
rect 220728 341216 220780 341222
rect 220728 341158 220780 341164
rect 220726 340640 220782 340649
rect 220726 340575 220782 340584
rect 220740 339590 220768 340575
rect 220728 339584 220780 339590
rect 220728 339526 220780 339532
rect 220360 302932 220412 302938
rect 220360 302874 220412 302880
rect 220358 243536 220414 243545
rect 220358 243471 220414 243480
rect 220266 236872 220322 236881
rect 220266 236807 220322 236816
rect 220082 236736 220138 236745
rect 220082 236671 220138 236680
rect 218794 235784 218850 235793
rect 218794 235719 218850 235728
rect 211894 235648 211950 235657
rect 211894 235583 211950 235592
rect 189724 234592 189776 234598
rect 189724 234534 189776 234540
rect 192484 234592 192536 234598
rect 192484 234534 192536 234540
rect 192496 207058 192524 234534
rect 216126 225040 216182 225049
rect 216126 224975 216182 224984
rect 199382 209808 199438 209817
rect 199382 209743 199438 209752
rect 192484 207052 192536 207058
rect 192484 206994 192536 207000
rect 197360 207052 197412 207058
rect 197360 206994 197412 207000
rect 197372 202162 197400 206994
rect 197360 202156 197412 202162
rect 197360 202098 197412 202104
rect 188342 195664 188398 195673
rect 188342 195599 188398 195608
rect 186962 177168 187018 177177
rect 186962 177103 187018 177112
rect 178682 157584 178738 157593
rect 178682 157519 178738 157528
rect 180246 115152 180302 115161
rect 180246 115087 180302 115096
rect 176658 114472 176714 114481
rect 176658 114407 176714 114416
rect 166078 114336 166134 114345
rect 166078 114271 166134 114280
rect 162490 114200 162546 114209
rect 162490 114135 162546 114144
rect 159362 109984 159418 109993
rect 159362 109919 159418 109928
rect 155406 108352 155462 108361
rect 155406 108287 155462 108296
rect 151818 73808 151874 73817
rect 151818 73743 151874 73752
rect 151082 16144 151138 16153
rect 151082 16079 151138 16088
rect 151832 480 151860 73743
rect 155420 480 155448 108287
rect 158902 91896 158958 91905
rect 158902 91831 158958 91840
rect 158916 480 158944 91831
rect 162504 480 162532 114135
rect 166092 480 166120 114271
rect 170402 112840 170458 112849
rect 170402 112775 170458 112784
rect 170416 3641 170444 112775
rect 173162 79520 173218 79529
rect 173162 79455 173218 79464
rect 169574 3632 169630 3641
rect 169574 3567 169630 3576
rect 170402 3632 170458 3641
rect 170402 3567 170458 3576
rect 169588 480 169616 3567
rect 173176 480 173204 79455
rect 176672 480 176700 114407
rect 180260 480 180288 115087
rect 186976 112713 187004 177103
rect 186962 112704 187018 112713
rect 186962 112639 187018 112648
rect 183742 111344 183798 111353
rect 183742 111279 183798 111288
rect 183756 480 183784 111279
rect 187330 101688 187386 101697
rect 187330 101623 187386 101632
rect 187344 480 187372 101623
rect 188356 13297 188384 195599
rect 198002 186960 198058 186969
rect 198002 186895 198058 186904
rect 191746 117192 191802 117201
rect 191746 117127 191802 117136
rect 191760 117094 191788 117127
rect 191748 117088 191800 117094
rect 191748 117030 191800 117036
rect 190826 116784 190882 116793
rect 190826 116719 190882 116728
rect 188342 13288 188398 13297
rect 188342 13223 188398 13232
rect 190840 480 190868 116719
rect 195242 109984 195298 109993
rect 195242 109919 195298 109928
rect 195256 3641 195284 109919
rect 197910 107128 197966 107137
rect 197910 107063 197966 107072
rect 194414 3632 194470 3641
rect 194414 3567 194470 3576
rect 195242 3632 195298 3641
rect 195242 3567 195298 3576
rect 194428 480 194456 3567
rect 197924 480 197952 107063
rect 198016 5137 198044 186895
rect 199396 57361 199424 209743
rect 211802 207496 211858 207505
rect 211802 207431 211858 207440
rect 209042 201104 209098 201113
rect 209042 201039 209098 201048
rect 206282 191312 206338 191321
rect 206282 191247 206338 191256
rect 205086 112704 205142 112713
rect 205086 112639 205142 112648
rect 201498 94752 201554 94761
rect 201498 94687 201554 94696
rect 199382 57352 199438 57361
rect 199382 57287 199438 57296
rect 198002 5128 198058 5137
rect 198002 5063 198058 5072
rect 201512 480 201540 94687
rect 205100 480 205128 112639
rect 206296 20097 206324 191247
rect 208582 108624 208638 108633
rect 208582 108559 208638 108568
rect 206282 20088 206338 20097
rect 206282 20023 206338 20032
rect 208596 480 208624 108559
rect 209056 94625 209084 201039
rect 210422 189136 210478 189145
rect 210422 189071 210478 189080
rect 209042 94616 209098 94625
rect 209042 94551 209098 94560
rect 210436 32745 210464 189071
rect 211816 103057 211844 207431
rect 216140 198121 216168 224975
rect 216126 198112 216182 198121
rect 216126 198047 216182 198056
rect 215942 197840 215998 197849
rect 215942 197775 215998 197784
rect 214562 196752 214618 196761
rect 214562 196687 214618 196696
rect 213182 182608 213238 182617
rect 213182 182543 213238 182552
rect 212448 117020 212500 117026
rect 212448 116962 212500 116968
rect 212460 116385 212488 116962
rect 212446 116376 212502 116385
rect 212446 116311 212502 116320
rect 212170 116240 212226 116249
rect 212170 116175 212226 116184
rect 211802 103048 211858 103057
rect 211802 102983 211858 102992
rect 210422 32736 210478 32745
rect 210422 32671 210478 32680
rect 212184 480 212212 116175
rect 213196 97209 213224 182543
rect 213182 97200 213238 97209
rect 213182 97135 213238 97144
rect 214576 14793 214604 196687
rect 215666 115016 215722 115025
rect 215666 114951 215722 114960
rect 214562 14784 214618 14793
rect 214562 14719 214618 14728
rect 215680 480 215708 114951
rect 215956 51513 215984 197775
rect 220082 194576 220138 194585
rect 220082 194511 220138 194520
rect 219254 105768 219310 105777
rect 219254 105703 219310 105712
rect 215942 51504 215998 51513
rect 215942 51439 215998 51448
rect 219268 480 219296 105703
rect 220096 11937 220124 194511
rect 220372 191185 220400 243471
rect 221476 235385 221504 350882
rect 221648 349172 221700 349178
rect 221648 349114 221700 349120
rect 221554 347848 221610 347857
rect 221554 347783 221610 347792
rect 221462 235376 221518 235385
rect 221462 235311 221518 235320
rect 221568 234569 221596 347783
rect 221660 238678 221688 349114
rect 221740 342848 221792 342854
rect 221740 342790 221792 342796
rect 221752 238746 221780 342790
rect 221844 303006 221872 387466
rect 222106 351792 222162 351801
rect 222106 351727 222162 351736
rect 222014 351384 222070 351393
rect 222014 351319 222070 351328
rect 222028 345014 222056 351319
rect 222120 350606 222148 351727
rect 222108 350600 222160 350606
rect 222108 350542 222160 350548
rect 222212 350169 222240 390116
rect 223486 381712 223542 381721
rect 223486 381647 223542 381656
rect 223394 376272 223450 376281
rect 223394 376207 223450 376216
rect 222198 350160 222254 350169
rect 222198 350095 222254 350104
rect 222106 348800 222162 348809
rect 222106 348735 222162 348744
rect 222120 348090 222148 348735
rect 222108 348084 222160 348090
rect 222108 348026 222160 348032
rect 223302 347576 223358 347585
rect 223302 347511 223358 347520
rect 223316 346594 223344 347511
rect 223304 346588 223356 346594
rect 223304 346530 223356 346536
rect 223210 346216 223266 346225
rect 223210 346151 223266 346160
rect 223118 346080 223174 346089
rect 223118 346015 223174 346024
rect 223026 345944 223082 345953
rect 223026 345879 223082 345888
rect 222842 345128 222898 345137
rect 222842 345063 222898 345072
rect 222028 344986 222148 345014
rect 221924 339788 221976 339794
rect 221924 339730 221976 339736
rect 221936 339561 221964 339730
rect 222016 339720 222068 339726
rect 222014 339688 222016 339697
rect 222068 339688 222070 339697
rect 222014 339623 222070 339632
rect 221922 339552 221978 339561
rect 221922 339487 221978 339496
rect 221832 303000 221884 303006
rect 221832 302942 221884 302948
rect 222120 255377 222148 344986
rect 222106 255368 222162 255377
rect 222106 255303 222162 255312
rect 221740 238740 221792 238746
rect 221740 238682 221792 238688
rect 221648 238672 221700 238678
rect 221648 238614 221700 238620
rect 222856 237153 222884 345063
rect 223040 237289 223068 345879
rect 223132 345166 223160 346015
rect 223224 345506 223252 346151
rect 223302 345808 223358 345817
rect 223302 345743 223358 345752
rect 223212 345500 223264 345506
rect 223212 345442 223264 345448
rect 223316 345302 223344 345743
rect 223304 345296 223356 345302
rect 223304 345238 223356 345244
rect 223120 345160 223172 345166
rect 223120 345102 223172 345108
rect 223302 341864 223358 341873
rect 223302 341799 223358 341808
rect 223316 341358 223344 341799
rect 223304 341352 223356 341358
rect 223304 341294 223356 341300
rect 223408 292505 223436 376207
rect 223394 292496 223450 292505
rect 223394 292431 223450 292440
rect 223500 290329 223528 381647
rect 223960 369481 223988 390116
rect 224774 389872 224830 389881
rect 224774 389807 224830 389816
rect 223946 369472 224002 369481
rect 223946 369407 224002 369416
rect 224222 351656 224278 351665
rect 224222 351591 224278 351600
rect 224236 350878 224264 351591
rect 224682 351520 224738 351529
rect 224604 351478 224682 351506
rect 224224 350872 224276 350878
rect 224224 350814 224276 350820
rect 224222 348664 224278 348673
rect 224222 348599 224278 348608
rect 224236 347818 224264 348599
rect 224406 348256 224462 348265
rect 224328 348214 224406 348242
rect 224224 347812 224276 347818
rect 224224 347754 224276 347760
rect 224224 346724 224276 346730
rect 224224 346666 224276 346672
rect 224236 346633 224264 346666
rect 224222 346624 224278 346633
rect 224222 346559 224278 346568
rect 224222 344584 224278 344593
rect 224222 344519 224278 344528
rect 224236 343874 224264 344519
rect 224224 343868 224276 343874
rect 224224 343810 224276 343816
rect 224224 342780 224276 342786
rect 224224 342722 224276 342728
rect 224236 342553 224264 342722
rect 224222 342544 224278 342553
rect 224222 342479 224278 342488
rect 224222 340232 224278 340241
rect 224222 340167 224278 340176
rect 224236 339697 224264 340167
rect 224222 339688 224278 339697
rect 224222 339623 224278 339632
rect 224328 335354 224356 348214
rect 224406 348191 224462 348200
rect 224604 335354 224632 351478
rect 224682 351455 224738 351464
rect 224684 351008 224736 351014
rect 224684 350950 224736 350956
rect 224236 335326 224356 335354
rect 224420 335326 224632 335354
rect 223486 290320 223542 290329
rect 223486 290255 223542 290264
rect 224236 259457 224264 335326
rect 224314 326360 224370 326369
rect 224314 326295 224370 326304
rect 224222 259448 224278 259457
rect 224222 259383 224278 259392
rect 223026 237280 223082 237289
rect 223026 237215 223082 237224
rect 222842 237144 222898 237153
rect 222842 237079 222898 237088
rect 221554 234560 221610 234569
rect 221554 234495 221610 234504
rect 222842 202056 222898 202065
rect 222842 201991 222898 202000
rect 220358 191176 220414 191185
rect 220358 191111 220414 191120
rect 222750 111480 222806 111489
rect 222750 111415 222806 111424
rect 220082 11928 220138 11937
rect 220082 11863 220138 11872
rect 222764 480 222792 111415
rect 222856 108497 222884 201991
rect 224222 192400 224278 192409
rect 224222 192335 224278 192344
rect 222842 108488 222898 108497
rect 222842 108423 222898 108432
rect 224236 9217 224264 192335
rect 224328 164121 224356 326295
rect 224420 261089 224448 335326
rect 224406 261080 224462 261089
rect 224406 261015 224462 261024
rect 224696 256737 224724 350950
rect 224788 293593 224816 389807
rect 225708 387025 225736 390116
rect 225694 387016 225750 387025
rect 225694 386951 225750 386960
rect 226246 376000 226302 376009
rect 226246 375935 226302 375944
rect 226154 373280 226210 373289
rect 226154 373215 226210 373224
rect 224866 351928 224922 351937
rect 224866 351863 224922 351872
rect 224774 293584 224830 293593
rect 224774 293519 224830 293528
rect 224682 256728 224738 256737
rect 224682 256663 224738 256672
rect 224880 254017 224908 351863
rect 225050 347440 225106 347449
rect 225050 347375 225106 347384
rect 224958 347032 225014 347041
rect 224958 346967 225014 346976
rect 224972 346458 225000 346967
rect 225064 346526 225092 347375
rect 225786 347032 225842 347041
rect 225786 346967 225842 346976
rect 225052 346520 225104 346526
rect 225052 346462 225104 346468
rect 224960 346452 225012 346458
rect 224960 346394 225012 346400
rect 225800 345014 225828 346967
rect 226064 346792 226116 346798
rect 226064 346734 226116 346740
rect 225880 345772 225932 345778
rect 225880 345714 225932 345720
rect 225892 345409 225920 345714
rect 225878 345400 225934 345409
rect 225878 345335 225934 345344
rect 225800 344986 226012 345014
rect 224958 341728 225014 341737
rect 224958 341663 225014 341672
rect 224972 341494 225000 341663
rect 224960 341488 225012 341494
rect 224960 341430 225012 341436
rect 225984 289785 226012 344986
rect 225970 289776 226026 289785
rect 225970 289711 226026 289720
rect 226076 282305 226104 346734
rect 226168 299033 226196 373215
rect 226154 299024 226210 299033
rect 226154 298959 226210 298968
rect 226260 295769 226288 375935
rect 227456 364313 227484 390116
rect 227626 387968 227682 387977
rect 227626 387903 227682 387912
rect 227534 376408 227590 376417
rect 227534 376343 227590 376352
rect 227442 364304 227498 364313
rect 227442 364239 227498 364248
rect 226338 350432 226394 350441
rect 226338 350367 226340 350376
rect 226392 350367 226394 350376
rect 226340 350338 226392 350344
rect 227350 349616 227406 349625
rect 227350 349551 227406 349560
rect 227166 349480 227222 349489
rect 227166 349415 227222 349424
rect 226982 349344 227038 349353
rect 226982 349279 227038 349288
rect 226430 348528 226486 348537
rect 226430 348463 226486 348472
rect 226524 348492 226576 348498
rect 226444 348226 226472 348463
rect 226524 348434 226576 348440
rect 226432 348220 226484 348226
rect 226432 348162 226484 348168
rect 226340 348152 226392 348158
rect 226340 348094 226392 348100
rect 226352 347993 226380 348094
rect 226338 347984 226394 347993
rect 226338 347919 226394 347928
rect 226536 347857 226564 348434
rect 226522 347848 226578 347857
rect 226522 347783 226578 347792
rect 226338 345536 226394 345545
rect 226338 345471 226394 345480
rect 226352 345370 226380 345471
rect 226340 345364 226392 345370
rect 226340 345306 226392 345312
rect 226246 295760 226302 295769
rect 226246 295695 226302 295704
rect 226062 282296 226118 282305
rect 226062 282231 226118 282240
rect 226996 277409 227024 349279
rect 227074 348664 227130 348673
rect 227074 348599 227130 348608
rect 227088 283937 227116 348599
rect 227074 283928 227130 283937
rect 227074 283863 227130 283872
rect 227180 279041 227208 349415
rect 227364 292097 227392 349551
rect 227548 318753 227576 376343
rect 227534 318744 227590 318753
rect 227534 318679 227590 318688
rect 227350 292088 227406 292097
rect 227350 292023 227406 292032
rect 227166 279032 227222 279041
rect 227166 278967 227222 278976
rect 226982 277400 227038 277409
rect 226982 277335 227038 277344
rect 224866 254008 224922 254017
rect 224866 253943 224922 253952
rect 227166 240272 227222 240281
rect 227166 240207 227222 240216
rect 226064 202156 226116 202162
rect 226064 202098 226116 202104
rect 226076 194546 226104 202098
rect 227180 199345 227208 240207
rect 227166 199336 227222 199345
rect 227166 199271 227222 199280
rect 226982 198928 227038 198937
rect 226982 198863 227038 198872
rect 226064 194540 226116 194546
rect 226064 194482 226116 194488
rect 224314 164112 224370 164121
rect 224314 164047 224370 164056
rect 226996 111217 227024 198863
rect 227640 149025 227668 387903
rect 227720 386368 227772 386374
rect 227720 386310 227772 386316
rect 227732 380186 227760 386310
rect 229006 382936 229062 382945
rect 229006 382871 229062 382880
rect 227720 380180 227772 380186
rect 227720 380122 227772 380128
rect 228914 378856 228970 378865
rect 228914 378791 228970 378800
rect 228822 377360 228878 377369
rect 228822 377295 228878 377304
rect 228730 376136 228786 376145
rect 228730 376071 228786 376080
rect 227720 345840 227772 345846
rect 227720 345782 227772 345788
rect 227732 345137 227760 345782
rect 228364 345432 228416 345438
rect 228364 345374 228416 345380
rect 227718 345128 227774 345137
rect 227718 345063 227774 345072
rect 228272 343936 228324 343942
rect 228272 343878 228324 343884
rect 228284 317422 228312 343878
rect 228272 317416 228324 317422
rect 228272 317358 228324 317364
rect 228376 219337 228404 345374
rect 228456 344412 228508 344418
rect 228456 344354 228508 344360
rect 228468 238610 228496 344354
rect 228548 341420 228600 341426
rect 228548 341362 228600 341368
rect 228560 300801 228588 341362
rect 228640 338496 228692 338502
rect 228640 338438 228692 338444
rect 228652 300830 228680 338438
rect 228744 326505 228772 376071
rect 228730 326496 228786 326505
rect 228730 326431 228786 326440
rect 228836 323649 228864 377295
rect 228822 323640 228878 323649
rect 228822 323575 228878 323584
rect 228928 311137 228956 378791
rect 228914 311128 228970 311137
rect 228914 311063 228970 311072
rect 228640 300824 228692 300830
rect 228546 300792 228602 300801
rect 228640 300766 228692 300772
rect 228546 300727 228602 300736
rect 229020 291417 229048 382871
rect 229204 371113 229232 390116
rect 230386 383752 230442 383761
rect 230386 383687 230442 383696
rect 230202 381168 230258 381177
rect 230202 381103 230258 381112
rect 230110 378992 230166 379001
rect 230110 378927 230166 378936
rect 230018 375456 230074 375465
rect 230018 375391 230074 375400
rect 229190 371104 229246 371113
rect 229190 371039 229246 371048
rect 229928 351144 229980 351150
rect 229926 351112 229928 351121
rect 229980 351112 229982 351121
rect 229926 351047 229982 351056
rect 229744 345908 229796 345914
rect 229744 345850 229796 345856
rect 229006 291408 229062 291417
rect 229006 291343 229062 291352
rect 228456 238604 228508 238610
rect 228456 238546 228508 238552
rect 228362 219328 228418 219337
rect 228362 219263 228418 219272
rect 228362 200016 228418 200025
rect 228362 199951 228418 199960
rect 227626 149016 227682 149025
rect 227626 148951 227682 148960
rect 226982 111208 227038 111217
rect 226982 111143 227038 111152
rect 226338 108488 226394 108497
rect 226338 108423 226394 108432
rect 224222 9208 224278 9217
rect 224222 9143 224278 9152
rect 226352 480 226380 108423
rect 228376 101561 228404 199951
rect 229756 187105 229784 345850
rect 229926 340504 229982 340513
rect 229926 340439 229982 340448
rect 229940 339862 229968 340439
rect 229928 339856 229980 339862
rect 229928 339798 229980 339804
rect 230032 320929 230060 375391
rect 230018 320920 230074 320929
rect 230018 320855 230074 320864
rect 230124 313177 230152 378927
rect 230110 313168 230166 313177
rect 230110 313103 230166 313112
rect 230216 307737 230244 381103
rect 230296 351076 230348 351082
rect 230296 351018 230348 351024
rect 230202 307728 230258 307737
rect 230202 307663 230258 307672
rect 229834 301472 229890 301481
rect 229834 301407 229890 301416
rect 229742 187096 229798 187105
rect 229742 187031 229798 187040
rect 229848 155922 229876 301407
rect 230308 252521 230336 351018
rect 230294 252512 230350 252521
rect 230294 252447 230350 252456
rect 230400 219609 230428 383687
rect 230952 352481 230980 390116
rect 231766 387832 231822 387841
rect 231766 387767 231822 387776
rect 231674 384432 231730 384441
rect 231674 384367 231730 384376
rect 231582 384296 231638 384305
rect 231582 384231 231638 384240
rect 231490 381576 231546 381585
rect 231490 381511 231546 381520
rect 231398 381032 231454 381041
rect 231398 380967 231454 380976
rect 231306 378720 231362 378729
rect 231306 378655 231362 378664
rect 231216 376032 231268 376038
rect 231216 375974 231268 375980
rect 230938 352472 230994 352481
rect 230938 352407 230994 352416
rect 231124 344072 231176 344078
rect 231124 344014 231176 344020
rect 231136 343346 231164 344014
rect 231044 343318 231164 343346
rect 231044 335354 231072 343318
rect 231124 343256 231176 343262
rect 231124 343198 231176 343204
rect 231136 342825 231164 343198
rect 231122 342816 231178 342825
rect 231122 342751 231178 342760
rect 231124 341624 231176 341630
rect 231124 341566 231176 341572
rect 231136 341057 231164 341566
rect 231122 341048 231178 341057
rect 231122 340983 231178 340992
rect 231122 338872 231178 338881
rect 231122 338807 231178 338816
rect 231136 338502 231164 338807
rect 231124 338496 231176 338502
rect 231124 338438 231176 338444
rect 231044 335326 231164 335354
rect 231136 302841 231164 335326
rect 231228 326369 231256 375974
rect 231214 326360 231270 326369
rect 231214 326295 231270 326304
rect 231320 312225 231348 378655
rect 231306 312216 231362 312225
rect 231306 312151 231362 312160
rect 231412 306649 231440 380967
rect 231398 306640 231454 306649
rect 231398 306575 231454 306584
rect 231122 302832 231178 302841
rect 231122 302767 231178 302776
rect 231504 301209 231532 381511
rect 231490 301200 231546 301209
rect 231490 301135 231546 301144
rect 230386 219600 230442 219609
rect 230386 219535 230442 219544
rect 231596 218521 231624 384231
rect 231582 218512 231638 218521
rect 231582 218447 231638 218456
rect 231596 217705 231624 218447
rect 231582 217696 231638 217705
rect 231582 217631 231638 217640
rect 231688 217433 231716 384367
rect 231674 217424 231730 217433
rect 231674 217359 231730 217368
rect 229928 194540 229980 194546
rect 229928 194482 229980 194488
rect 229836 155916 229888 155922
rect 229836 155858 229888 155864
rect 229940 154562 229968 194482
rect 229928 154556 229980 154562
rect 229928 154498 229980 154504
rect 231780 151065 231808 387767
rect 232700 373153 232728 390116
rect 233146 388104 233202 388113
rect 233146 388039 233202 388048
rect 233054 384160 233110 384169
rect 233054 384095 233110 384104
rect 232778 383208 232834 383217
rect 232778 383143 232834 383152
rect 232686 373144 232742 373153
rect 232686 373079 232742 373088
rect 232594 367840 232650 367849
rect 232594 367775 232650 367784
rect 232504 350532 232556 350538
rect 232504 350474 232556 350480
rect 232516 317393 232544 350474
rect 232502 317384 232558 317393
rect 232502 317319 232558 317328
rect 232608 285977 232636 367775
rect 232688 348288 232740 348294
rect 232688 348230 232740 348236
rect 232594 285968 232650 285977
rect 232594 285903 232650 285912
rect 232700 255513 232728 348230
rect 232792 288153 232820 383143
rect 232962 362808 233018 362817
rect 232962 362743 233018 362752
rect 232870 359408 232926 359417
rect 232870 359343 232926 359352
rect 232778 288144 232834 288153
rect 232778 288079 232834 288088
rect 232884 256601 232912 359343
rect 232976 257689 233004 362743
rect 233068 258777 233096 384095
rect 233054 258768 233110 258777
rect 233054 258703 233110 258712
rect 232962 257680 233018 257689
rect 232962 257615 233018 257624
rect 232870 256592 232926 256601
rect 232870 256527 232926 256536
rect 232686 255504 232742 255513
rect 232686 255439 232742 255448
rect 231766 151056 231822 151065
rect 231766 150991 231822 151000
rect 233160 150113 233188 388039
rect 234342 381440 234398 381449
rect 234342 381375 234398 381384
rect 233606 378584 233662 378593
rect 233606 378519 233662 378528
rect 233620 275097 233648 378519
rect 234158 374912 234214 374921
rect 234158 374847 234214 374856
rect 233882 370696 233938 370705
rect 233882 370631 233938 370640
rect 233790 361312 233846 361321
rect 233790 361247 233846 361256
rect 233698 355872 233754 355881
rect 233698 355807 233754 355816
rect 233712 282713 233740 355807
rect 233698 282704 233754 282713
rect 233698 282639 233754 282648
rect 233804 279449 233832 361247
rect 233896 281625 233924 370631
rect 234066 369200 234122 369209
rect 234066 369135 234122 369144
rect 233976 348560 234028 348566
rect 233976 348502 234028 348508
rect 233882 281616 233938 281625
rect 233882 281551 233938 281560
rect 233790 279440 233846 279449
rect 233790 279375 233846 279384
rect 233606 275088 233662 275097
rect 233606 275023 233662 275032
rect 233988 254425 234016 348502
rect 234080 274009 234108 369135
rect 234172 278361 234200 374847
rect 234250 372192 234306 372201
rect 234250 372127 234306 372136
rect 234158 278352 234214 278361
rect 234158 278287 234214 278296
rect 234066 274000 234122 274009
rect 234066 273935 234122 273944
rect 234264 272921 234292 372127
rect 234356 277273 234384 381375
rect 234448 375329 234476 390116
rect 234618 384976 234674 384985
rect 234618 384911 234674 384920
rect 234632 383722 234660 384911
rect 235814 384840 235870 384849
rect 235814 384775 235870 384784
rect 234620 383716 234672 383722
rect 234620 383658 234672 383664
rect 235828 383654 235856 384775
rect 235828 383626 235948 383654
rect 235814 377904 235870 377913
rect 235814 377839 235870 377848
rect 235630 377768 235686 377777
rect 235630 377703 235686 377712
rect 234620 376712 234672 376718
rect 234620 376654 234672 376660
rect 234632 375465 234660 376654
rect 234618 375456 234674 375465
rect 234618 375391 234674 375400
rect 234434 375320 234490 375329
rect 234434 375255 234490 375264
rect 235538 373960 235594 373969
rect 235538 373895 235594 373904
rect 234526 368112 234582 368121
rect 234526 368047 234582 368056
rect 234342 277264 234398 277273
rect 234342 277199 234398 277208
rect 234250 272912 234306 272921
rect 234250 272847 234306 272856
rect 234540 259865 234568 368047
rect 235078 364032 235134 364041
rect 235078 363967 235134 363976
rect 235092 360194 235120 363967
rect 235446 362672 235502 362681
rect 235446 362607 235502 362616
rect 235092 360166 235212 360194
rect 235078 355192 235134 355201
rect 235000 355150 235078 355178
rect 235000 351830 235028 355150
rect 235078 355127 235134 355136
rect 235078 352880 235134 352889
rect 235078 352815 235134 352824
rect 234988 351824 235040 351830
rect 234988 351766 235040 351772
rect 234988 349308 235040 349314
rect 234988 349250 235040 349256
rect 235000 349217 235028 349250
rect 234986 349208 235042 349217
rect 234986 349143 235042 349152
rect 235092 270745 235120 352815
rect 235184 276185 235212 360166
rect 235262 353696 235318 353705
rect 235262 353631 235318 353640
rect 235170 276176 235226 276185
rect 235170 276111 235226 276120
rect 235078 270736 235134 270745
rect 235078 270671 235134 270680
rect 235276 262041 235304 353631
rect 235354 353288 235410 353297
rect 235354 353223 235410 353232
rect 235368 351966 235396 353223
rect 235356 351960 235408 351966
rect 235356 351902 235408 351908
rect 235356 351824 235408 351830
rect 235356 351766 235408 351772
rect 235262 262032 235318 262041
rect 235262 261967 235318 261976
rect 235368 260953 235396 351766
rect 235460 264217 235488 362607
rect 235552 266393 235580 373895
rect 235644 269657 235672 377703
rect 235722 376680 235778 376689
rect 235722 376615 235778 376624
rect 235630 269648 235686 269657
rect 235630 269583 235686 269592
rect 235736 267481 235764 376615
rect 235722 267472 235778 267481
rect 235722 267407 235778 267416
rect 235538 266384 235594 266393
rect 235538 266319 235594 266328
rect 235446 264208 235502 264217
rect 235446 264143 235502 264152
rect 235828 263129 235856 377839
rect 235920 265305 235948 383626
rect 236000 380180 236052 380186
rect 236000 380122 236052 380128
rect 236012 375426 236040 380122
rect 236000 375420 236052 375426
rect 236000 375362 236052 375368
rect 236196 372473 236224 390116
rect 237286 380760 237342 380769
rect 237286 380695 237342 380704
rect 236734 374640 236790 374649
rect 236734 374575 236790 374584
rect 236182 372464 236238 372473
rect 236182 372399 236238 372408
rect 236642 354240 236698 354249
rect 236642 354175 236698 354184
rect 236550 354104 236606 354113
rect 236550 354039 236606 354048
rect 235998 344448 236054 344457
rect 235998 344383 236054 344392
rect 236012 344214 236040 344383
rect 236000 344208 236052 344214
rect 236000 344150 236052 344156
rect 236366 343768 236422 343777
rect 236366 343703 236422 343712
rect 235998 342136 236054 342145
rect 235998 342071 236054 342080
rect 236012 341290 236040 342071
rect 236000 341284 236052 341290
rect 236000 341226 236052 341232
rect 235906 265296 235962 265305
rect 235906 265231 235962 265240
rect 235814 263120 235870 263129
rect 235814 263055 235870 263064
rect 235354 260944 235410 260953
rect 235354 260879 235410 260888
rect 234526 259856 234582 259865
rect 234526 259791 234582 259800
rect 233974 254416 234030 254425
rect 233974 254351 234030 254360
rect 236380 253337 236408 343703
rect 236564 303385 236592 354039
rect 236550 303376 236606 303385
rect 236550 303311 236606 303320
rect 236656 302297 236684 354175
rect 236748 319841 236776 374575
rect 236826 372736 236882 372745
rect 236826 372671 236882 372680
rect 236734 319832 236790 319841
rect 236734 319767 236790 319776
rect 236840 305561 236868 372671
rect 237194 365528 237250 365537
rect 237194 365463 237250 365472
rect 237102 355056 237158 355065
rect 236932 355014 237102 355042
rect 236932 350534 236960 355014
rect 237102 354991 237158 355000
rect 237010 354512 237066 354521
rect 237010 354447 237066 354456
rect 237024 353326 237052 354447
rect 237102 354376 237158 354385
rect 237102 354311 237158 354320
rect 237116 353394 237144 354311
rect 237104 353388 237156 353394
rect 237104 353330 237156 353336
rect 237012 353320 237064 353326
rect 237012 353262 237064 353268
rect 236932 350506 237144 350534
rect 237010 341728 237066 341737
rect 237010 341663 237066 341672
rect 236920 340332 236972 340338
rect 236920 340274 236972 340280
rect 236826 305552 236882 305561
rect 236826 305487 236882 305496
rect 236642 302288 236698 302297
rect 236642 302223 236698 302232
rect 236366 253328 236422 253337
rect 236366 253263 236422 253272
rect 236932 250073 236960 340274
rect 237024 251161 237052 341663
rect 237116 323105 237144 350506
rect 237102 323096 237158 323105
rect 237102 323031 237158 323040
rect 237208 268569 237236 365463
rect 237300 271833 237328 380695
rect 237944 369073 237972 390116
rect 238666 388512 238722 388521
rect 238666 388447 238722 388456
rect 238482 388376 238538 388385
rect 238482 388311 238538 388320
rect 237930 369064 237986 369073
rect 237930 368999 237986 369008
rect 238298 363760 238354 363769
rect 238298 363695 238354 363704
rect 238036 355570 238248 355586
rect 238036 355564 238260 355570
rect 238036 355558 238208 355564
rect 237748 355360 237800 355366
rect 237748 355302 237800 355308
rect 237760 327457 237788 355302
rect 237840 354000 237892 354006
rect 237840 353942 237892 353948
rect 237852 340241 237880 353942
rect 237932 350668 237984 350674
rect 237932 350610 237984 350616
rect 237838 340232 237894 340241
rect 237838 340167 237894 340176
rect 237746 327448 237802 327457
rect 237746 327383 237802 327392
rect 237746 326496 237802 326505
rect 237746 326431 237802 326440
rect 237760 296857 237788 326431
rect 237838 323640 237894 323649
rect 237838 323575 237894 323584
rect 237746 296848 237802 296857
rect 237746 296783 237802 296792
rect 237852 294681 237880 323575
rect 237944 321473 237972 350610
rect 238036 325281 238064 355558
rect 238208 355506 238260 355512
rect 238206 355464 238262 355473
rect 238206 355399 238262 355408
rect 238114 354920 238170 354929
rect 238114 354855 238170 354864
rect 238022 325272 238078 325281
rect 238022 325207 238078 325216
rect 238128 324193 238156 354855
rect 238114 324184 238170 324193
rect 238114 324119 238170 324128
rect 237930 321464 237986 321473
rect 237930 321399 237986 321408
rect 238220 317665 238248 355399
rect 238206 317656 238262 317665
rect 238206 317591 238262 317600
rect 238022 317384 238078 317393
rect 238022 317319 238078 317328
rect 238036 297945 238064 317319
rect 238312 314401 238340 363695
rect 238390 356008 238446 356017
rect 238390 355943 238392 355952
rect 238444 355943 238446 355952
rect 238392 355914 238444 355920
rect 238392 340264 238444 340270
rect 238392 340206 238444 340212
rect 238298 314392 238354 314401
rect 238298 314327 238354 314336
rect 238022 297936 238078 297945
rect 238022 297871 238078 297880
rect 237838 294672 237894 294681
rect 237838 294607 237894 294616
rect 238404 280537 238432 340206
rect 238496 308825 238524 388311
rect 238574 379128 238630 379137
rect 238574 379063 238630 379072
rect 238588 315489 238616 379063
rect 238574 315480 238630 315489
rect 238574 315415 238630 315424
rect 238574 313984 238630 313993
rect 238574 313919 238630 313928
rect 238482 308816 238538 308825
rect 238482 308751 238538 308760
rect 238390 280528 238446 280537
rect 238390 280463 238446 280472
rect 237286 271824 237342 271833
rect 237286 271759 237342 271768
rect 237194 268560 237250 268569
rect 237194 268495 237250 268504
rect 237010 251152 237066 251161
rect 237010 251087 237066 251096
rect 236918 250064 236974 250073
rect 236918 249999 236974 250008
rect 233882 241360 233938 241369
rect 233882 241295 233938 241304
rect 233896 202201 233924 241295
rect 237378 236056 237434 236065
rect 237378 235991 237434 236000
rect 237392 229094 237420 235991
rect 238206 229392 238262 229401
rect 238206 229327 238262 229336
rect 237300 229066 237420 229094
rect 233882 202192 233938 202201
rect 233882 202127 233938 202136
rect 233882 193488 233938 193497
rect 233882 193423 233938 193432
rect 233146 150104 233202 150113
rect 233146 150039 233202 150048
rect 233422 104408 233478 104417
rect 233422 104343 233478 104352
rect 228362 101552 228418 101561
rect 228362 101487 228418 101496
rect 229834 3904 229890 3913
rect 229834 3839 229890 3848
rect 229848 480 229876 3839
rect 233436 480 233464 104343
rect 233896 17513 233924 193423
rect 235906 172816 235962 172825
rect 235906 172751 235962 172760
rect 235722 156632 235778 156641
rect 235722 156567 235778 156576
rect 235354 153232 235410 153241
rect 235354 153167 235410 153176
rect 235262 136912 235318 136921
rect 235262 136847 235318 136856
rect 235276 118833 235304 136847
rect 235368 120465 235396 153167
rect 235736 140321 235764 156567
rect 235814 155952 235870 155961
rect 235814 155887 235870 155896
rect 235722 140312 235778 140321
rect 235722 140247 235778 140256
rect 235828 128354 235856 155887
rect 235644 128326 235856 128354
rect 235354 120456 235410 120465
rect 235354 120391 235410 120400
rect 235644 120306 235672 128326
rect 235920 120986 235948 172751
rect 237300 152153 237328 229066
rect 238114 228304 238170 228313
rect 238114 228239 238170 228248
rect 238022 227216 238078 227225
rect 238022 227151 238078 227160
rect 237470 217424 237526 217433
rect 237470 217359 237526 217368
rect 237378 216336 237434 216345
rect 237378 216271 237434 216280
rect 237392 215393 237420 216271
rect 237378 215384 237434 215393
rect 237378 215319 237434 215328
rect 237484 197985 237512 217359
rect 237470 197976 237526 197985
rect 237470 197911 237526 197920
rect 238036 192681 238064 227151
rect 238128 194041 238156 228239
rect 238220 196625 238248 229327
rect 238588 226409 238616 313919
rect 238680 289241 238708 388447
rect 239692 382265 239720 390116
rect 239956 384328 240008 384334
rect 239956 384270 240008 384276
rect 239678 382256 239734 382265
rect 239678 382191 239734 382200
rect 239312 378208 239364 378214
rect 239312 378150 239364 378156
rect 238852 375420 238904 375426
rect 238852 375362 238904 375368
rect 238864 373318 238892 375362
rect 238852 373312 238904 373318
rect 238852 373254 238904 373260
rect 239324 360194 239352 378150
rect 239494 361176 239550 361185
rect 239494 361111 239550 361120
rect 239140 360166 239352 360194
rect 239140 352730 239168 360166
rect 239402 355328 239458 355337
rect 239324 355286 239402 355314
rect 239324 353002 239352 355286
rect 239402 355263 239458 355272
rect 239402 354648 239458 354657
rect 239402 354583 239458 354592
rect 239416 353462 239444 354583
rect 239404 353456 239456 353462
rect 239404 353398 239456 353404
rect 239324 352974 239444 353002
rect 239140 352702 239352 352730
rect 239220 342984 239272 342990
rect 239220 342926 239272 342932
rect 239232 341578 239260 342926
rect 239140 341550 239260 341578
rect 239140 338638 239168 341550
rect 239218 341456 239274 341465
rect 239218 341391 239274 341400
rect 239232 339153 239260 341391
rect 239218 339144 239274 339153
rect 239218 339079 239274 339088
rect 239128 338632 239180 338638
rect 239128 338574 239180 338580
rect 239324 313993 239352 352702
rect 239416 322017 239444 352974
rect 239402 322008 239458 322017
rect 239402 321943 239458 321952
rect 239508 316577 239536 361111
rect 239678 354376 239734 354385
rect 239678 354311 239734 354320
rect 239588 351348 239640 351354
rect 239588 351290 239640 351296
rect 239494 316568 239550 316577
rect 239494 316503 239550 316512
rect 239310 313984 239366 313993
rect 239310 313919 239366 313928
rect 239600 304473 239628 351290
rect 239586 304464 239642 304473
rect 239586 304399 239642 304408
rect 239692 300121 239720 354311
rect 239864 351280 239916 351286
rect 239864 351222 239916 351228
rect 239770 339416 239826 339425
rect 239770 339351 239826 339360
rect 239784 338745 239812 339351
rect 239770 338736 239826 338745
rect 239770 338671 239826 338680
rect 239772 338632 239824 338638
rect 239772 338574 239824 338580
rect 239678 300112 239734 300121
rect 239678 300047 239734 300056
rect 238666 289232 238722 289241
rect 238666 289167 238722 289176
rect 239784 252249 239812 338574
rect 239770 252240 239826 252249
rect 239770 252175 239826 252184
rect 238574 226400 238630 226409
rect 238574 226335 238630 226344
rect 238298 226128 238354 226137
rect 238298 226063 238354 226072
rect 238206 196616 238262 196625
rect 238206 196551 238262 196560
rect 238114 194032 238170 194041
rect 238114 193967 238170 193976
rect 238022 192672 238078 192681
rect 238022 192607 238078 192616
rect 238206 187912 238262 187921
rect 238206 187847 238262 187856
rect 238022 185056 238078 185065
rect 238022 184991 238078 185000
rect 238036 173913 238064 184991
rect 238114 181520 238170 181529
rect 238114 181455 238170 181464
rect 238022 173904 238078 173913
rect 238022 173839 238078 173848
rect 237380 155916 237432 155922
rect 237380 155858 237432 155864
rect 237392 155417 237420 155858
rect 237378 155408 237434 155417
rect 237378 155343 237434 155352
rect 237380 154556 237432 154562
rect 237380 154498 237432 154504
rect 237392 154329 237420 154498
rect 237378 154320 237434 154329
rect 237378 154255 237434 154264
rect 237286 152144 237342 152153
rect 237286 152079 237342 152088
rect 238022 123584 238078 123593
rect 238022 123519 238078 123528
rect 235736 120958 235948 120986
rect 235736 120601 235764 120958
rect 235814 120864 235870 120873
rect 235814 120799 235870 120808
rect 235828 120698 235856 120799
rect 235906 120728 235962 120737
rect 235816 120692 235868 120698
rect 235906 120663 235962 120672
rect 235816 120634 235868 120640
rect 235920 120630 235948 120663
rect 235908 120624 235960 120630
rect 235722 120592 235778 120601
rect 235908 120566 235960 120572
rect 235722 120527 235778 120536
rect 235814 120320 235870 120329
rect 235644 120278 235814 120306
rect 235814 120255 235870 120264
rect 237286 120320 237342 120329
rect 237562 120320 237618 120329
rect 237342 120278 237562 120306
rect 237286 120255 237342 120264
rect 237562 120255 237618 120264
rect 235816 119604 235868 119610
rect 235816 119546 235868 119552
rect 235828 118969 235856 119546
rect 235908 119536 235960 119542
rect 235908 119478 235960 119484
rect 235920 119241 235948 119478
rect 235906 119232 235962 119241
rect 235906 119167 235962 119176
rect 235814 118960 235870 118969
rect 235814 118895 235870 118904
rect 235262 118824 235318 118833
rect 235262 118759 235318 118768
rect 234620 118652 234672 118658
rect 234620 118594 234672 118600
rect 234632 117337 234660 118594
rect 237564 118584 237616 118590
rect 237564 118526 237616 118532
rect 237380 118176 237432 118182
rect 237380 118118 237432 118124
rect 237392 117881 237420 118118
rect 237472 118108 237524 118114
rect 237472 118050 237524 118056
rect 237378 117872 237434 117881
rect 237378 117807 237434 117816
rect 237484 117745 237512 118050
rect 237470 117736 237526 117745
rect 237470 117671 237526 117680
rect 237576 117473 237604 118526
rect 238036 118250 238064 123519
rect 238024 118244 238076 118250
rect 238024 118186 238076 118192
rect 237562 117464 237618 117473
rect 237562 117399 237618 117408
rect 234618 117328 234674 117337
rect 234618 117263 234674 117272
rect 234620 115796 234672 115802
rect 234620 115738 234672 115744
rect 234632 115297 234660 115738
rect 234618 115288 234674 115297
rect 234618 115223 234674 115232
rect 233882 17504 233938 17513
rect 233882 17439 233938 17448
rect 237010 7712 237066 7721
rect 237010 7647 237066 7656
rect 237024 480 237052 7647
rect 238128 6361 238156 181455
rect 238220 118386 238248 187847
rect 238312 185745 238340 226063
rect 238574 216336 238630 216345
rect 238574 216271 238630 216280
rect 238482 187776 238538 187785
rect 238482 187711 238538 187720
rect 238392 186992 238444 186998
rect 238392 186934 238444 186940
rect 238298 185736 238354 185745
rect 238298 185671 238354 185680
rect 238404 156505 238432 186934
rect 238496 158681 238524 187711
rect 238482 158672 238538 158681
rect 238482 158607 238538 158616
rect 238390 156496 238446 156505
rect 238390 156431 238446 156440
rect 238482 139088 238538 139097
rect 238482 139023 238538 139032
rect 238390 138000 238446 138009
rect 238390 137935 238446 137944
rect 238404 122058 238432 137935
rect 238392 122052 238444 122058
rect 238392 121994 238444 122000
rect 238298 120048 238354 120057
rect 238298 119983 238354 119992
rect 238312 119678 238340 119983
rect 238300 119672 238352 119678
rect 238300 119614 238352 119620
rect 238208 118380 238260 118386
rect 238208 118322 238260 118328
rect 238496 118318 238524 139023
rect 238588 119746 238616 216271
rect 238666 215248 238722 215257
rect 238666 215183 238722 215192
rect 238680 187921 238708 215183
rect 238666 187912 238722 187921
rect 238666 187847 238722 187856
rect 238666 173904 238722 173913
rect 238666 173839 238722 173848
rect 238576 119740 238628 119746
rect 238576 119682 238628 119688
rect 238574 119504 238630 119513
rect 238574 119439 238576 119448
rect 238628 119439 238630 119448
rect 238576 119410 238628 119416
rect 238680 118697 238708 173839
rect 239876 147869 239904 351222
rect 239862 147860 239918 147869
rect 239862 147795 239918 147804
rect 239862 146772 239918 146781
rect 239968 146758 239996 384270
rect 240048 382220 240100 382226
rect 240048 382162 240100 382168
rect 240060 381177 240088 382162
rect 240046 381168 240102 381177
rect 240046 381103 240102 381112
rect 240048 354680 240100 354686
rect 240048 354622 240100 354628
rect 240060 353433 240088 354622
rect 240046 353424 240102 353433
rect 240046 353359 240102 353368
rect 240048 353252 240100 353258
rect 240048 353194 240100 353200
rect 240060 350538 240088 353194
rect 240048 350532 240100 350538
rect 240048 350474 240100 350480
rect 240048 342236 240100 342242
rect 240048 342178 240100 342184
rect 240060 341737 240088 342178
rect 240046 341728 240102 341737
rect 240046 341663 240102 341672
rect 241440 340218 241468 390116
rect 242990 359544 243046 359553
rect 242990 359479 243046 359488
rect 241440 340190 241560 340218
rect 241426 340096 241482 340105
rect 241532 340082 241560 340190
rect 241610 340096 241666 340105
rect 241532 340054 241610 340082
rect 241426 340031 241482 340040
rect 241610 340031 241666 340040
rect 242360 340066 242480 340082
rect 242360 340060 242492 340066
rect 242360 340054 242440 340060
rect 241440 339998 241468 340031
rect 241428 339992 241480 339998
rect 242360 339946 242388 340054
rect 242440 340002 242492 340008
rect 241428 339934 241480 339940
rect 242098 339918 242388 339946
rect 243004 339932 243032 359479
rect 243188 344457 243216 390116
rect 243542 347032 243598 347041
rect 243542 346967 243598 346976
rect 244094 347032 244150 347041
rect 244094 346967 244150 346976
rect 243556 346866 243584 346967
rect 243544 346860 243596 346866
rect 243544 346802 243596 346808
rect 243544 345024 243596 345030
rect 243544 344966 243596 344972
rect 243174 344448 243230 344457
rect 243174 344383 243230 344392
rect 243556 343777 243584 344966
rect 243542 343768 243598 343777
rect 243542 343703 243598 343712
rect 244108 339946 244136 346967
rect 244278 345808 244334 345817
rect 244278 345743 244334 345752
rect 244292 345574 244320 345743
rect 244280 345568 244332 345574
rect 244280 345510 244332 345516
rect 244830 345128 244886 345137
rect 244830 345063 244886 345072
rect 244278 343632 244334 343641
rect 244278 343567 244334 343576
rect 244292 342446 244320 343567
rect 244280 342440 244332 342446
rect 244280 342382 244332 342388
rect 243938 339918 244136 339946
rect 244844 339932 244872 345063
rect 244936 342961 244964 390116
rect 245750 357912 245806 357921
rect 245750 357847 245806 357856
rect 244922 342952 244978 342961
rect 244922 342887 244978 342896
rect 245764 339932 245792 357847
rect 246684 357649 246712 390116
rect 247590 359272 247646 359281
rect 247590 359207 247646 359216
rect 246762 358592 246818 358601
rect 246762 358527 246818 358536
rect 246670 357640 246726 357649
rect 246670 357575 246726 357584
rect 246776 339946 246804 358527
rect 246698 339918 246804 339946
rect 247604 339932 247632 359207
rect 248432 349194 248460 390116
rect 248510 360088 248566 360097
rect 248510 360023 248566 360032
rect 248340 349166 248460 349194
rect 248340 348537 248368 349166
rect 248326 348528 248382 348537
rect 248326 348463 248382 348472
rect 248524 339932 248552 360023
rect 249430 359952 249486 359961
rect 249430 359887 249486 359896
rect 249444 339932 249472 359887
rect 249706 349072 249762 349081
rect 249706 349007 249762 349016
rect 249720 348362 249748 349007
rect 249708 348356 249760 348362
rect 249708 348298 249760 348304
rect 250180 344321 250208 390116
rect 251928 360777 251956 390116
rect 251914 360768 251970 360777
rect 251914 360703 251970 360712
rect 252190 359816 252246 359825
rect 252190 359751 252246 359760
rect 251270 359000 251326 359009
rect 251270 358935 251326 358944
rect 251086 344720 251142 344729
rect 251086 344655 251142 344664
rect 251100 344350 251128 344655
rect 251088 344344 251140 344350
rect 250166 344312 250222 344321
rect 251088 344286 251140 344292
rect 250166 344247 250222 344256
rect 250352 343052 250404 343058
rect 250352 342994 250404 343000
rect 250364 339932 250392 342994
rect 250996 339992 251048 339998
rect 250996 339934 251048 339940
rect 250904 339924 250956 339930
rect 250904 339866 250956 339872
rect 250916 339425 250944 339866
rect 251008 339561 251036 339934
rect 251284 339932 251312 358935
rect 252204 339932 252232 359751
rect 252374 359680 252430 359689
rect 252374 359615 252430 359624
rect 252650 359680 252706 359689
rect 252650 359615 252706 359624
rect 252388 358834 252416 359615
rect 252466 359136 252522 359145
rect 252466 359071 252522 359080
rect 252480 358902 252508 359071
rect 252664 359009 252692 359615
rect 253204 359576 253256 359582
rect 253204 359518 253256 359524
rect 252650 359000 252706 359009
rect 252650 358935 252706 358944
rect 252468 358896 252520 358902
rect 252468 358838 252520 358844
rect 252376 358828 252428 358834
rect 252376 358770 252428 358776
rect 253112 346316 253164 346322
rect 253112 346258 253164 346264
rect 253124 345953 253152 346258
rect 253110 345944 253166 345953
rect 253110 345879 253166 345888
rect 253216 343058 253244 359518
rect 253676 345817 253704 390116
rect 254950 357368 255006 357377
rect 254950 357303 255006 357312
rect 254030 356552 254086 356561
rect 254030 356487 254086 356496
rect 253662 345808 253718 345817
rect 253662 345743 253718 345752
rect 253204 343052 253256 343058
rect 253204 342994 253256 343000
rect 253480 343052 253532 343058
rect 253480 342994 253532 343000
rect 253492 339946 253520 342994
rect 253138 339918 253520 339946
rect 254044 339932 254072 356487
rect 254584 349376 254636 349382
rect 254584 349318 254636 349324
rect 254596 344418 254624 349318
rect 254584 344412 254636 344418
rect 254584 344354 254636 344360
rect 254964 339932 254992 357303
rect 255318 344992 255374 345001
rect 255318 344927 255374 344936
rect 255332 344282 255360 344927
rect 255320 344276 255372 344282
rect 255320 344218 255372 344224
rect 255424 343233 255452 390116
rect 255870 357232 255926 357241
rect 255870 357167 255926 357176
rect 255410 343224 255466 343233
rect 255410 343159 255466 343168
rect 255884 339932 255912 357167
rect 256790 357096 256846 357105
rect 256790 357031 256846 357040
rect 256698 342000 256754 342009
rect 256698 341935 256754 341944
rect 256712 341698 256740 341935
rect 256700 341692 256752 341698
rect 256700 341634 256752 341640
rect 256804 339932 256832 357031
rect 257172 341873 257200 390116
rect 257710 356960 257766 356969
rect 257710 356895 257766 356904
rect 257158 341864 257214 341873
rect 257158 341799 257214 341808
rect 257724 339932 257752 356895
rect 258630 356824 258686 356833
rect 258630 356759 258686 356768
rect 258644 339932 258672 356759
rect 258920 348809 258948 390116
rect 260472 356856 260524 356862
rect 260472 356798 260524 356804
rect 259550 356688 259606 356697
rect 259550 356623 259606 356632
rect 258906 348800 258962 348809
rect 258906 348735 258962 348744
rect 259368 348628 259420 348634
rect 259368 348570 259420 348576
rect 259380 348401 259408 348570
rect 259366 348392 259422 348401
rect 259366 348327 259422 348336
rect 259564 339932 259592 356623
rect 259642 348800 259698 348809
rect 259642 348735 259698 348744
rect 259656 348401 259684 348735
rect 259642 348392 259698 348401
rect 259642 348327 259698 348336
rect 260484 339932 260512 356798
rect 260668 345953 260696 390116
rect 262416 387161 262444 390116
rect 262402 387152 262458 387161
rect 262402 387087 262458 387096
rect 263230 380624 263286 380633
rect 263230 380559 263286 380568
rect 262954 359816 263010 359825
rect 262692 359774 262954 359802
rect 262692 359689 262720 359774
rect 262954 359751 263010 359760
rect 262678 359680 262734 359689
rect 262678 359615 262734 359624
rect 261392 356788 261444 356794
rect 261392 356730 261444 356736
rect 260748 346384 260800 346390
rect 260748 346326 260800 346332
rect 260654 345944 260710 345953
rect 260654 345879 260710 345888
rect 260760 345137 260788 346326
rect 260746 345128 260802 345137
rect 260746 345063 260802 345072
rect 261404 339932 261432 356730
rect 262312 343120 262364 343126
rect 262312 343062 262364 343068
rect 262324 339932 262352 343062
rect 263244 339932 263272 380559
rect 264164 373425 264192 390116
rect 265912 386345 265940 390116
rect 265898 386336 265954 386345
rect 265898 386271 265954 386280
rect 265070 385928 265126 385937
rect 265070 385863 265126 385872
rect 264150 373416 264206 373425
rect 264150 373351 264206 373360
rect 264980 373312 265032 373318
rect 264980 373254 265032 373260
rect 264992 369170 265020 373254
rect 264980 369164 265032 369170
rect 264980 369106 265032 369112
rect 264150 365120 264206 365129
rect 264150 365055 264206 365064
rect 264164 339932 264192 365055
rect 265084 339932 265112 385863
rect 266360 382152 266412 382158
rect 266360 382094 266412 382100
rect 266910 382120 266966 382129
rect 266372 381041 266400 382094
rect 266910 382055 266966 382064
rect 266358 381032 266414 381041
rect 266358 380967 266414 380976
rect 265990 363896 266046 363905
rect 265990 363831 266046 363840
rect 266004 339932 266032 363831
rect 266360 346996 266412 347002
rect 266360 346938 266412 346944
rect 266372 346497 266400 346938
rect 266358 346488 266414 346497
rect 266358 346423 266414 346432
rect 266924 339932 266952 382055
rect 267660 347449 267688 390116
rect 268750 357776 268806 357785
rect 268750 357711 268806 357720
rect 267830 355736 267886 355745
rect 267830 355671 267886 355680
rect 267646 347440 267702 347449
rect 267646 347375 267702 347384
rect 267844 339932 267872 355671
rect 268382 340368 268438 340377
rect 268382 340303 268438 340312
rect 268396 339969 268424 340303
rect 268382 339960 268438 339969
rect 268764 339932 268792 357711
rect 269028 355836 269080 355842
rect 269028 355778 269080 355784
rect 269040 354929 269068 355778
rect 269026 354920 269082 354929
rect 269026 354855 269082 354864
rect 269408 341737 269436 390116
rect 269670 358320 269726 358329
rect 269670 358255 269726 358264
rect 269394 341728 269450 341737
rect 269394 341663 269450 341672
rect 269684 339932 269712 358255
rect 270590 358184 270646 358193
rect 270590 358119 270646 358128
rect 270408 341760 270460 341766
rect 270408 341702 270460 341708
rect 270420 341329 270448 341702
rect 270406 341320 270462 341329
rect 270406 341255 270462 341264
rect 270604 339932 270632 358119
rect 271156 344593 271184 390116
rect 272904 387705 272932 390116
rect 273904 390040 273956 390046
rect 273904 389982 273956 389988
rect 272890 387696 272946 387705
rect 272890 387631 272946 387640
rect 273916 382294 273944 389982
rect 273904 382288 273956 382294
rect 273904 382230 273956 382236
rect 271786 358728 271842 358737
rect 271786 358663 271788 358672
rect 271840 358663 271842 358672
rect 271788 358634 271840 358640
rect 272432 358624 272484 358630
rect 272432 358566 272484 358572
rect 271786 358456 271842 358465
rect 271786 358391 271842 358400
rect 271510 358048 271566 358057
rect 271510 357983 271566 357992
rect 271142 344584 271198 344593
rect 271142 344519 271198 344528
rect 271524 339932 271552 357983
rect 271800 357474 271828 358391
rect 271788 357468 271840 357474
rect 271788 357410 271840 357416
rect 271788 344412 271840 344418
rect 271788 344354 271840 344360
rect 271800 344185 271828 344354
rect 271786 344176 271842 344185
rect 271786 344111 271842 344120
rect 272444 339932 272472 358566
rect 273352 358556 273404 358562
rect 273352 358498 273404 358504
rect 273260 346928 273312 346934
rect 273260 346870 273312 346876
rect 273272 346322 273300 346870
rect 273260 346316 273312 346322
rect 273260 346258 273312 346264
rect 273364 339932 273392 358498
rect 274272 358488 274324 358494
rect 274272 358430 274324 358436
rect 274284 339932 274312 358430
rect 274652 346089 274680 390116
rect 274732 389972 274784 389978
rect 274732 389914 274784 389920
rect 274744 384402 274772 389914
rect 274732 384396 274784 384402
rect 274732 384338 274784 384344
rect 276020 373992 276072 373998
rect 276020 373934 276072 373940
rect 276032 372745 276060 373934
rect 276018 372736 276074 372745
rect 276018 372671 276074 372680
rect 276020 369164 276072 369170
rect 276020 369106 276072 369112
rect 276032 366722 276060 369106
rect 276020 366716 276072 366722
rect 276020 366658 276072 366664
rect 275192 358420 275244 358426
rect 275192 358362 275244 358368
rect 274638 346080 274694 346089
rect 274638 346015 274694 346024
rect 274638 345672 274694 345681
rect 274638 345607 274640 345616
rect 274692 345607 274694 345616
rect 274640 345578 274692 345584
rect 275204 339932 275232 358362
rect 276400 356017 276428 390116
rect 276664 382288 276716 382294
rect 276664 382230 276716 382236
rect 276676 371249 276704 382230
rect 277030 373688 277086 373697
rect 277030 373623 277086 373632
rect 276662 371240 276718 371249
rect 276662 371175 276718 371184
rect 276386 356008 276442 356017
rect 276386 355943 276442 355952
rect 276020 355904 276072 355910
rect 276020 355846 276072 355852
rect 276032 355065 276060 355846
rect 276018 355056 276074 355065
rect 276018 354991 276074 355000
rect 276112 343188 276164 343194
rect 276112 343130 276164 343136
rect 276020 342848 276072 342854
rect 276020 342790 276072 342796
rect 276032 340406 276060 342790
rect 276020 340400 276072 340406
rect 276020 340342 276072 340348
rect 275744 340060 275796 340066
rect 275744 340002 275796 340008
rect 268382 339895 268438 339904
rect 275756 339561 275784 340002
rect 276124 339932 276152 343130
rect 277044 339932 277072 373623
rect 277952 350940 278004 350946
rect 277952 350882 278004 350888
rect 277964 339932 277992 350882
rect 278044 348492 278096 348498
rect 278044 348434 278096 348440
rect 278056 340474 278084 348434
rect 278148 345014 278176 390116
rect 279606 387696 279662 387705
rect 279606 387631 279662 387640
rect 279422 387016 279478 387025
rect 279422 386951 279478 386960
rect 278964 345840 279016 345846
rect 278964 345782 279016 345788
rect 278976 345014 279004 345782
rect 279436 345014 279464 386951
rect 279620 364334 279648 387631
rect 279620 364306 279740 364334
rect 279712 345014 279740 364306
rect 279896 345014 279924 390116
rect 280066 387152 280122 387161
rect 280066 387087 280122 387096
rect 278148 344986 278452 345014
rect 278976 344986 279096 345014
rect 279436 344986 279648 345014
rect 279712 344986 279832 345014
rect 279896 344986 280016 345014
rect 278044 340468 278096 340474
rect 278044 340410 278096 340416
rect 250994 339552 251050 339561
rect 275742 339552 275798 339561
rect 250994 339487 251050 339496
rect 274640 339516 274692 339522
rect 275742 339487 275798 339496
rect 274640 339458 274692 339464
rect 274652 339425 274680 339458
rect 278424 339425 278452 344986
rect 279068 340134 279096 344986
rect 279332 344344 279384 344350
rect 279332 344286 279384 344292
rect 279056 340128 279108 340134
rect 279056 340070 279108 340076
rect 279344 339454 279372 344286
rect 279514 343768 279570 343777
rect 279514 343703 279570 343712
rect 279424 342712 279476 342718
rect 279424 342654 279476 342660
rect 279436 339454 279464 342654
rect 279528 339454 279556 343703
rect 279620 339454 279648 344986
rect 279804 339998 279832 344986
rect 279792 339992 279844 339998
rect 279792 339934 279844 339940
rect 279988 339946 280016 344986
rect 280080 340066 280108 387087
rect 281644 384849 281672 390116
rect 283392 386889 283420 390116
rect 283378 386880 283434 386889
rect 283378 386815 283434 386824
rect 282182 385656 282238 385665
rect 282182 385591 282238 385600
rect 282092 385008 282144 385014
rect 282092 384950 282144 384956
rect 281630 384840 281686 384849
rect 281630 384775 281686 384784
rect 282104 383761 282132 384950
rect 282090 383752 282146 383761
rect 282090 383687 282146 383696
rect 280894 373416 280950 373425
rect 280894 373351 280950 373360
rect 280802 369064 280858 369073
rect 280802 368999 280858 369008
rect 280434 351384 280490 351393
rect 280434 351319 280490 351328
rect 280252 351144 280304 351150
rect 280252 351086 280304 351092
rect 280160 345908 280212 345914
rect 280160 345850 280212 345856
rect 280172 345681 280200 345850
rect 280158 345672 280214 345681
rect 280158 345607 280214 345616
rect 280068 340060 280120 340066
rect 280068 340002 280120 340008
rect 279988 339918 280200 339946
rect 280066 339824 280122 339833
rect 280066 339759 280122 339768
rect 279332 339448 279384 339454
rect 250902 339416 250958 339425
rect 250902 339351 250958 339360
rect 274638 339416 274694 339425
rect 274638 339351 274694 339360
rect 278410 339416 278466 339425
rect 279332 339390 279384 339396
rect 279424 339448 279476 339454
rect 279424 339390 279476 339396
rect 279516 339448 279568 339454
rect 279516 339390 279568 339396
rect 279608 339448 279660 339454
rect 279976 339448 280028 339454
rect 279608 339390 279660 339396
rect 279974 339416 279976 339425
rect 280028 339416 280030 339425
rect 278410 339351 278466 339360
rect 279974 339351 280030 339360
rect 280080 339266 280108 339759
rect 280172 339425 280200 339918
rect 280158 339416 280214 339425
rect 280158 339351 280214 339360
rect 280080 339238 280200 339266
rect 280066 339144 280122 339153
rect 280066 339079 280122 339088
rect 280080 338774 280108 339079
rect 280172 338978 280200 339238
rect 280160 338972 280212 338978
rect 280160 338914 280212 338920
rect 280068 338768 280120 338774
rect 280068 338710 280120 338716
rect 280066 338464 280122 338473
rect 280122 338422 280200 338450
rect 280066 338399 280122 338408
rect 280066 338328 280122 338337
rect 280172 338298 280200 338422
rect 280066 338263 280122 338272
rect 280160 338292 280212 338298
rect 280080 338230 280108 338263
rect 280160 338234 280212 338240
rect 280068 338224 280120 338230
rect 280068 338166 280120 338172
rect 280066 338056 280122 338065
rect 280066 337991 280122 338000
rect 280080 336705 280108 337991
rect 280158 337920 280214 337929
rect 280158 337855 280214 337864
rect 280066 336696 280122 336705
rect 280066 336631 280122 336640
rect 280172 336297 280200 337855
rect 280158 336288 280214 336297
rect 280158 336223 280214 336232
rect 280160 336184 280212 336190
rect 280160 336126 280212 336132
rect 280172 268569 280200 336126
rect 280264 303929 280292 351086
rect 280344 351008 280396 351014
rect 280344 350950 280396 350956
rect 280356 304473 280384 350950
rect 280448 305561 280476 351319
rect 280528 346792 280580 346798
rect 280528 346734 280580 346740
rect 280434 305552 280490 305561
rect 280434 305487 280490 305496
rect 280342 304464 280398 304473
rect 280342 304399 280398 304408
rect 280250 303920 280306 303929
rect 280250 303855 280306 303864
rect 280540 302841 280568 346734
rect 280712 343256 280764 343262
rect 280712 343198 280764 343204
rect 280620 341624 280672 341630
rect 280620 341566 280672 341572
rect 280632 307193 280660 341566
rect 280724 308825 280752 343198
rect 280710 308816 280766 308825
rect 280710 308751 280766 308760
rect 280618 307184 280674 307193
rect 280618 307119 280674 307128
rect 280526 302832 280582 302841
rect 280526 302767 280582 302776
rect 280816 301481 280844 368999
rect 280908 317801 280936 373351
rect 280986 357640 281042 357649
rect 280986 357575 281042 357584
rect 280894 317792 280950 317801
rect 280894 317727 280950 317736
rect 281000 306921 281028 357575
rect 282092 353184 282144 353190
rect 282092 353126 282144 353132
rect 282000 351416 282052 351422
rect 282000 351358 282052 351364
rect 281078 344040 281134 344049
rect 281078 343975 281134 343984
rect 281092 336190 281120 343975
rect 281356 340128 281408 340134
rect 281356 340070 281408 340076
rect 281172 340060 281224 340066
rect 281172 340002 281224 340008
rect 281080 336184 281132 336190
rect 281080 336126 281132 336132
rect 281184 336025 281212 340002
rect 281264 339992 281316 339998
rect 281264 339934 281316 339940
rect 281276 338745 281304 339934
rect 281262 338736 281318 338745
rect 281262 338671 281318 338680
rect 281368 336161 281396 340070
rect 281906 338872 281962 338881
rect 281906 338807 281962 338816
rect 281920 338473 281948 338807
rect 281906 338464 281962 338473
rect 281906 338399 281962 338408
rect 281354 336152 281410 336161
rect 281354 336087 281410 336096
rect 281170 336016 281226 336025
rect 281170 335951 281226 335960
rect 281816 307760 281868 307766
rect 281814 307728 281816 307737
rect 281868 307728 281870 307737
rect 281814 307663 281870 307672
rect 280986 306912 281042 306921
rect 280986 306847 281042 306856
rect 280802 301472 280858 301481
rect 280802 301407 280858 301416
rect 281906 298480 281962 298489
rect 281906 298415 281962 298424
rect 281920 298178 281948 298415
rect 281908 298172 281960 298178
rect 281908 298114 281960 298120
rect 281814 293040 281870 293049
rect 281814 292975 281870 292984
rect 281828 292602 281856 292975
rect 281816 292596 281868 292602
rect 281816 292538 281868 292544
rect 281906 292496 281962 292505
rect 281906 292431 281962 292440
rect 281920 291242 281948 292431
rect 281908 291236 281960 291242
rect 281908 291178 281960 291184
rect 281906 290864 281962 290873
rect 281906 290799 281962 290808
rect 281920 289882 281948 290799
rect 281908 289876 281960 289882
rect 281908 289818 281960 289824
rect 281906 289776 281962 289785
rect 281906 289711 281962 289720
rect 281920 288454 281948 289711
rect 281908 288448 281960 288454
rect 281908 288390 281960 288396
rect 282012 287065 282040 351358
rect 281998 287056 282054 287065
rect 281998 286991 282054 287000
rect 282104 284889 282132 353126
rect 282090 284880 282146 284889
rect 282090 284815 282146 284824
rect 282196 281625 282224 385591
rect 282552 378888 282604 378894
rect 282552 378830 282604 378836
rect 282276 378820 282328 378826
rect 282276 378762 282328 378768
rect 282288 285433 282316 378762
rect 282460 376100 282512 376106
rect 282460 376042 282512 376048
rect 282366 371920 282422 371929
rect 282366 371855 282422 371864
rect 282274 285424 282330 285433
rect 282274 285359 282330 285368
rect 282182 281616 282238 281625
rect 282182 281551 282238 281560
rect 282380 279993 282408 371855
rect 282472 283801 282500 376042
rect 282564 286521 282592 378830
rect 284942 372328 284998 372337
rect 284942 372263 284998 372272
rect 282642 362400 282698 362409
rect 282642 362335 282698 362344
rect 282550 286512 282606 286521
rect 282550 286447 282606 286456
rect 282458 283792 282514 283801
rect 282458 283727 282514 283736
rect 282366 279984 282422 279993
rect 282366 279919 282422 279928
rect 282656 277817 282684 362335
rect 282920 358692 282972 358698
rect 282920 358634 282972 358640
rect 282932 357513 282960 358634
rect 282918 357504 282974 357513
rect 282918 357439 282974 357448
rect 284300 355972 284352 355978
rect 284300 355914 284352 355920
rect 284312 355065 284340 355914
rect 284298 355056 284354 355065
rect 284298 354991 284354 355000
rect 283102 351928 283158 351937
rect 283102 351863 283158 351872
rect 282826 351112 282882 351121
rect 282826 351047 282882 351056
rect 283012 351076 283064 351082
rect 282736 350328 282788 350334
rect 282736 350270 282788 350276
rect 282748 278905 282776 350270
rect 282840 282713 282868 351047
rect 283012 351018 283064 351024
rect 282918 349072 282974 349081
rect 282918 349007 282974 349016
rect 282932 348566 282960 349007
rect 282920 348560 282972 348566
rect 282920 348502 282972 348508
rect 282920 342780 282972 342786
rect 282920 342722 282972 342728
rect 282932 308281 282960 342722
rect 282918 308272 282974 308281
rect 282918 308207 282974 308216
rect 283024 302297 283052 351018
rect 283116 305017 283144 351863
rect 284758 349480 284814 349489
rect 284758 349415 284814 349424
rect 283380 349240 283432 349246
rect 283380 349182 283432 349188
rect 283286 348664 283342 348673
rect 283286 348599 283342 348608
rect 283196 346860 283248 346866
rect 283196 346802 283248 346808
rect 283208 306649 283236 346802
rect 283194 306640 283250 306649
rect 283194 306575 283250 306584
rect 283102 305008 283158 305017
rect 283102 304943 283158 304952
rect 283010 302288 283066 302297
rect 283010 302223 283066 302232
rect 283010 293584 283066 293593
rect 283010 293519 283066 293528
rect 282826 282704 282882 282713
rect 282826 282639 282882 282648
rect 282734 278896 282790 278905
rect 282734 278831 282790 278840
rect 282642 277808 282698 277817
rect 282642 277743 282698 277752
rect 282090 269104 282146 269113
rect 282090 269039 282092 269048
rect 282144 269039 282146 269048
rect 282092 269010 282144 269016
rect 282828 269000 282880 269006
rect 282828 268942 282880 268948
rect 280158 268560 280214 268569
rect 280158 268495 280214 268504
rect 282840 268025 282868 268942
rect 282826 268016 282882 268025
rect 282826 267951 282882 267960
rect 282828 266348 282880 266354
rect 282828 266290 282880 266296
rect 282840 265305 282868 266290
rect 282826 265296 282882 265305
rect 282826 265231 282882 265240
rect 282828 264920 282880 264926
rect 282828 264862 282880 264868
rect 282840 264217 282868 264862
rect 282826 264208 282882 264217
rect 282826 264143 282882 264152
rect 282736 263560 282788 263566
rect 282736 263502 282788 263508
rect 282748 262585 282776 263502
rect 282828 263492 282880 263498
rect 282828 263434 282880 263440
rect 282840 263129 282868 263434
rect 282826 263120 282882 263129
rect 282826 263055 282882 263064
rect 282734 262576 282790 262585
rect 282734 262511 282790 262520
rect 282828 262200 282880 262206
rect 282828 262142 282880 262148
rect 282840 262041 282868 262142
rect 282826 262032 282882 262041
rect 282826 261967 282882 261976
rect 282828 260840 282880 260846
rect 282828 260782 282880 260788
rect 282840 259865 282868 260782
rect 282826 259856 282882 259865
rect 282826 259791 282882 259800
rect 282828 259412 282880 259418
rect 282828 259354 282880 259360
rect 282644 259344 282696 259350
rect 282840 259321 282868 259354
rect 282644 259286 282696 259292
rect 282826 259312 282882 259321
rect 282656 258777 282684 259286
rect 282736 259276 282788 259282
rect 282826 259247 282882 259256
rect 282736 259218 282788 259224
rect 282642 258768 282698 258777
rect 282642 258703 282698 258712
rect 282748 258233 282776 259218
rect 282734 258224 282790 258233
rect 282734 258159 282790 258168
rect 282736 258052 282788 258058
rect 282736 257994 282788 258000
rect 282748 257145 282776 257994
rect 282828 257984 282880 257990
rect 282828 257926 282880 257932
rect 282840 257689 282868 257926
rect 282826 257680 282882 257689
rect 282826 257615 282882 257624
rect 282734 257136 282790 257145
rect 282734 257071 282790 257080
rect 282644 256692 282696 256698
rect 282644 256634 282696 256640
rect 282656 256057 282684 256634
rect 282828 256624 282880 256630
rect 282826 256592 282828 256601
rect 282880 256592 282882 256601
rect 282736 256556 282788 256562
rect 282826 256527 282882 256536
rect 282736 256498 282788 256504
rect 282642 256048 282698 256057
rect 282642 255983 282698 255992
rect 282748 255513 282776 256498
rect 282734 255504 282790 255513
rect 282734 255439 282790 255448
rect 282828 255196 282880 255202
rect 282828 255138 282880 255144
rect 282840 254425 282868 255138
rect 282826 254416 282882 254425
rect 282826 254351 282882 254360
rect 282644 253904 282696 253910
rect 282644 253846 282696 253852
rect 282826 253872 282882 253881
rect 282656 253337 282684 253846
rect 282736 253836 282788 253842
rect 282826 253807 282882 253816
rect 282736 253778 282788 253784
rect 282642 253328 282698 253337
rect 282642 253263 282698 253272
rect 282748 252793 282776 253778
rect 282840 253774 282868 253807
rect 282828 253768 282880 253774
rect 282828 253710 282880 253716
rect 282734 252784 282790 252793
rect 282734 252719 282790 252728
rect 282736 252544 282788 252550
rect 282736 252486 282788 252492
rect 282748 251705 282776 252486
rect 282828 252476 282880 252482
rect 282828 252418 282880 252424
rect 282840 252249 282868 252418
rect 282826 252240 282882 252249
rect 282826 252175 282882 252184
rect 282734 251696 282790 251705
rect 282734 251631 282790 251640
rect 282828 251184 282880 251190
rect 282826 251152 282828 251161
rect 282880 251152 282882 251161
rect 282736 251116 282788 251122
rect 282826 251087 282882 251096
rect 282736 251058 282788 251064
rect 282552 251048 282604 251054
rect 282552 250990 282604 250996
rect 282564 250073 282592 250990
rect 282748 250617 282776 251058
rect 282734 250608 282790 250617
rect 282734 250543 282790 250552
rect 282550 250064 282606 250073
rect 282550 249999 282606 250008
rect 282828 249756 282880 249762
rect 282828 249698 282880 249704
rect 282736 249688 282788 249694
rect 282736 249630 282788 249636
rect 282748 248441 282776 249630
rect 282840 248985 282868 249698
rect 282826 248976 282882 248985
rect 282826 248911 282882 248920
rect 282734 248432 282790 248441
rect 282734 248367 282790 248376
rect 282644 248124 282696 248130
rect 282644 248066 282696 248072
rect 282656 247897 282684 248066
rect 282642 247888 282698 247897
rect 282642 247823 282698 247832
rect 282828 247036 282880 247042
rect 282828 246978 282880 246984
rect 282840 246809 282868 246978
rect 282826 246800 282882 246809
rect 282826 246735 282882 246744
rect 282828 238740 282880 238746
rect 282828 238682 282880 238688
rect 282840 237561 282868 238682
rect 282826 237552 282882 237561
rect 282826 237487 282882 237496
rect 281540 235952 281592 235958
rect 281538 235920 281540 235929
rect 281592 235920 281594 235929
rect 281538 235855 281594 235864
rect 280250 229392 280306 229401
rect 280250 229327 280306 229336
rect 280158 223408 280214 223417
rect 280158 223343 280214 223352
rect 280066 192944 280122 192953
rect 280066 192879 280122 192888
rect 239918 146730 239996 146758
rect 239862 146707 239918 146716
rect 280080 135153 280108 192879
rect 280066 135144 280122 135153
rect 280066 135079 280122 135088
rect 280066 134736 280122 134745
rect 280066 134671 280122 134680
rect 239956 122052 240008 122058
rect 239956 121994 240008 122000
rect 238850 119368 238906 119377
rect 238850 119303 238906 119312
rect 238864 118833 238892 119303
rect 238850 118824 238906 118833
rect 238850 118759 238906 118768
rect 238666 118688 238722 118697
rect 238666 118623 238722 118632
rect 239968 118454 239996 121994
rect 279976 120556 280028 120562
rect 279976 120498 280028 120504
rect 279988 120329 280016 120498
rect 279974 120320 280030 120329
rect 279974 120255 280030 120264
rect 279698 120184 279754 120193
rect 279698 120119 279754 120128
rect 240902 120006 241008 120034
rect 242098 120006 242204 120034
rect 243294 120006 243400 120034
rect 239956 118448 240008 118454
rect 239956 118390 240008 118396
rect 238484 118312 238536 118318
rect 238484 118254 238536 118260
rect 240506 116240 240562 116249
rect 240506 116175 240562 116184
rect 238114 6352 238170 6361
rect 238114 6287 238170 6296
rect 240520 480 240548 116175
rect 240980 103514 241008 120006
rect 241428 116952 241480 116958
rect 241426 116920 241428 116929
rect 241480 116920 241482 116929
rect 241426 116855 241482 116864
rect 242176 103514 242204 120006
rect 243372 107001 243400 120006
rect 244292 120006 244490 120034
rect 245686 120006 245792 120034
rect 244292 117774 244320 120006
rect 245764 118658 245792 120006
rect 246592 120006 246882 120034
rect 247696 120006 248078 120034
rect 248984 120006 249274 120034
rect 250088 120006 250470 120034
rect 251376 120006 251666 120034
rect 252862 120006 252968 120034
rect 254058 120006 254164 120034
rect 255254 120006 255360 120034
rect 256450 120006 256556 120034
rect 257646 120006 257752 120034
rect 258842 120006 258948 120034
rect 260038 120006 260144 120034
rect 261234 120006 261340 120034
rect 262430 120006 262536 120034
rect 263626 120006 263732 120034
rect 264822 120006 264928 120034
rect 266018 120006 266124 120034
rect 267214 120006 267320 120034
rect 268410 120006 268516 120034
rect 269606 120006 269712 120034
rect 270802 120006 270908 120034
rect 271998 120006 272104 120034
rect 245752 118652 245804 118658
rect 245752 118594 245804 118600
rect 246592 118590 246620 120006
rect 247040 118652 247092 118658
rect 247040 118594 247092 118600
rect 246580 118584 246632 118590
rect 246580 118526 246632 118532
rect 244280 117768 244332 117774
rect 244280 117710 244332 117716
rect 247052 117609 247080 118594
rect 247696 118114 247724 120006
rect 247774 118280 247830 118289
rect 247774 118215 247830 118224
rect 247684 118108 247736 118114
rect 247684 118050 247736 118056
rect 247038 117600 247094 117609
rect 247038 117535 247094 117544
rect 243358 106992 243414 107001
rect 243358 106927 243414 106936
rect 247788 103514 247816 118215
rect 248984 118182 249012 120006
rect 250088 118658 250116 120006
rect 250076 118652 250128 118658
rect 250076 118594 250128 118600
rect 248972 118176 249024 118182
rect 248972 118118 249024 118124
rect 251376 118017 251404 120006
rect 251362 118008 251418 118017
rect 251362 117943 251418 117952
rect 252468 114504 252520 114510
rect 252468 114446 252520 114452
rect 251178 113656 251234 113665
rect 251178 113591 251234 113600
rect 240888 103486 241008 103514
rect 242084 103486 242204 103514
rect 247696 103486 247816 103514
rect 240888 100065 240916 103486
rect 240874 100056 240930 100065
rect 240874 99991 240930 100000
rect 242084 6225 242112 103486
rect 242070 6216 242126 6225
rect 242070 6151 242126 6160
rect 247696 3913 247724 103486
rect 247682 3904 247738 3913
rect 247682 3839 247738 3848
rect 247590 3768 247646 3777
rect 247590 3703 247646 3712
rect 244094 3632 244150 3641
rect 244094 3567 244150 3576
rect 244108 480 244136 3567
rect 247604 480 247632 3703
rect 251192 480 251220 113591
rect 252480 113257 252508 114446
rect 252466 113248 252522 113257
rect 252466 113183 252522 113192
rect 252940 103514 252968 120006
rect 254136 103514 254164 120006
rect 255332 119898 255360 120006
rect 252848 103486 252968 103514
rect 254044 103486 254164 103514
rect 255240 119870 255360 119898
rect 252848 22953 252876 103486
rect 254044 36689 254072 103486
rect 254030 36680 254086 36689
rect 254030 36615 254086 36624
rect 255240 35329 255268 119870
rect 256528 103514 256556 120006
rect 257724 103514 257752 120006
rect 258920 103514 258948 120006
rect 260116 103514 260144 120006
rect 261312 103514 261340 120006
rect 261758 117736 261814 117745
rect 261758 117671 261814 117680
rect 256436 103486 256556 103514
rect 257632 103486 257752 103514
rect 258828 103486 258948 103514
rect 260024 103486 260144 103514
rect 261220 103486 261340 103514
rect 255226 35320 255282 35329
rect 255226 35255 255282 35264
rect 256436 24313 256464 103486
rect 257632 33969 257660 103486
rect 257618 33960 257674 33969
rect 257618 33895 257674 33904
rect 258828 25673 258856 103486
rect 260024 27033 260052 103486
rect 261220 31113 261248 103486
rect 261206 31104 261262 31113
rect 261206 31039 261262 31048
rect 260010 27024 260066 27033
rect 260010 26959 260066 26968
rect 258814 25664 258870 25673
rect 258814 25599 258870 25608
rect 256422 24304 256478 24313
rect 256422 24239 256478 24248
rect 252834 22944 252890 22953
rect 252834 22879 252890 22888
rect 258262 4040 258318 4049
rect 258262 3975 258318 3984
rect 254674 3904 254730 3913
rect 254674 3839 254730 3848
rect 254688 480 254716 3839
rect 258276 480 258304 3975
rect 261772 480 261800 117671
rect 262508 103514 262536 120006
rect 263704 103514 263732 120006
rect 264900 103514 264928 120006
rect 264980 118176 265032 118182
rect 264980 118118 265032 118124
rect 264992 117473 265020 118118
rect 265346 118008 265402 118017
rect 265346 117943 265402 117952
rect 264978 117464 265034 117473
rect 264978 117399 265034 117408
rect 262416 103486 262536 103514
rect 263612 103486 263732 103514
rect 264808 103486 264928 103514
rect 262416 28393 262444 103486
rect 262402 28384 262458 28393
rect 262402 28319 262458 28328
rect 263612 6497 263640 103486
rect 264808 29889 264836 103486
rect 264794 29880 264850 29889
rect 264794 29815 264850 29824
rect 263598 6488 263654 6497
rect 263598 6423 263654 6432
rect 265360 480 265388 117943
rect 266096 103514 266124 120006
rect 267292 103514 267320 120006
rect 268488 103514 268516 120006
rect 269684 103514 269712 120006
rect 270880 104281 270908 120006
rect 271786 118416 271842 118425
rect 271786 118351 271842 118360
rect 271800 118114 271828 118351
rect 271788 118108 271840 118114
rect 271788 118050 271840 118056
rect 271142 117328 271198 117337
rect 271142 117263 271198 117272
rect 270866 104272 270922 104281
rect 270866 104207 270922 104216
rect 266004 103486 266124 103514
rect 267200 103486 267320 103514
rect 268396 103486 268516 103514
rect 269592 103486 269712 103514
rect 266004 98977 266032 103486
rect 265990 98968 266046 98977
rect 265990 98903 266046 98912
rect 267200 95849 267228 103486
rect 268396 102921 268424 103486
rect 268382 102912 268438 102921
rect 268382 102847 268438 102856
rect 269592 97345 269620 103486
rect 269578 97336 269634 97345
rect 269578 97271 269634 97280
rect 267186 95840 267242 95849
rect 267186 95775 267242 95784
rect 271156 89185 271184 117263
rect 272076 105641 272104 120006
rect 272904 120006 273194 120034
rect 274390 120006 274496 120034
rect 275586 120006 275692 120034
rect 272904 117337 272932 120006
rect 272890 117328 272946 117337
rect 272890 117263 272946 117272
rect 273902 117328 273958 117337
rect 273902 117263 273958 117272
rect 272062 105632 272118 105641
rect 272062 105567 272118 105576
rect 273916 93129 273944 117263
rect 274468 103514 274496 120006
rect 275664 103514 275692 120006
rect 276400 120006 276782 120034
rect 277688 120006 277978 120034
rect 279174 120006 279464 120034
rect 276400 117337 276428 120006
rect 277688 118153 277716 120006
rect 279436 118153 279464 120006
rect 277674 118144 277730 118153
rect 277674 118079 277730 118088
rect 279422 118144 279478 118153
rect 279422 118079 279478 118088
rect 276386 117328 276442 117337
rect 276386 117263 276442 117272
rect 279712 103514 279740 120119
rect 274376 103486 274496 103514
rect 275572 103486 275692 103514
rect 279436 103486 279740 103514
rect 273902 93120 273958 93129
rect 273902 93055 273958 93064
rect 274376 90545 274404 103486
rect 275572 91769 275600 103486
rect 275558 91760 275614 91769
rect 275558 91695 275614 91704
rect 274362 90536 274418 90545
rect 274362 90471 274418 90480
rect 271142 89176 271198 89185
rect 271142 89111 271198 89120
rect 275282 86048 275338 86057
rect 275282 85983 275338 85992
rect 271142 85912 271198 85921
rect 271142 85847 271198 85856
rect 267002 54496 267058 54505
rect 267002 54431 267058 54440
rect 267016 6225 267044 54431
rect 268842 49328 268898 49337
rect 268842 49263 268898 49272
rect 267002 6216 267058 6225
rect 267002 6151 267058 6160
rect 268856 480 268884 49263
rect 271156 3641 271184 85847
rect 275296 16574 275324 85983
rect 278042 69456 278098 69465
rect 278042 69391 278098 69400
rect 275296 16546 275968 16574
rect 271788 4140 271840 4146
rect 271788 4082 271840 4088
rect 271142 3632 271198 3641
rect 271142 3567 271198 3576
rect 270590 3496 270646 3505
rect 271050 3496 271106 3505
rect 270646 3454 271050 3482
rect 270590 3431 270646 3440
rect 271050 3431 271106 3440
rect 271800 2825 271828 4082
rect 272430 3632 272486 3641
rect 272430 3567 272486 3576
rect 271786 2816 271842 2825
rect 271786 2751 271842 2760
rect 272444 480 272472 3567
rect 275940 3074 275968 16546
rect 278056 5681 278084 69391
rect 278042 5672 278098 5681
rect 278042 5607 278098 5616
rect 279436 3369 279464 103486
rect 279514 4856 279570 4865
rect 279514 4791 279570 4800
rect 279422 3360 279478 3369
rect 279422 3295 279478 3304
rect 275940 3046 276060 3074
rect 276032 480 276060 3046
rect 279528 480 279556 4791
rect 280080 3233 280108 134671
rect 280172 111489 280200 223343
rect 280264 117745 280292 229327
rect 282550 228848 282606 228857
rect 282550 228783 282606 228792
rect 281538 228304 281594 228313
rect 281538 228239 281594 228248
rect 280342 226128 280398 226137
rect 280342 226063 280398 226072
rect 280250 117736 280306 117745
rect 280250 117671 280306 117680
rect 280356 116249 280384 226063
rect 280526 222320 280582 222329
rect 280526 222255 280582 222264
rect 280434 220688 280490 220697
rect 280434 220623 280490 220632
rect 280342 116240 280398 116249
rect 280342 116175 280398 116184
rect 280448 112713 280476 220623
rect 280540 115025 280568 222255
rect 280618 221776 280674 221785
rect 280618 221711 280674 221720
rect 280632 116385 280660 221711
rect 280894 218512 280950 218521
rect 280894 218447 280950 218456
rect 280710 216336 280766 216345
rect 280710 216271 280766 216280
rect 280618 116376 280674 116385
rect 280618 116311 280674 116320
rect 280526 115016 280582 115025
rect 280526 114951 280582 114960
rect 280724 114481 280752 216271
rect 280802 214568 280858 214577
rect 280802 214503 280858 214512
rect 280710 114472 280766 114481
rect 280710 114407 280766 114416
rect 280434 112704 280490 112713
rect 280434 112639 280490 112648
rect 280158 111480 280214 111489
rect 280158 111415 280214 111424
rect 280816 3913 280844 214503
rect 280908 116793 280936 218447
rect 281552 214577 281580 228239
rect 281630 227216 281686 227225
rect 281630 227151 281686 227160
rect 281538 214568 281594 214577
rect 281538 214503 281594 214512
rect 281644 209774 281672 227151
rect 281998 226672 282054 226681
rect 281998 226607 282054 226616
rect 281814 219056 281870 219065
rect 281814 218991 281870 219000
rect 281722 217968 281778 217977
rect 281722 217903 281778 217912
rect 281552 209746 281672 209774
rect 281552 204218 281580 209746
rect 281000 204190 281580 204218
rect 280894 116784 280950 116793
rect 280894 116719 280950 116728
rect 280802 3904 280858 3913
rect 280802 3839 280858 3848
rect 281000 3777 281028 204190
rect 281630 203280 281686 203289
rect 281630 203215 281686 203224
rect 281644 87553 281672 203215
rect 281736 101697 281764 217903
rect 281828 109993 281856 218991
rect 281906 217424 281962 217433
rect 281906 217359 281962 217368
rect 281920 111353 281948 217359
rect 282012 120193 282040 226607
rect 282090 224496 282146 224505
rect 282090 224431 282146 224440
rect 281998 120184 282054 120193
rect 281998 120119 282054 120128
rect 282104 118289 282132 224431
rect 282274 216880 282330 216889
rect 282274 216815 282330 216824
rect 282182 215248 282238 215257
rect 282182 215183 282238 215192
rect 282090 118280 282146 118289
rect 282090 118215 282146 118224
rect 282196 112849 282224 215183
rect 282288 115161 282316 216815
rect 282366 198384 282422 198393
rect 282366 198319 282422 198328
rect 282274 115152 282330 115161
rect 282274 115087 282330 115096
rect 282182 112840 282238 112849
rect 282182 112775 282238 112784
rect 281906 111344 281962 111353
rect 281906 111279 281962 111288
rect 281814 109984 281870 109993
rect 281814 109919 281870 109928
rect 281722 101688 281778 101697
rect 281722 101623 281778 101632
rect 282380 100201 282408 198319
rect 282564 197441 282592 228783
rect 282734 215792 282790 215801
rect 282734 215727 282790 215736
rect 282550 197432 282606 197441
rect 282550 197367 282606 197376
rect 282460 168360 282512 168366
rect 282460 168302 282512 168308
rect 282472 167385 282500 168302
rect 282642 167920 282698 167929
rect 282642 167855 282698 167864
rect 282458 167376 282514 167385
rect 282458 167311 282514 167320
rect 282656 167074 282684 167855
rect 282644 167068 282696 167074
rect 282644 167010 282696 167016
rect 282644 164144 282696 164150
rect 282644 164086 282696 164092
rect 282656 163033 282684 164086
rect 282642 163024 282698 163033
rect 282642 162959 282698 162968
rect 282644 162852 282696 162858
rect 282644 162794 282696 162800
rect 282656 161945 282684 162794
rect 282642 161936 282698 161945
rect 282642 161871 282698 161880
rect 282366 100192 282422 100201
rect 282366 100127 282422 100136
rect 281630 87544 281686 87553
rect 281630 87479 281686 87488
rect 282182 84824 282238 84833
rect 282182 84759 282238 84768
rect 280986 3768 281042 3777
rect 280986 3703 281042 3712
rect 282196 3369 282224 84759
rect 282748 79529 282776 215727
rect 282918 197432 282974 197441
rect 282918 197367 282974 197376
rect 282826 192400 282882 192409
rect 282826 192335 282882 192344
rect 282840 191894 282868 192335
rect 282828 191888 282880 191894
rect 282828 191830 282880 191836
rect 282826 170640 282882 170649
rect 282826 170575 282882 170584
rect 282840 169794 282868 170575
rect 282828 169788 282880 169794
rect 282828 169730 282880 169736
rect 282826 168464 282882 168473
rect 282826 168399 282828 168408
rect 282880 168399 282882 168408
rect 282828 168370 282880 168376
rect 282828 167000 282880 167006
rect 282828 166942 282880 166948
rect 282840 166841 282868 166942
rect 282826 166832 282882 166841
rect 282826 166767 282882 166776
rect 282828 165572 282880 165578
rect 282828 165514 282880 165520
rect 282840 165209 282868 165514
rect 282826 165200 282882 165209
rect 282826 165135 282882 165144
rect 282828 164212 282880 164218
rect 282828 164154 282880 164160
rect 282840 163577 282868 164154
rect 282826 163568 282882 163577
rect 282826 163503 282882 163512
rect 282828 162784 282880 162790
rect 282828 162726 282880 162732
rect 282840 162489 282868 162726
rect 282826 162480 282882 162489
rect 282826 162415 282882 162424
rect 282828 161424 282880 161430
rect 282826 161392 282828 161401
rect 282880 161392 282882 161401
rect 282826 161327 282882 161336
rect 282734 79520 282790 79529
rect 282734 79455 282790 79464
rect 282932 4049 282960 197367
rect 283024 119649 283052 293519
rect 283194 291952 283250 291961
rect 283194 291887 283250 291896
rect 283102 290320 283158 290329
rect 283102 290255 283158 290264
rect 283116 119814 283144 290255
rect 283208 120698 283236 291887
rect 283300 244633 283328 348599
rect 283392 260953 283420 349182
rect 284298 348936 284354 348945
rect 284298 348871 284354 348880
rect 284312 348294 284340 348871
rect 284300 348288 284352 348294
rect 284300 348230 284352 348236
rect 284666 348256 284722 348265
rect 284666 348191 284722 348200
rect 283654 347304 283710 347313
rect 283654 347239 283710 347248
rect 283470 342680 283526 342689
rect 283470 342615 283526 342624
rect 283484 266393 283512 342615
rect 283564 339788 283616 339794
rect 283564 339730 283616 339736
rect 283576 306105 283604 339730
rect 283562 306096 283618 306105
rect 283562 306031 283618 306040
rect 283562 295352 283618 295361
rect 283562 295287 283618 295296
rect 283470 266384 283526 266393
rect 283470 266319 283526 266328
rect 283378 260944 283434 260953
rect 283378 260879 283434 260888
rect 283286 244624 283342 244633
rect 283286 244559 283342 244568
rect 283576 237017 283604 295287
rect 283668 290601 283696 347239
rect 284300 345772 284352 345778
rect 284300 345714 284352 345720
rect 284312 345681 284340 345714
rect 284298 345672 284354 345681
rect 284298 345607 284354 345616
rect 284300 339720 284352 339726
rect 284300 339662 284352 339668
rect 283748 339448 283800 339454
rect 283748 339390 283800 339396
rect 283838 339416 283894 339425
rect 283654 290592 283710 290601
rect 283654 290527 283710 290536
rect 283562 237008 283618 237017
rect 283562 236943 283618 236952
rect 283760 235958 283788 339390
rect 283838 339351 283894 339360
rect 283852 338881 283880 339351
rect 283838 338872 283894 338881
rect 283838 338807 283894 338816
rect 284312 307766 284340 339662
rect 284300 307760 284352 307766
rect 284300 307702 284352 307708
rect 284390 294672 284446 294681
rect 284390 294607 284446 294616
rect 284300 292596 284352 292602
rect 284300 292538 284352 292544
rect 283748 235952 283800 235958
rect 283748 235894 283800 235900
rect 283562 219600 283618 219609
rect 283562 219535 283618 219544
rect 283378 209808 283434 209817
rect 283378 209743 283434 209752
rect 283286 179072 283342 179081
rect 283286 179007 283342 179016
rect 283300 178673 283328 179007
rect 283286 178664 283342 178673
rect 283286 178599 283342 178608
rect 283286 169824 283342 169833
rect 283286 169759 283342 169768
rect 283196 120692 283248 120698
rect 283196 120634 283248 120640
rect 283104 119808 283156 119814
rect 283104 119750 283156 119756
rect 283010 119640 283066 119649
rect 283010 119575 283066 119584
rect 283102 6216 283158 6225
rect 283102 6151 283158 6160
rect 282918 4040 282974 4049
rect 282918 3975 282974 3984
rect 282182 3360 282238 3369
rect 282182 3295 282238 3304
rect 280066 3224 280122 3233
rect 280066 3159 280122 3168
rect 283116 480 283144 6151
rect 283300 3505 283328 169759
rect 283392 76537 283420 209743
rect 283470 209264 283526 209273
rect 283470 209199 283526 209208
rect 283484 77897 283512 209199
rect 283576 107137 283604 219535
rect 283746 213072 283802 213081
rect 283746 213007 283802 213016
rect 283654 193488 283710 193497
rect 283654 193423 283710 193432
rect 283562 107128 283618 107137
rect 283562 107063 283618 107072
rect 283668 89049 283696 193423
rect 283760 108361 283788 213007
rect 284312 120170 284340 292538
rect 284404 121009 284432 294607
rect 284484 291236 284536 291242
rect 284484 291178 284536 291184
rect 284390 121000 284446 121009
rect 284390 120935 284446 120944
rect 284312 120142 284432 120170
rect 284298 120048 284354 120057
rect 284298 119983 284354 119992
rect 284312 119882 284340 119983
rect 284300 119876 284352 119882
rect 284300 119818 284352 119824
rect 284404 119542 284432 120142
rect 284392 119536 284444 119542
rect 284392 119478 284444 119484
rect 284496 119474 284524 291178
rect 284576 289876 284628 289882
rect 284576 289818 284628 289824
rect 284588 119610 284616 289818
rect 284680 236473 284708 348191
rect 284772 243001 284800 349415
rect 284852 339244 284904 339250
rect 284852 339186 284904 339192
rect 284864 269074 284892 339186
rect 284956 285161 284984 372263
rect 285036 344208 285088 344214
rect 285036 344150 285088 344156
rect 284942 285152 284998 285161
rect 284942 285087 284998 285096
rect 285048 277370 285076 344150
rect 285140 337385 285168 390116
rect 286690 386880 286746 386889
rect 286690 386815 286746 386824
rect 286506 384704 286562 384713
rect 286506 384639 286562 384648
rect 286322 379264 286378 379273
rect 286322 379199 286378 379208
rect 285218 347168 285274 347177
rect 285218 347103 285274 347112
rect 285126 337376 285182 337385
rect 285126 337311 285182 337320
rect 285232 289513 285260 347103
rect 285772 346996 285824 347002
rect 285772 346938 285824 346944
rect 285310 344584 285366 344593
rect 285310 344519 285366 344528
rect 285324 322153 285352 344519
rect 285402 341728 285458 341737
rect 285402 341663 285458 341672
rect 285310 322144 285366 322153
rect 285310 322079 285366 322088
rect 285416 321065 285444 341663
rect 285680 341556 285732 341562
rect 285680 341498 285732 341504
rect 285692 341193 285720 341498
rect 285678 341184 285734 341193
rect 285678 341119 285734 341128
rect 285784 335354 285812 346938
rect 285954 342408 286010 342417
rect 285954 342343 286010 342352
rect 285864 341692 285916 341698
rect 285864 341634 285916 341640
rect 285692 335326 285812 335354
rect 285402 321056 285458 321065
rect 285402 320991 285458 321000
rect 285218 289504 285274 289513
rect 285218 289439 285274 289448
rect 285036 277364 285088 277370
rect 285036 277306 285088 277312
rect 284852 269068 284904 269074
rect 284852 269010 284904 269016
rect 285692 251054 285720 335326
rect 285770 295760 285826 295769
rect 285770 295695 285826 295704
rect 285680 251048 285732 251054
rect 285680 250990 285732 250996
rect 284758 242992 284814 243001
rect 284758 242927 284814 242936
rect 284666 236464 284722 236473
rect 284666 236399 284722 236408
rect 285034 227760 285090 227769
rect 285034 227695 285090 227704
rect 284758 220144 284814 220153
rect 284758 220079 284814 220088
rect 284666 203824 284722 203833
rect 284666 203759 284722 203768
rect 284576 119604 284628 119610
rect 284576 119546 284628 119552
rect 284484 119468 284536 119474
rect 284484 119410 284536 119416
rect 283746 108352 283802 108361
rect 283746 108287 283802 108296
rect 283654 89040 283710 89049
rect 283654 88975 283710 88984
rect 283470 77888 283526 77897
rect 283470 77823 283526 77832
rect 283378 76528 283434 76537
rect 283378 76463 283434 76472
rect 284680 64161 284708 203759
rect 284772 94761 284800 220079
rect 284850 213616 284906 213625
rect 284850 213551 284906 213560
rect 284758 94752 284814 94761
rect 284758 94687 284814 94696
rect 284864 91905 284892 213551
rect 284942 210896 284998 210905
rect 284942 210831 284998 210840
rect 284956 93265 284984 210831
rect 285048 113665 285076 227695
rect 285678 225584 285734 225593
rect 285678 225519 285734 225528
rect 285126 221232 285182 221241
rect 285126 221167 285182 221176
rect 285034 113656 285090 113665
rect 285034 113591 285090 113600
rect 285140 108633 285168 221167
rect 285126 108624 285182 108633
rect 285126 108559 285182 108568
rect 284942 93256 284998 93265
rect 284942 93191 284998 93200
rect 284850 91896 284906 91905
rect 284850 91831 284906 91840
rect 284666 64152 284722 64161
rect 284666 64087 284722 64096
rect 284942 43616 284998 43625
rect 284942 43551 284998 43560
rect 284956 3641 284984 43551
rect 285692 7721 285720 225519
rect 285784 121145 285812 295695
rect 285876 248130 285904 341634
rect 285968 266937 285996 342343
rect 285954 266928 286010 266937
rect 285954 266863 286010 266872
rect 285864 248124 285916 248130
rect 285864 248066 285916 248072
rect 286230 229936 286286 229945
rect 286230 229871 286286 229880
rect 285954 225040 286010 225049
rect 285954 224975 286010 224984
rect 285862 212528 285918 212537
rect 285862 212463 285918 212472
rect 285770 121136 285826 121145
rect 285770 121071 285826 121080
rect 285876 73817 285904 212463
rect 285968 104417 285996 224975
rect 286138 223952 286194 223961
rect 286138 223887 286194 223896
rect 286046 222864 286102 222873
rect 286046 222799 286102 222808
rect 286060 105777 286088 222799
rect 286152 108497 286180 223887
rect 286244 118017 286272 229871
rect 286336 229673 286364 379199
rect 286414 365256 286470 365265
rect 286414 365191 286470 365200
rect 286322 229664 286378 229673
rect 286322 229599 286378 229608
rect 286428 219881 286456 365191
rect 286520 248169 286548 384639
rect 286600 342644 286652 342650
rect 286600 342586 286652 342592
rect 286612 255270 286640 342586
rect 286704 329769 286732 386815
rect 286782 345808 286838 345817
rect 286782 345743 286838 345752
rect 286690 329760 286746 329769
rect 286690 329695 286746 329704
rect 286796 311273 286824 345743
rect 286888 337521 286916 390116
rect 288162 386336 288218 386345
rect 288162 386271 288218 386280
rect 287704 384396 287756 384402
rect 287704 384338 287756 384344
rect 287716 375358 287744 384338
rect 287704 375352 287756 375358
rect 287704 375294 287756 375300
rect 288070 370968 288126 370977
rect 288070 370903 288126 370912
rect 287702 355600 287758 355609
rect 287702 355535 287758 355544
rect 287150 351520 287206 351529
rect 287150 351455 287206 351464
rect 287058 349344 287114 349353
rect 287058 349279 287114 349288
rect 286874 337512 286930 337521
rect 286874 337447 286930 337456
rect 286782 311264 286838 311273
rect 286782 311199 286838 311208
rect 286600 255264 286652 255270
rect 286600 255206 286652 255212
rect 286506 248160 286562 248169
rect 286506 248095 286562 248104
rect 287072 242457 287100 349279
rect 287164 295361 287192 351455
rect 287244 344412 287296 344418
rect 287244 344354 287296 344360
rect 287150 295352 287206 295361
rect 287150 295287 287206 295296
rect 287150 295216 287206 295225
rect 287150 295151 287206 295160
rect 287058 242448 287114 242457
rect 287058 242383 287114 242392
rect 286414 219872 286470 219881
rect 286414 219807 286470 219816
rect 286414 211984 286470 211993
rect 286414 211919 286470 211928
rect 286322 211440 286378 211449
rect 286322 211375 286378 211384
rect 286230 118008 286286 118017
rect 286230 117943 286286 117952
rect 286336 109857 286364 211375
rect 286428 114073 286456 211919
rect 286506 205456 286562 205465
rect 286506 205391 286562 205400
rect 286520 116521 286548 205391
rect 287058 201104 287114 201113
rect 287058 201039 287114 201048
rect 286506 116512 286562 116521
rect 286506 116447 286562 116456
rect 286414 114064 286470 114073
rect 286414 113999 286470 114008
rect 286322 109848 286378 109857
rect 286322 109783 286378 109792
rect 286138 108488 286194 108497
rect 286138 108423 286194 108432
rect 286046 105768 286102 105777
rect 286046 105703 286102 105712
rect 285954 104408 286010 104417
rect 285954 104343 286010 104352
rect 285862 73808 285918 73817
rect 285862 73743 285918 73752
rect 285678 7712 285734 7721
rect 285678 7647 285734 7656
rect 286598 5672 286654 5681
rect 286598 5607 286654 5616
rect 284942 3632 284998 3641
rect 284942 3567 284998 3576
rect 283286 3496 283342 3505
rect 283286 3431 283342 3440
rect 286612 480 286640 5607
rect 287072 5001 287100 201039
rect 287164 119105 287192 295151
rect 287256 269006 287284 344354
rect 287244 269000 287296 269006
rect 287244 268942 287296 268948
rect 287610 206544 287666 206553
rect 287610 206479 287666 206488
rect 287518 204368 287574 204377
rect 287518 204303 287574 204312
rect 287426 202736 287482 202745
rect 287426 202671 287482 202680
rect 287334 201648 287390 201657
rect 287334 201583 287390 201592
rect 287242 200560 287298 200569
rect 287242 200495 287298 200504
rect 287150 119096 287206 119105
rect 287150 119031 287206 119040
rect 287256 46209 287284 200495
rect 287348 50289 287376 201583
rect 287440 72457 287468 202671
rect 287532 105505 287560 204303
rect 287624 111081 287652 206479
rect 287716 198121 287744 355535
rect 287886 349752 287942 349761
rect 287886 349687 287942 349696
rect 287796 348016 287848 348022
rect 287796 347958 287848 347964
rect 287702 198112 287758 198121
rect 287702 198047 287758 198056
rect 287808 195974 287836 347958
rect 287900 215529 287928 349687
rect 287980 342576 288032 342582
rect 287980 342518 288032 342524
rect 287992 218006 288020 342518
rect 288084 263401 288112 370903
rect 288176 318889 288204 386271
rect 288440 351960 288492 351966
rect 288440 351902 288492 351908
rect 288254 341864 288310 341873
rect 288254 341799 288310 341808
rect 288162 318880 288218 318889
rect 288162 318815 288218 318824
rect 288268 313449 288296 341799
rect 288254 313440 288310 313449
rect 288254 313375 288310 313384
rect 288070 263392 288126 263401
rect 288070 263327 288126 263336
rect 287980 218000 288032 218006
rect 287980 217942 288032 217948
rect 287886 215520 287942 215529
rect 287886 215455 287942 215464
rect 287886 202192 287942 202201
rect 287886 202127 287942 202136
rect 287796 195968 287848 195974
rect 287796 195910 287848 195916
rect 287900 112577 287928 202127
rect 288452 162790 288480 351902
rect 288530 349616 288586 349625
rect 288530 349551 288586 349560
rect 288544 247353 288572 349551
rect 288636 337929 288664 390116
rect 289174 381848 289230 381857
rect 289174 381783 289230 381792
rect 289084 358896 289136 358902
rect 289084 358838 289136 358844
rect 288716 350804 288768 350810
rect 288716 350746 288768 350752
rect 288622 337920 288678 337929
rect 288622 337855 288678 337864
rect 288728 262206 288756 350746
rect 288716 262200 288768 262206
rect 288716 262142 288768 262148
rect 288530 247344 288586 247353
rect 288530 247279 288586 247288
rect 288714 208176 288770 208185
rect 288714 208111 288770 208120
rect 288622 207632 288678 207641
rect 288622 207567 288678 207576
rect 288530 207088 288586 207097
rect 288530 207023 288586 207032
rect 288440 162784 288492 162790
rect 288440 162726 288492 162732
rect 287886 112568 287942 112577
rect 287886 112503 287942 112512
rect 287610 111072 287666 111081
rect 287610 111007 287666 111016
rect 287518 105496 287574 105505
rect 287518 105431 287574 105440
rect 287426 72448 287482 72457
rect 287426 72383 287482 72392
rect 288544 58721 288572 207023
rect 288636 60081 288664 207567
rect 288728 61441 288756 208111
rect 289096 205630 289124 358838
rect 289188 236201 289216 381783
rect 289450 352744 289506 352753
rect 289450 352679 289506 352688
rect 289268 346656 289320 346662
rect 289268 346598 289320 346604
rect 289174 236192 289230 236201
rect 289174 236127 289230 236136
rect 289280 206990 289308 346598
rect 289360 345500 289412 345506
rect 289360 345442 289412 345448
rect 289372 208350 289400 345442
rect 289464 218793 289492 352679
rect 290094 348120 290150 348129
rect 290094 348055 290150 348064
rect 289544 339856 289596 339862
rect 289544 339798 289596 339804
rect 289556 273222 289584 339798
rect 289912 338292 289964 338298
rect 289912 338234 289964 338240
rect 289544 273216 289596 273222
rect 289544 273158 289596 273164
rect 289924 247042 289952 338234
rect 290002 338056 290058 338065
rect 290002 337991 290058 338000
rect 289912 247036 289964 247042
rect 289912 246978 289964 246984
rect 290016 246265 290044 337991
rect 290108 260409 290136 348055
rect 290384 334121 290412 390116
rect 292132 387598 292160 390116
rect 292120 387592 292172 387598
rect 292120 387534 292172 387540
rect 293880 387054 293908 390116
rect 294604 389904 294656 389910
rect 294604 389846 294656 389852
rect 293868 387048 293920 387054
rect 293868 386990 293920 386996
rect 292118 384840 292174 384849
rect 292118 384775 292174 384784
rect 292026 383344 292082 383353
rect 292026 383279 292082 383288
rect 291842 380488 291898 380497
rect 291842 380423 291898 380432
rect 290738 375320 290794 375329
rect 290738 375255 290794 375264
rect 290462 373824 290518 373833
rect 290462 373759 290518 373768
rect 290370 334112 290426 334121
rect 290370 334047 290426 334056
rect 290186 299432 290242 299441
rect 290186 299367 290242 299376
rect 290094 260400 290150 260409
rect 290094 260335 290150 260344
rect 290002 246256 290058 246265
rect 290002 246191 290058 246200
rect 289450 218784 289506 218793
rect 289450 218719 289506 218728
rect 289910 214160 289966 214169
rect 289910 214095 289966 214104
rect 289360 208344 289412 208350
rect 289360 208286 289412 208292
rect 289268 206984 289320 206990
rect 289268 206926 289320 206932
rect 289084 205624 289136 205630
rect 289084 205566 289136 205572
rect 288898 196208 288954 196217
rect 288898 196143 288954 196152
rect 288806 195120 288862 195129
rect 288806 195055 288862 195064
rect 288820 90409 288848 195055
rect 288912 102785 288940 196143
rect 289082 195664 289138 195673
rect 289082 195599 289138 195608
rect 288990 194576 289046 194585
rect 288990 194511 289046 194520
rect 288898 102776 288954 102785
rect 288898 102711 288954 102720
rect 289004 101425 289032 194511
rect 289096 106865 289124 195599
rect 289820 167068 289872 167074
rect 289820 167010 289872 167016
rect 289832 119950 289860 167010
rect 289820 119944 289872 119950
rect 289820 119886 289872 119892
rect 289924 114209 289952 214095
rect 290004 169788 290056 169794
rect 290004 169730 290056 169736
rect 290016 114510 290044 169730
rect 290096 168428 290148 168434
rect 290096 168370 290148 168376
rect 290108 120562 290136 168370
rect 290200 161430 290228 299367
rect 290476 240553 290504 373759
rect 290556 350872 290608 350878
rect 290556 350814 290608 350820
rect 290462 240544 290518 240553
rect 290462 240479 290518 240488
rect 290568 223582 290596 350814
rect 290648 348220 290700 348226
rect 290648 348162 290700 348168
rect 290660 270502 290688 348162
rect 290752 299305 290780 375255
rect 291568 350736 291620 350742
rect 291568 350678 291620 350684
rect 291200 346724 291252 346730
rect 291200 346666 291252 346672
rect 290738 299296 290794 299305
rect 290738 299231 290794 299240
rect 290648 270496 290700 270502
rect 290648 270438 290700 270444
rect 290556 223576 290608 223582
rect 290556 223518 290608 223524
rect 291212 168366 291240 346666
rect 291476 338224 291528 338230
rect 291476 338166 291528 338172
rect 291382 301200 291438 301209
rect 291382 301135 291438 301144
rect 291290 294128 291346 294137
rect 291290 294063 291346 294072
rect 291200 168360 291252 168366
rect 291200 168302 291252 168308
rect 290188 161424 290240 161430
rect 290188 161366 290240 161372
rect 290096 120556 290148 120562
rect 290096 120498 290148 120504
rect 291304 119377 291332 294063
rect 291396 131209 291424 301135
rect 291488 238746 291516 338166
rect 291580 263498 291608 350678
rect 291568 263492 291620 263498
rect 291568 263434 291620 263440
rect 291476 238740 291528 238746
rect 291476 238682 291528 238688
rect 291474 199472 291530 199481
rect 291474 199407 291530 199416
rect 291382 131200 291438 131209
rect 291382 131135 291438 131144
rect 291290 119368 291346 119377
rect 291290 119303 291346 119312
rect 290004 114504 290056 114510
rect 290004 114446 290056 114452
rect 289910 114200 289966 114209
rect 289910 114135 289966 114144
rect 289082 106856 289138 106865
rect 289082 106791 289138 106800
rect 288990 101416 289046 101425
rect 288990 101351 289046 101360
rect 288806 90400 288862 90409
rect 288806 90335 288862 90344
rect 288714 61432 288770 61441
rect 288714 61367 288770 61376
rect 288622 60072 288678 60081
rect 288622 60007 288678 60016
rect 288530 58712 288586 58721
rect 288530 58647 288586 58656
rect 287702 55720 287758 55729
rect 287702 55655 287758 55664
rect 287334 50280 287390 50289
rect 287334 50215 287390 50224
rect 287242 46200 287298 46209
rect 287242 46135 287298 46144
rect 287058 4992 287114 5001
rect 287058 4927 287114 4936
rect 287716 4865 287744 55655
rect 291488 49201 291516 199407
rect 291856 197033 291884 380423
rect 291934 370832 291990 370841
rect 291934 370767 291990 370776
rect 291948 232937 291976 370767
rect 292040 267753 292068 383279
rect 292132 328681 292160 384775
rect 294616 382974 294644 389846
rect 294694 383072 294750 383081
rect 294694 383007 294750 383016
rect 294604 382968 294656 382974
rect 294604 382910 294656 382916
rect 293222 377632 293278 377641
rect 293222 377567 293278 377576
rect 292580 349376 292632 349382
rect 292580 349318 292632 349324
rect 292302 345944 292358 345953
rect 292302 345879 292358 345888
rect 292210 344448 292266 344457
rect 292210 344383 292266 344392
rect 292118 328672 292174 328681
rect 292118 328607 292174 328616
rect 292224 304745 292252 344383
rect 292316 315625 292344 345879
rect 292302 315616 292358 315625
rect 292302 315551 292358 315560
rect 292210 304736 292266 304745
rect 292210 304671 292266 304680
rect 292026 267744 292082 267753
rect 292026 267679 292082 267688
rect 292592 253774 292620 349318
rect 292856 347880 292908 347886
rect 292856 347822 292908 347828
rect 292764 344276 292816 344282
rect 292764 344218 292816 344224
rect 292672 298172 292724 298178
rect 292672 298114 292724 298120
rect 292580 253768 292632 253774
rect 292580 253710 292632 253716
rect 291934 232928 291990 232937
rect 291934 232863 291990 232872
rect 291842 197024 291898 197033
rect 291842 196959 291898 196968
rect 292580 191888 292632 191894
rect 292580 191830 292632 191836
rect 291566 170096 291622 170105
rect 291566 170031 291622 170040
rect 291580 118833 291608 170031
rect 291842 160712 291898 160721
rect 291842 160647 291898 160656
rect 291856 153241 291884 160647
rect 291842 153232 291898 153241
rect 291842 153167 291898 153176
rect 291566 118824 291622 118833
rect 291566 118759 291622 118768
rect 291842 118144 291898 118153
rect 291842 118079 291898 118088
rect 291856 100609 291884 118079
rect 291842 100600 291898 100609
rect 291842 100535 291898 100544
rect 291474 49192 291530 49201
rect 291474 49127 291530 49136
rect 289082 42256 289138 42265
rect 289082 42191 289138 42200
rect 287702 4856 287758 4865
rect 287702 4791 287758 4800
rect 289096 3505 289124 42191
rect 290186 19952 290242 19961
rect 290186 19887 290242 19896
rect 289082 3496 289138 3505
rect 289082 3431 289138 3440
rect 290200 480 290228 19887
rect 292592 4146 292620 191830
rect 292684 118114 292712 298114
rect 292776 249694 292804 344218
rect 292868 259282 292896 347822
rect 292948 338360 293000 338366
rect 292948 338302 293000 338308
rect 292960 263566 292988 338302
rect 292948 263560 293000 263566
rect 292948 263502 293000 263508
rect 292856 259276 292908 259282
rect 292856 259218 292908 259224
rect 292764 249688 292816 249694
rect 292764 249630 292816 249636
rect 293236 234025 293264 377567
rect 294604 375352 294656 375358
rect 294604 375294 294656 375300
rect 294616 366722 294644 375294
rect 293592 366716 293644 366722
rect 293592 366658 293644 366664
rect 294604 366716 294656 366722
rect 294604 366658 294656 366664
rect 293498 362944 293554 362953
rect 293498 362879 293554 362888
rect 293406 350024 293462 350033
rect 293406 349959 293462 349968
rect 293316 344140 293368 344146
rect 293316 344082 293368 344088
rect 293328 235958 293356 344082
rect 293420 262313 293448 349959
rect 293512 284073 293540 362879
rect 293604 344350 293632 366658
rect 294604 358828 294656 358834
rect 294604 358770 294656 358776
rect 293592 344344 293644 344350
rect 293592 344286 293644 344292
rect 294142 342272 294198 342281
rect 294142 342207 294198 342216
rect 293958 299024 294014 299033
rect 293958 298959 294014 298968
rect 293498 284064 293554 284073
rect 293498 283999 293554 284008
rect 293406 262304 293462 262313
rect 293406 262239 293462 262248
rect 293316 235952 293368 235958
rect 293316 235894 293368 235900
rect 293222 234016 293278 234025
rect 293222 233951 293278 233960
rect 292762 210352 292818 210361
rect 292762 210287 292818 210296
rect 292672 118108 292724 118114
rect 292672 118050 292724 118056
rect 292776 113937 292804 210287
rect 293972 125497 294000 298959
rect 294052 288448 294104 288454
rect 294052 288390 294104 288396
rect 293958 125488 294014 125497
rect 293958 125423 294014 125432
rect 294064 118182 294092 288390
rect 294156 267481 294184 342207
rect 294234 341456 294290 341465
rect 294234 341391 294290 341400
rect 294142 267472 294198 267481
rect 294142 267407 294198 267416
rect 294248 265849 294276 341391
rect 294328 338972 294380 338978
rect 294328 338914 294380 338920
rect 294234 265840 294290 265849
rect 294234 265775 294290 265784
rect 294340 264926 294368 338914
rect 294328 264920 294380 264926
rect 294328 264862 294380 264868
rect 294142 206000 294198 206009
rect 294142 205935 294198 205944
rect 294052 118176 294104 118182
rect 294052 118118 294104 118124
rect 292762 113928 292818 113937
rect 292762 113863 292818 113872
rect 294156 113801 294184 205935
rect 294616 201482 294644 358770
rect 294708 238377 294736 383007
rect 294878 378040 294934 378049
rect 294878 377975 294934 377984
rect 294788 339652 294840 339658
rect 294788 339594 294840 339600
rect 294694 238368 294750 238377
rect 294694 238303 294750 238312
rect 294800 226302 294828 339594
rect 294892 266665 294920 377975
rect 294970 372464 295026 372473
rect 294970 372399 295026 372408
rect 294984 300393 295012 372399
rect 295340 353388 295392 353394
rect 295340 353330 295392 353336
rect 295062 346080 295118 346089
rect 295062 346015 295118 346024
rect 295076 324329 295104 346015
rect 295062 324320 295118 324329
rect 295062 324255 295118 324264
rect 294970 300384 295026 300393
rect 294970 300319 295026 300328
rect 294878 266656 294934 266665
rect 294878 266591 294934 266600
rect 294788 226296 294840 226302
rect 294788 226238 294840 226244
rect 294604 201476 294656 201482
rect 294604 201418 294656 201424
rect 295352 164150 295380 353330
rect 295524 345636 295576 345642
rect 295524 345578 295576 345584
rect 295430 337920 295486 337929
rect 295430 337855 295486 337864
rect 295444 333033 295472 337855
rect 295430 333024 295486 333033
rect 295430 332959 295486 332968
rect 295430 299568 295486 299577
rect 295430 299503 295486 299512
rect 295340 164144 295392 164150
rect 295340 164086 295392 164092
rect 295444 120601 295472 299503
rect 295536 249762 295564 345578
rect 295524 249756 295576 249762
rect 295524 249698 295576 249704
rect 295628 146985 295656 390116
rect 296166 381984 296222 381993
rect 296166 381919 296222 381928
rect 295982 376544 296038 376553
rect 295982 376479 296038 376488
rect 295708 341760 295760 341766
rect 295708 341702 295760 341708
rect 295720 266354 295748 341702
rect 295798 336288 295854 336297
rect 295798 336223 295854 336232
rect 295708 266348 295760 266354
rect 295708 266290 295760 266296
rect 295812 263673 295840 336223
rect 295798 263664 295854 263673
rect 295798 263599 295854 263608
rect 295996 241641 296024 376479
rect 296076 348084 296128 348090
rect 296076 348026 296128 348032
rect 295982 241632 296038 241641
rect 295982 241567 296038 241576
rect 296088 224942 296116 348026
rect 296180 265577 296208 381919
rect 296812 353456 296864 353462
rect 296812 353398 296864 353404
rect 296720 353320 296772 353326
rect 296720 353262 296772 353268
rect 296258 352472 296314 352481
rect 296258 352407 296314 352416
rect 296272 297129 296300 352407
rect 296258 297120 296314 297129
rect 296258 297055 296314 297064
rect 296166 265568 296222 265577
rect 296166 265503 296222 265512
rect 296076 224936 296128 224942
rect 296076 224878 296128 224884
rect 296732 164218 296760 353262
rect 296824 165578 296852 353398
rect 296994 345264 297050 345273
rect 296904 345228 296956 345234
rect 296994 345199 297050 345208
rect 296904 345170 296956 345176
rect 296916 256562 296944 345170
rect 297008 269657 297036 345199
rect 296994 269648 297050 269657
rect 296994 269583 297050 269592
rect 296904 256556 296956 256562
rect 296904 256498 296956 256504
rect 296812 165572 296864 165578
rect 296812 165514 296864 165520
rect 296720 164212 296772 164218
rect 296720 164154 296772 164160
rect 297376 147393 297404 390116
rect 297454 369336 297510 369345
rect 297454 369271 297510 369280
rect 297468 274281 297496 369271
rect 298742 367704 298798 367713
rect 298742 367639 298798 367648
rect 298100 350396 298152 350402
rect 298100 350338 298152 350344
rect 298112 349217 298140 350338
rect 298098 349208 298154 349217
rect 298098 349143 298154 349152
rect 298284 346928 298336 346934
rect 298284 346870 298336 346876
rect 298192 345568 298244 345574
rect 298192 345510 298244 345516
rect 298100 339516 298152 339522
rect 298100 339458 298152 339464
rect 297546 339144 297602 339153
rect 297546 339079 297602 339088
rect 297560 326505 297588 339079
rect 297546 326496 297602 326505
rect 297546 326431 297602 326440
rect 297454 274272 297510 274281
rect 297454 274207 297510 274216
rect 298112 251122 298140 339458
rect 298204 256630 298232 345510
rect 298296 257990 298324 346870
rect 298376 338904 298428 338910
rect 298376 338846 298428 338852
rect 298284 257984 298336 257990
rect 298284 257926 298336 257932
rect 298192 256624 298244 256630
rect 298192 256566 298244 256572
rect 298388 253842 298416 338846
rect 298376 253836 298428 253842
rect 298376 253778 298428 253784
rect 298100 251116 298152 251122
rect 298100 251058 298152 251064
rect 298756 227497 298784 367639
rect 299018 366752 299074 366761
rect 299018 366687 299074 366696
rect 298926 365392 298982 365401
rect 298926 365327 298982 365336
rect 298836 347948 298888 347954
rect 298836 347890 298888 347896
rect 298742 227488 298798 227497
rect 298742 227423 298798 227432
rect 298848 212498 298876 347890
rect 298940 249257 298968 365327
rect 299032 286249 299060 366687
rect 299018 286240 299074 286249
rect 299018 286175 299074 286184
rect 298926 249248 298982 249257
rect 298926 249183 298982 249192
rect 299124 244934 299152 390116
rect 300122 385792 300178 385801
rect 300122 385727 300178 385736
rect 299572 348152 299624 348158
rect 299572 348094 299624 348100
rect 299480 345432 299532 345438
rect 299480 345374 299532 345380
rect 299202 343224 299258 343233
rect 299202 343159 299258 343168
rect 299216 312361 299244 343159
rect 299202 312352 299258 312361
rect 299202 312287 299258 312296
rect 299492 256698 299520 345374
rect 299584 259350 299612 348094
rect 299662 336152 299718 336161
rect 299662 336087 299718 336096
rect 299572 259344 299624 259350
rect 299572 259286 299624 259292
rect 299676 258058 299704 336087
rect 299664 258052 299716 258058
rect 299664 257994 299716 258000
rect 299480 256692 299532 256698
rect 299480 256634 299532 256640
rect 299112 244928 299164 244934
rect 299112 244870 299164 244876
rect 300136 213353 300164 385727
rect 300490 364304 300546 364313
rect 300490 364239 300546 364248
rect 300306 361448 300362 361457
rect 300306 361383 300362 361392
rect 300214 349888 300270 349897
rect 300214 349823 300270 349832
rect 300228 231849 300256 349823
rect 300320 251433 300348 361383
rect 300400 341488 300452 341494
rect 300400 341430 300452 341436
rect 300412 256698 300440 341430
rect 300504 294953 300532 364239
rect 300582 347440 300638 347449
rect 300582 347375 300638 347384
rect 300596 319977 300624 347375
rect 300582 319968 300638 319977
rect 300582 319903 300638 319912
rect 300872 299441 300900 390116
rect 302634 390102 302924 390130
rect 306130 390116 306328 390130
rect 307878 390116 308168 390130
rect 302896 386442 302924 390102
rect 304368 389065 304396 390116
rect 306116 390102 306328 390116
rect 307864 390102 308168 390116
rect 309626 390102 309824 390130
rect 304354 389056 304410 389065
rect 304354 388991 304410 389000
rect 302884 386436 302936 386442
rect 302884 386378 302936 386384
rect 301594 372056 301650 372065
rect 301594 371991 301650 372000
rect 301502 353016 301558 353025
rect 301502 352951 301558 352960
rect 301134 350568 301190 350577
rect 301134 350503 301190 350512
rect 301044 348356 301096 348362
rect 301044 348298 301096 348304
rect 300952 339924 301004 339930
rect 300952 339866 301004 339872
rect 300858 299432 300914 299441
rect 300858 299367 300914 299376
rect 300490 294944 300546 294953
rect 300490 294879 300546 294888
rect 300400 256692 300452 256698
rect 300400 256634 300452 256640
rect 300964 252482 300992 339866
rect 301056 260846 301084 348298
rect 301148 264761 301176 350503
rect 301228 338836 301280 338842
rect 301228 338778 301280 338784
rect 301134 264752 301190 264761
rect 301134 264687 301190 264696
rect 301044 260840 301096 260846
rect 301044 260782 301096 260788
rect 301240 255202 301268 338778
rect 301228 255196 301280 255202
rect 301228 255138 301280 255144
rect 300952 252476 301004 252482
rect 300952 252418 301004 252424
rect 300306 251424 300362 251433
rect 300306 251359 300362 251368
rect 301516 245993 301544 352951
rect 301608 268841 301636 371991
rect 302240 358352 302292 358358
rect 302240 358294 302292 358300
rect 301594 268832 301650 268841
rect 301594 268767 301650 268776
rect 301502 245984 301558 245993
rect 301502 245919 301558 245928
rect 300214 231840 300270 231849
rect 300214 231775 300270 231784
rect 300122 213344 300178 213353
rect 300122 213279 300178 213288
rect 298836 212492 298888 212498
rect 298836 212434 298888 212440
rect 298742 187776 298798 187785
rect 298742 187711 298798 187720
rect 298756 160313 298784 187711
rect 302252 162858 302280 358294
rect 302606 350704 302662 350713
rect 302606 350639 302662 350648
rect 302332 349172 302384 349178
rect 302332 349114 302384 349120
rect 302344 253910 302372 349114
rect 302516 348628 302568 348634
rect 302516 348570 302568 348576
rect 302424 340400 302476 340406
rect 302424 340342 302476 340348
rect 302332 253904 302384 253910
rect 302332 253846 302384 253852
rect 302436 251190 302464 340342
rect 302528 259418 302556 348570
rect 302620 261497 302648 350639
rect 302896 343670 302924 386378
rect 304262 380352 304318 380361
rect 304262 380287 304318 380296
rect 303250 369472 303306 369481
rect 303250 369407 303306 369416
rect 302974 366344 303030 366353
rect 302974 366279 303030 366288
rect 302884 343664 302936 343670
rect 302884 343606 302936 343612
rect 302606 261488 302662 261497
rect 302606 261423 302662 261432
rect 302516 259412 302568 259418
rect 302516 259354 302568 259360
rect 302424 251184 302476 251190
rect 302424 251126 302476 251132
rect 302896 164898 302924 343606
rect 302988 228585 303016 366279
rect 303158 364168 303214 364177
rect 303158 364103 303214 364112
rect 303068 346588 303120 346594
rect 303068 346530 303120 346536
rect 302974 228576 303030 228585
rect 302974 228511 303030 228520
rect 303080 215286 303108 346530
rect 303172 252521 303200 364103
rect 303264 292777 303292 369407
rect 303620 357468 303672 357474
rect 303620 357410 303672 357416
rect 303250 292768 303306 292777
rect 303250 292703 303306 292712
rect 303158 252512 303214 252521
rect 303158 252447 303214 252456
rect 303068 215280 303120 215286
rect 303068 215222 303120 215228
rect 303526 191720 303582 191729
rect 303526 191655 303582 191664
rect 303540 187785 303568 191655
rect 303526 187776 303582 187785
rect 303526 187711 303582 187720
rect 303632 167006 303660 357410
rect 303712 340468 303764 340474
rect 303712 340410 303764 340416
rect 303724 252550 303752 340410
rect 304170 337512 304226 337521
rect 304170 337447 304226 337456
rect 304184 331945 304212 337447
rect 304170 331936 304226 331945
rect 304170 331871 304226 331880
rect 303712 252544 303764 252550
rect 303712 252486 303764 252492
rect 304276 199209 304304 380287
rect 304368 345710 304396 388991
rect 305734 379400 305790 379409
rect 305734 379335 305790 379344
rect 304446 362536 304502 362545
rect 304446 362471 304502 362480
rect 304356 345704 304408 345710
rect 304356 345646 304408 345652
rect 304262 199200 304318 199209
rect 304262 199135 304318 199144
rect 304368 167657 304396 345646
rect 304460 253609 304488 362471
rect 304998 350976 305054 350985
rect 304998 350911 305054 350920
rect 304540 344344 304592 344350
rect 304540 344286 304592 344292
rect 304552 322930 304580 344286
rect 304540 322924 304592 322930
rect 304540 322866 304592 322872
rect 305012 254969 305040 350911
rect 305644 342508 305696 342514
rect 305644 342450 305696 342456
rect 304998 254960 305054 254969
rect 304998 254895 305054 254904
rect 304446 253600 304502 253609
rect 304446 253535 304502 253544
rect 305656 175982 305684 342450
rect 305748 259049 305776 379335
rect 305918 371104 305974 371113
rect 305918 371039 305974 371048
rect 305828 345296 305880 345302
rect 305828 345238 305880 345244
rect 305734 259040 305790 259049
rect 305734 258975 305790 258984
rect 305840 240106 305868 345238
rect 305932 296041 305960 371039
rect 306012 366716 306064 366722
rect 306012 366658 306064 366664
rect 306024 303618 306052 366658
rect 306116 342514 306144 390102
rect 307022 386064 307078 386073
rect 307022 385999 307078 386008
rect 306378 350840 306434 350849
rect 306378 350775 306434 350784
rect 306104 342508 306156 342514
rect 306104 342450 306156 342456
rect 306012 303612 306064 303618
rect 306012 303554 306064 303560
rect 305918 296032 305974 296041
rect 305918 295967 305974 295976
rect 305828 240100 305880 240106
rect 305828 240042 305880 240048
rect 306392 232665 306420 350775
rect 307036 237289 307064 385999
rect 307206 375048 307262 375057
rect 307206 374983 307262 374992
rect 307116 344004 307168 344010
rect 307116 343946 307168 343952
rect 307022 237280 307078 237289
rect 307022 237215 307078 237224
rect 306378 232656 306434 232665
rect 306378 232591 306434 232600
rect 307128 222154 307156 343946
rect 307220 264489 307248 374983
rect 307300 345364 307352 345370
rect 307300 345306 307352 345312
rect 307312 271862 307340 345306
rect 307864 341086 307892 390102
rect 308140 390046 308168 390102
rect 308128 390040 308180 390046
rect 308128 389982 308180 389988
rect 309796 389162 309824 390102
rect 311176 390102 311374 390130
rect 312556 390102 313122 390130
rect 309784 389156 309836 389162
rect 309784 389098 309836 389104
rect 308496 382968 308548 382974
rect 308496 382910 308548 382916
rect 307852 341080 307904 341086
rect 307852 341022 307904 341028
rect 308404 341080 308456 341086
rect 308404 341022 308456 341028
rect 307300 271856 307352 271862
rect 307300 271798 307352 271804
rect 307206 264480 307262 264489
rect 307206 264415 307262 264424
rect 307116 222148 307168 222154
rect 307116 222090 307168 222096
rect 305644 175976 305696 175982
rect 305644 175918 305696 175924
rect 308416 170406 308444 341022
rect 308508 218074 308536 382910
rect 308586 351248 308642 351257
rect 308586 351183 308642 351192
rect 308600 278633 308628 351183
rect 309796 341018 309824 389098
rect 311176 389094 311204 390102
rect 311164 389088 311216 389094
rect 311164 389030 311216 389036
rect 309874 375864 309930 375873
rect 309874 375799 309930 375808
rect 309784 341012 309836 341018
rect 309784 340954 309836 340960
rect 308680 322924 308732 322930
rect 308680 322866 308732 322872
rect 308586 278624 308642 278633
rect 308586 278559 308642 278568
rect 308692 250510 308720 322866
rect 309048 303612 309100 303618
rect 309048 303554 309100 303560
rect 309060 298110 309088 303554
rect 309048 298104 309100 298110
rect 309048 298046 309100 298052
rect 308680 250504 308732 250510
rect 308680 250446 308732 250452
rect 308496 218068 308548 218074
rect 308496 218010 308548 218016
rect 309046 195936 309102 195945
rect 309046 195871 309102 195880
rect 309060 191865 309088 195871
rect 309046 191856 309102 191865
rect 309046 191791 309102 191800
rect 308404 170400 308456 170406
rect 308404 170342 308456 170348
rect 308402 169824 308458 169833
rect 308402 169759 308458 169768
rect 304354 167648 304410 167657
rect 304354 167583 304410 167592
rect 303620 167000 303672 167006
rect 303620 166942 303672 166948
rect 302884 164892 302936 164898
rect 302884 164834 302936 164840
rect 308416 162897 308444 169759
rect 308402 162888 308458 162897
rect 302240 162852 302292 162858
rect 308402 162823 308458 162832
rect 302240 162794 302292 162800
rect 303986 162752 304042 162761
rect 303986 162687 304042 162696
rect 304000 160857 304028 162687
rect 303986 160848 304042 160857
rect 303986 160783 304042 160792
rect 309796 160750 309824 340954
rect 309888 275369 309916 375799
rect 311176 341154 311204 389030
rect 312556 386345 312584 390102
rect 314856 387666 314884 390116
rect 314844 387660 314896 387666
rect 314844 387602 314896 387608
rect 315304 387660 315356 387666
rect 315304 387602 315356 387608
rect 312542 386336 312598 386345
rect 312542 386271 312598 386280
rect 311438 365664 311494 365673
rect 311438 365599 311494 365608
rect 311256 350600 311308 350606
rect 311256 350542 311308 350548
rect 311164 341148 311216 341154
rect 311164 341090 311216 341096
rect 309968 339584 310020 339590
rect 309968 339526 310020 339532
rect 309874 275360 309930 275369
rect 309874 275295 309930 275304
rect 309980 251190 310008 339526
rect 310426 337376 310482 337385
rect 310426 337311 310482 337320
rect 310440 330857 310468 337311
rect 310426 330848 310482 330857
rect 310426 330783 310482 330792
rect 309968 251184 310020 251190
rect 309968 251126 310020 251132
rect 310518 175264 310574 175273
rect 310518 175199 310574 175208
rect 310532 171134 310560 175199
rect 310440 171106 310560 171134
rect 310440 169833 310468 171106
rect 310426 169824 310482 169833
rect 310426 169759 310482 169768
rect 309784 160744 309836 160750
rect 309784 160686 309836 160692
rect 298742 160304 298798 160313
rect 298742 160239 298798 160248
rect 311176 149734 311204 341090
rect 311268 201414 311296 350542
rect 311348 342372 311400 342378
rect 311348 342314 311400 342320
rect 311360 226234 311388 342314
rect 311452 279721 311480 365599
rect 312556 348430 312584 386271
rect 313924 383716 313976 383722
rect 313924 383658 313976 383664
rect 312544 348424 312596 348430
rect 312544 348366 312596 348372
rect 312556 302841 312584 348366
rect 312542 302832 312598 302841
rect 312542 302767 312598 302776
rect 311438 279712 311494 279721
rect 311438 279647 311494 279656
rect 311348 226228 311400 226234
rect 311348 226170 311400 226176
rect 313936 204270 313964 383658
rect 314198 367976 314254 367985
rect 314198 367911 314254 367920
rect 314108 346520 314160 346526
rect 314108 346462 314160 346468
rect 314016 343800 314068 343806
rect 314016 343742 314068 343748
rect 314028 209778 314056 343742
rect 314120 231810 314148 346462
rect 314212 256873 314240 367911
rect 315316 340950 315344 387602
rect 315394 373552 315450 373561
rect 315394 373487 315450 373496
rect 315304 340944 315356 340950
rect 315304 340886 315356 340892
rect 314198 256864 314254 256873
rect 314198 256799 314254 256808
rect 314108 231804 314160 231810
rect 314108 231746 314160 231752
rect 314660 218068 314712 218074
rect 314660 218010 314712 218016
rect 314672 211818 314700 218010
rect 314660 211812 314712 211818
rect 314660 211754 314712 211760
rect 314016 209772 314068 209778
rect 314016 209714 314068 209720
rect 313924 204264 313976 204270
rect 313924 204206 313976 204212
rect 311256 201408 311308 201414
rect 311256 201350 311308 201356
rect 315316 169250 315344 340886
rect 315408 202473 315436 373487
rect 316604 364334 316632 390215
rect 321834 390144 321890 390153
rect 318076 390102 318366 390130
rect 319732 390102 320114 390130
rect 318076 388929 318104 390102
rect 318062 388920 318118 388929
rect 319732 388890 319760 390102
rect 321834 390079 321890 390088
rect 318062 388855 318118 388864
rect 319720 388884 319772 388890
rect 316604 364306 316724 364334
rect 315486 350160 315542 350169
rect 315486 350095 315542 350104
rect 315500 291689 315528 350095
rect 316696 344078 316724 364306
rect 318076 350674 318104 388855
rect 319720 388826 319772 388832
rect 318154 384568 318210 384577
rect 318154 384503 318210 384512
rect 318064 350668 318116 350674
rect 318064 350610 318116 350616
rect 316684 344072 316736 344078
rect 316684 344014 316736 344020
rect 315580 298104 315632 298110
rect 315580 298046 315632 298052
rect 315486 291680 315542 291689
rect 315486 291615 315542 291624
rect 315592 275330 315620 298046
rect 315580 275324 315632 275330
rect 315580 275266 315632 275272
rect 315394 202464 315450 202473
rect 315394 202399 315450 202408
rect 315394 188456 315450 188465
rect 315394 188391 315450 188400
rect 315408 175409 315436 188391
rect 315394 175400 315450 175409
rect 315394 175335 315450 175344
rect 315304 169244 315356 169250
rect 315304 169186 315356 169192
rect 311164 149728 311216 149734
rect 311164 149670 311216 149676
rect 316696 148345 316724 344014
rect 316774 198792 316830 198801
rect 316774 198727 316830 198736
rect 316788 188465 316816 198727
rect 316774 188456 316830 188465
rect 316774 188391 316830 188400
rect 318076 148481 318104 350610
rect 318168 242729 318196 384503
rect 319732 373994 319760 388826
rect 321098 382256 321154 382265
rect 321098 382191 321154 382200
rect 320914 380896 320970 380905
rect 320914 380831 320970 380840
rect 319456 373966 319760 373994
rect 318246 361584 318302 361593
rect 318246 361519 318302 361528
rect 318260 282849 318288 361519
rect 319456 343942 319484 373966
rect 319626 368248 319682 368257
rect 319626 368183 319682 368192
rect 319444 343936 319496 343942
rect 319444 343878 319496 343884
rect 318246 282840 318302 282849
rect 318246 282775 318302 282784
rect 318248 275324 318300 275330
rect 318248 275266 318300 275272
rect 318260 260846 318288 275266
rect 318248 260840 318300 260846
rect 318248 260782 318300 260788
rect 318154 242720 318210 242729
rect 318154 242655 318210 242664
rect 318154 208584 318210 208593
rect 318154 208519 318210 208528
rect 318168 196081 318196 208519
rect 318338 208448 318394 208457
rect 318338 208383 318394 208392
rect 318352 198801 318380 208383
rect 318338 198792 318394 198801
rect 318338 198727 318394 198736
rect 318154 196072 318210 196081
rect 318154 196007 318210 196016
rect 318156 151836 318208 151842
rect 318156 151778 318208 151784
rect 318062 148472 318118 148481
rect 318062 148407 318118 148416
rect 316682 148336 316738 148345
rect 316682 148271 316738 148280
rect 297362 147384 297418 147393
rect 297362 147319 297418 147328
rect 295614 146976 295670 146985
rect 295614 146911 295670 146920
rect 295982 146976 296038 146985
rect 295982 146911 296038 146920
rect 295430 120592 295486 120601
rect 295430 120527 295486 120536
rect 295996 115938 296024 146911
rect 295984 115932 296036 115938
rect 295984 115874 296036 115880
rect 297376 115870 297404 147319
rect 318168 119678 318196 151778
rect 319456 148374 319484 343878
rect 319536 343868 319588 343874
rect 319536 343810 319588 343816
rect 319548 244186 319576 343810
rect 319640 280809 319668 368183
rect 320824 342304 320876 342310
rect 320824 342246 320876 342252
rect 319626 280800 319682 280809
rect 319626 280735 319682 280744
rect 319626 255368 319682 255377
rect 319626 255303 319682 255312
rect 319536 244180 319588 244186
rect 319536 244122 319588 244128
rect 319640 208457 319668 255303
rect 319720 250504 319772 250510
rect 319720 250446 319772 250452
rect 319732 212430 319760 250446
rect 320546 212528 320602 212537
rect 320546 212463 320602 212472
rect 319720 212424 319772 212430
rect 319720 212366 319772 212372
rect 320560 208593 320588 212463
rect 320836 211138 320864 342246
rect 320928 273193 320956 380831
rect 321008 341352 321060 341358
rect 321008 341294 321060 341300
rect 320914 273184 320970 273193
rect 320914 273119 320970 273128
rect 320914 263664 320970 263673
rect 320914 263599 320970 263608
rect 320928 255377 320956 263599
rect 320914 255368 320970 255377
rect 320914 255303 320970 255312
rect 321020 245614 321048 341294
rect 321112 302569 321140 382191
rect 321848 345014 321876 390079
rect 322386 386200 322442 386209
rect 322386 386135 322442 386144
rect 322296 347812 322348 347818
rect 322296 347754 322348 347760
rect 321848 344986 322244 345014
rect 322216 343738 322244 344986
rect 322204 343732 322256 343738
rect 322204 343674 322256 343680
rect 321098 302560 321154 302569
rect 321098 302495 321154 302504
rect 321008 245608 321060 245614
rect 321008 245550 321060 245556
rect 321928 212424 321980 212430
rect 321928 212366 321980 212372
rect 320824 211132 320876 211138
rect 320824 211074 320876 211080
rect 320546 208584 320602 208593
rect 320546 208519 320602 208528
rect 319626 208448 319682 208457
rect 319626 208383 319682 208392
rect 321940 204202 321968 212366
rect 321928 204196 321980 204202
rect 321928 204138 321980 204144
rect 320822 190768 320878 190777
rect 320822 190703 320878 190712
rect 319444 148368 319496 148374
rect 319444 148310 319496 148316
rect 318156 119672 318208 119678
rect 318156 119614 318208 119620
rect 297364 115864 297416 115870
rect 297364 115806 297416 115812
rect 294142 113792 294198 113801
rect 294142 113727 294198 113736
rect 320836 97889 320864 190703
rect 322216 148442 322244 343674
rect 322308 247042 322336 347754
rect 322400 288425 322428 386135
rect 323596 341426 323624 390351
rect 325516 390312 325568 390318
rect 325516 390254 325568 390260
rect 325528 390130 325556 390254
rect 343088 390176 343140 390182
rect 325358 390116 325556 390130
rect 325344 390102 325556 390116
rect 323674 366616 323730 366625
rect 323674 366551 323730 366560
rect 323584 341420 323636 341426
rect 323584 341362 323636 341368
rect 322386 288416 322442 288425
rect 322386 288351 322442 288360
rect 322296 247036 322348 247042
rect 322296 246978 322348 246984
rect 322294 230480 322350 230489
rect 322294 230415 322350 230424
rect 322308 212537 322336 230415
rect 322294 212528 322350 212537
rect 322294 212463 322350 212472
rect 322388 211812 322440 211818
rect 322388 211754 322440 211760
rect 322400 202162 322428 211754
rect 322388 202156 322440 202162
rect 322388 202098 322440 202104
rect 323596 148617 323624 341362
rect 323688 257961 323716 366551
rect 325344 354674 325372 390102
rect 326344 389836 326396 389842
rect 326344 389778 326396 389784
rect 324976 354646 325372 354674
rect 323766 340096 323822 340105
rect 323766 340031 323822 340040
rect 323780 303521 323808 340031
rect 324976 338774 325004 354646
rect 325056 346452 325108 346458
rect 325056 346394 325108 346400
rect 324964 338768 325016 338774
rect 324964 338710 325016 338716
rect 323766 303512 323822 303521
rect 323766 303447 323822 303456
rect 323768 260840 323820 260846
rect 323768 260782 323820 260788
rect 323674 257952 323730 257961
rect 323674 257887 323730 257896
rect 323674 252240 323730 252249
rect 323674 252175 323730 252184
rect 323688 230489 323716 252175
rect 323780 244254 323808 260782
rect 323768 244248 323820 244254
rect 323768 244190 323820 244196
rect 323674 230480 323730 230489
rect 323674 230415 323730 230424
rect 324976 162178 325004 338710
rect 325068 262206 325096 346394
rect 326356 330546 326384 389778
rect 327092 387462 327120 390116
rect 327080 387456 327132 387462
rect 327080 387398 327132 387404
rect 328840 387394 328868 390116
rect 328828 387388 328880 387394
rect 328828 387330 328880 387336
rect 330588 387326 330616 390116
rect 330576 387320 330628 387326
rect 330576 387262 330628 387268
rect 332336 387258 332364 390116
rect 332324 387252 332376 387258
rect 332324 387194 332376 387200
rect 334084 387190 334112 390116
rect 334072 387184 334124 387190
rect 334072 387126 334124 387132
rect 335832 387122 335860 390116
rect 337580 387734 337608 390116
rect 339328 387802 339356 390116
rect 341090 390102 341564 390130
rect 342838 390124 343088 390130
rect 342838 390118 343140 390124
rect 342838 390116 343128 390118
rect 339316 387796 339368 387802
rect 339316 387738 339368 387744
rect 337568 387728 337620 387734
rect 337568 387670 337620 387676
rect 339328 387122 339356 387738
rect 341536 387258 341564 390102
rect 342824 390102 343128 390116
rect 341524 387252 341576 387258
rect 341524 387194 341576 387200
rect 335820 387116 335872 387122
rect 335820 387058 335872 387064
rect 339316 387116 339368 387122
rect 339316 387058 339368 387064
rect 341536 371890 341564 387194
rect 341524 371884 341576 371890
rect 341524 371826 341576 371832
rect 341524 366648 341576 366654
rect 341524 366590 341576 366596
rect 333244 366580 333296 366586
rect 333244 366522 333296 366528
rect 329102 353152 329158 353161
rect 329102 353087 329158 353096
rect 327814 348528 327870 348537
rect 327814 348463 327870 348472
rect 327724 345160 327776 345166
rect 327724 345102 327776 345108
rect 326344 330540 326396 330546
rect 326344 330482 326396 330488
rect 325882 273048 325938 273057
rect 325804 273006 325882 273034
rect 325804 270494 325832 273006
rect 325882 272983 325938 272992
rect 325160 270466 325832 270494
rect 325160 263673 325188 270466
rect 325146 263664 325202 263673
rect 325146 263599 325202 263608
rect 325056 262200 325108 262206
rect 325056 262142 325108 262148
rect 326986 253872 327042 253881
rect 326986 253807 327042 253816
rect 327000 252249 327028 253807
rect 326986 252240 327042 252249
rect 326986 252175 327042 252184
rect 326344 244248 326396 244254
rect 326344 244190 326396 244196
rect 326356 202842 326384 244190
rect 327736 216646 327764 345102
rect 327828 308009 327856 348463
rect 327814 308000 327870 308009
rect 327814 307935 327870 307944
rect 327814 288280 327870 288289
rect 327814 288215 327870 288224
rect 327828 273057 327856 288215
rect 329116 277545 329144 353087
rect 331862 339552 331918 339561
rect 331862 339487 331918 339496
rect 329196 330540 329248 330546
rect 329196 330482 329248 330488
rect 329208 307766 329236 330482
rect 329196 307760 329248 307766
rect 329196 307702 329248 307708
rect 329930 291136 329986 291145
rect 329930 291071 329986 291080
rect 329944 288289 329972 291071
rect 329930 288280 329986 288289
rect 329930 288215 329986 288224
rect 330482 282296 330538 282305
rect 330482 282231 330538 282240
rect 329102 277536 329158 277545
rect 329102 277471 329158 277480
rect 330496 274689 330524 282231
rect 329102 274680 329158 274689
rect 329102 274615 329158 274624
rect 330482 274680 330538 274689
rect 330482 274615 330538 274624
rect 327814 273048 327870 273057
rect 327814 272983 327870 272992
rect 329116 253881 329144 274615
rect 329102 253872 329158 253881
rect 329102 253807 329158 253816
rect 327724 216640 327776 216646
rect 327724 216582 327776 216588
rect 326436 204196 326488 204202
rect 326436 204138 326488 204144
rect 326344 202836 326396 202842
rect 326344 202778 326396 202784
rect 326448 198762 326476 204138
rect 330484 202836 330536 202842
rect 330484 202778 330536 202784
rect 326436 198756 326488 198762
rect 326436 198698 326488 198704
rect 329104 198756 329156 198762
rect 329104 198698 329156 198704
rect 329116 189106 329144 198698
rect 329104 189100 329156 189106
rect 329104 189042 329156 189048
rect 330496 184210 330524 202778
rect 330484 184204 330536 184210
rect 330484 184146 330536 184152
rect 324964 162172 325016 162178
rect 324964 162114 325016 162120
rect 323582 148608 323638 148617
rect 323582 148543 323638 148552
rect 322204 148436 322256 148442
rect 322204 148378 322256 148384
rect 320822 97880 320878 97889
rect 320822 97815 320878 97824
rect 304354 86184 304410 86193
rect 304354 86119 304410 86128
rect 297270 32600 297326 32609
rect 297270 32535 297326 32544
rect 292580 4140 292632 4146
rect 292580 4082 292632 4088
rect 293682 3632 293738 3641
rect 293682 3567 293738 3576
rect 293696 480 293724 3567
rect 297284 480 297312 32535
rect 300766 3496 300822 3505
rect 300766 3431 300822 3440
rect 300780 480 300808 3431
rect 304368 480 304396 86119
rect 322110 85776 322166 85785
rect 322110 85711 322166 85720
rect 311438 82104 311494 82113
rect 311438 82039 311494 82048
rect 307114 59936 307170 59945
rect 307114 59871 307170 59880
rect 307128 53281 307156 59871
rect 307114 53272 307170 53281
rect 307114 53207 307170 53216
rect 307942 53136 307998 53145
rect 307942 53071 307998 53080
rect 307956 480 307984 53071
rect 311452 480 311480 82039
rect 318522 80744 318578 80753
rect 318522 80679 318578 80688
rect 315026 51776 315082 51785
rect 315026 51711 315082 51720
rect 315040 480 315068 51711
rect 318536 480 318564 80679
rect 322124 480 322152 85711
rect 329194 79384 329250 79393
rect 329194 79319 329250 79328
rect 324962 58576 325018 58585
rect 324962 58511 325018 58520
rect 324976 7721 325004 58511
rect 324962 7712 325018 7721
rect 324962 7647 325018 7656
rect 325606 7576 325662 7585
rect 325606 7511 325662 7520
rect 325620 480 325648 7511
rect 329208 480 329236 79319
rect 331876 6866 331904 339487
rect 331956 307760 332008 307766
rect 331956 307702 332008 307708
rect 331968 295390 331996 307702
rect 332046 300792 332102 300801
rect 332046 300727 332102 300736
rect 331956 295384 332008 295390
rect 331956 295326 332008 295332
rect 331954 292632 332010 292641
rect 331954 292567 332010 292576
rect 331968 282305 331996 292567
rect 332060 291145 332088 300727
rect 332046 291136 332102 291145
rect 332046 291071 332102 291080
rect 331954 282296 332010 282305
rect 331954 282231 332010 282240
rect 332508 202156 332560 202162
rect 332508 202098 332560 202104
rect 332520 198014 332548 202098
rect 332508 198008 332560 198014
rect 332508 197950 332560 197956
rect 333256 177682 333284 366522
rect 333428 364200 333480 364206
rect 333428 364142 333480 364148
rect 333336 363928 333388 363934
rect 333336 363870 333388 363876
rect 333244 177676 333296 177682
rect 333244 177618 333296 177624
rect 333348 177410 333376 363870
rect 333336 177404 333388 177410
rect 333336 177346 333388 177352
rect 333440 177274 333468 364142
rect 336004 364132 336056 364138
rect 336004 364074 336056 364080
rect 334624 345092 334676 345098
rect 334624 345034 334676 345040
rect 333518 343088 333574 343097
rect 333518 343023 333574 343032
rect 333532 300801 333560 343023
rect 333518 300792 333574 300801
rect 333518 300727 333574 300736
rect 334636 206922 334664 345034
rect 334714 342952 334770 342961
rect 334714 342887 334770 342896
rect 334728 305833 334756 342887
rect 334806 306504 334862 306513
rect 334806 306439 334862 306448
rect 334714 305824 334770 305833
rect 334714 305759 334770 305768
rect 334820 292641 334848 306439
rect 334806 292632 334862 292641
rect 334806 292567 334862 292576
rect 334624 206916 334676 206922
rect 334624 206858 334676 206864
rect 336016 178498 336044 364074
rect 338764 364064 338816 364070
rect 338764 364006 338816 364012
rect 336372 361412 336424 361418
rect 336372 361354 336424 361360
rect 336188 361344 336240 361350
rect 336188 361286 336240 361292
rect 336096 361140 336148 361146
rect 336096 361082 336148 361088
rect 336004 178492 336056 178498
rect 336004 178434 336056 178440
rect 336108 177857 336136 361082
rect 336094 177848 336150 177857
rect 336094 177783 336150 177792
rect 333428 177268 333480 177274
rect 333428 177210 333480 177216
rect 336200 177138 336228 361286
rect 336280 361276 336332 361282
rect 336280 361218 336332 361224
rect 336292 177206 336320 361218
rect 336384 180441 336412 361354
rect 336464 350260 336516 350266
rect 336464 350202 336516 350208
rect 336370 180432 336426 180441
rect 336370 180367 336426 180376
rect 336476 180334 336504 350202
rect 337382 347168 337438 347177
rect 337382 347103 337438 347112
rect 336556 341216 336608 341222
rect 336556 341158 336608 341164
rect 336568 222086 336596 341158
rect 336646 338872 336702 338881
rect 336646 338807 336702 338816
rect 336660 327593 336688 338807
rect 336646 327584 336702 327593
rect 336646 327519 336702 327528
rect 337396 306513 337424 347103
rect 337382 306504 337438 306513
rect 337382 306439 337438 306448
rect 337384 295384 337436 295390
rect 337384 295326 337436 295332
rect 337396 285734 337424 295326
rect 337384 285728 337436 285734
rect 337384 285670 337436 285676
rect 336556 222080 336608 222086
rect 336556 222022 336608 222028
rect 338028 189100 338080 189106
rect 338028 189042 338080 189048
rect 338040 181490 338068 189042
rect 338028 181484 338080 181490
rect 338028 181426 338080 181432
rect 336464 180328 336516 180334
rect 336464 180270 336516 180276
rect 338776 180198 338804 364006
rect 338856 361208 338908 361214
rect 338856 361150 338908 361156
rect 338764 180192 338816 180198
rect 338764 180134 338816 180140
rect 338868 178838 338896 361150
rect 338948 358284 339000 358290
rect 338948 358226 339000 358232
rect 338960 179081 338988 358226
rect 339040 350124 339092 350130
rect 339040 350066 339092 350072
rect 339052 180266 339080 350066
rect 339406 345128 339462 345137
rect 339406 345063 339462 345072
rect 339420 343097 339448 345063
rect 339406 343088 339462 343097
rect 339406 343023 339462 343032
rect 339224 342440 339276 342446
rect 339224 342382 339276 342388
rect 339130 302832 339186 302841
rect 339130 302767 339186 302776
rect 339040 180260 339092 180266
rect 339040 180202 339092 180208
rect 338946 179072 339002 179081
rect 338946 179007 339002 179016
rect 338856 178832 338908 178838
rect 338856 178774 338908 178780
rect 336280 177200 336332 177206
rect 336280 177142 336332 177148
rect 336188 177132 336240 177138
rect 336188 177074 336240 177080
rect 339144 151201 339172 302767
rect 339236 288386 339264 342382
rect 339224 288380 339276 288386
rect 339224 288322 339276 288328
rect 341536 179178 341564 366590
rect 341708 364268 341760 364274
rect 341708 364210 341760 364216
rect 341614 363624 341670 363633
rect 341614 363559 341670 363568
rect 341524 179172 341576 179178
rect 341524 179114 341576 179120
rect 341628 176633 341656 363559
rect 341720 179042 341748 364210
rect 341892 355768 341944 355774
rect 341892 355710 341944 355716
rect 341800 355700 341852 355706
rect 341800 355642 341852 355648
rect 341812 179314 341840 355642
rect 341904 179353 341932 355710
rect 342824 340814 342852 390102
rect 344572 387802 344600 390116
rect 346228 390114 346334 390130
rect 346216 390108 346334 390114
rect 346268 390102 346334 390108
rect 348082 390102 348464 390130
rect 349830 390102 350120 390130
rect 346216 390050 346268 390056
rect 343640 387796 343692 387802
rect 343640 387738 343692 387744
rect 344560 387796 344612 387802
rect 344560 387738 344612 387744
rect 343652 387530 343680 387738
rect 343640 387524 343692 387530
rect 343640 387466 343692 387472
rect 346228 383654 346256 390050
rect 346308 389020 346360 389026
rect 346308 388962 346360 388968
rect 346320 387977 346348 388962
rect 346306 387968 346362 387977
rect 346306 387903 346362 387912
rect 348436 387530 348464 390102
rect 349804 388952 349856 388958
rect 349804 388894 349856 388900
rect 349816 388113 349844 388894
rect 349802 388104 349858 388113
rect 349802 388039 349858 388048
rect 348424 387524 348476 387530
rect 348424 387466 348476 387472
rect 346228 383626 346348 383654
rect 344376 355632 344428 355638
rect 344376 355574 344428 355580
rect 344284 355496 344336 355502
rect 344284 355438 344336 355444
rect 342904 341284 342956 341290
rect 342904 341226 342956 341232
rect 342812 340808 342864 340814
rect 342812 340750 342864 340756
rect 342260 285728 342312 285734
rect 342260 285670 342312 285676
rect 342272 279478 342300 285670
rect 342916 282878 342944 341226
rect 342904 282872 342956 282878
rect 342904 282814 342956 282820
rect 342260 279472 342312 279478
rect 342260 279414 342312 279420
rect 341890 179344 341946 179353
rect 341800 179308 341852 179314
rect 341890 179279 341946 179288
rect 341800 179250 341852 179256
rect 341708 179036 341760 179042
rect 341708 178978 341760 178984
rect 344296 178770 344324 355438
rect 344388 178974 344416 355574
rect 344468 350192 344520 350198
rect 344468 350134 344520 350140
rect 344480 180402 344508 350134
rect 346214 349888 346270 349897
rect 346214 349823 346270 349832
rect 344560 347200 344612 347206
rect 344560 347142 344612 347148
rect 344572 180470 344600 347142
rect 346228 345137 346256 349823
rect 346214 345128 346270 345137
rect 346214 345063 346270 345072
rect 345662 344312 345718 344321
rect 345662 344247 345718 344256
rect 345676 309097 345704 344247
rect 346320 340202 346348 383626
rect 347044 363996 347096 364002
rect 347044 363938 347096 363944
rect 346308 340196 346360 340202
rect 346308 340138 346360 340144
rect 345662 309088 345718 309097
rect 345662 309023 345718 309032
rect 344560 180464 344612 180470
rect 344560 180406 344612 180412
rect 344468 180396 344520 180402
rect 344468 180338 344520 180344
rect 344376 178968 344428 178974
rect 344376 178910 344428 178916
rect 344284 178764 344336 178770
rect 344284 178706 344336 178712
rect 341614 176624 341670 176633
rect 347056 176594 347084 363938
rect 347136 363860 347188 363866
rect 347136 363802 347188 363808
rect 347148 180606 347176 363802
rect 347228 361072 347280 361078
rect 347228 361014 347280 361020
rect 347136 180600 347188 180606
rect 347136 180542 347188 180548
rect 347240 178022 347268 361014
rect 347320 358216 347372 358222
rect 347320 358158 347372 358164
rect 347228 178016 347280 178022
rect 347228 177958 347280 177964
rect 347332 176662 347360 358158
rect 347504 353048 347556 353054
rect 347504 352990 347556 352996
rect 347412 352980 347464 352986
rect 347412 352922 347464 352928
rect 347424 179110 347452 352922
rect 347516 179246 347544 352990
rect 347594 352608 347650 352617
rect 347594 352543 347650 352552
rect 347608 180305 347636 352543
rect 348436 340882 348464 387466
rect 350092 387025 350120 390102
rect 351564 387297 351592 390116
rect 353312 387433 353340 390116
rect 353298 387424 353354 387433
rect 353298 387359 353354 387368
rect 351550 387288 351606 387297
rect 351550 387223 351606 387232
rect 350078 387016 350134 387025
rect 350078 386951 350134 386960
rect 353942 387016 353998 387025
rect 353942 386951 353998 386960
rect 350446 360768 350502 360777
rect 350446 360703 350502 360712
rect 349896 358148 349948 358154
rect 349896 358090 349948 358096
rect 349804 358080 349856 358086
rect 349804 358022 349856 358028
rect 348424 340876 348476 340882
rect 348424 340818 348476 340824
rect 347594 180296 347650 180305
rect 347594 180231 347650 180240
rect 347504 179240 347556 179246
rect 347504 179182 347556 179188
rect 347412 179104 347464 179110
rect 347412 179046 347464 179052
rect 349816 177585 349844 358022
rect 349908 178945 349936 358090
rect 350080 353116 350132 353122
rect 350080 353058 350132 353064
rect 349988 352776 350040 352782
rect 349988 352718 350040 352724
rect 349894 178936 349950 178945
rect 349894 178871 349950 178880
rect 350000 177750 350028 352718
rect 350092 177818 350120 353058
rect 350264 347268 350316 347274
rect 350264 347210 350316 347216
rect 350172 347132 350224 347138
rect 350172 347074 350224 347080
rect 350184 180674 350212 347074
rect 350172 180668 350224 180674
rect 350172 180610 350224 180616
rect 350276 180130 350304 347210
rect 350356 342916 350408 342922
rect 350356 342858 350408 342864
rect 350368 180538 350396 342858
rect 350460 310185 350488 360703
rect 352656 352912 352708 352918
rect 352656 352854 352708 352860
rect 352564 352708 352616 352714
rect 352564 352650 352616 352656
rect 351182 348392 351238 348401
rect 351182 348327 351238 348336
rect 351196 314537 351224 348327
rect 351182 314528 351238 314537
rect 351182 314463 351238 314472
rect 350446 310176 350502 310185
rect 350446 310111 350502 310120
rect 351184 279472 351236 279478
rect 351184 279414 351236 279420
rect 351196 189786 351224 279414
rect 351184 189780 351236 189786
rect 351184 189722 351236 189728
rect 351184 184204 351236 184210
rect 351184 184146 351236 184152
rect 350356 180532 350408 180538
rect 350356 180474 350408 180480
rect 350264 180124 350316 180130
rect 350264 180066 350316 180072
rect 351196 179926 351224 184146
rect 351184 179920 351236 179926
rect 351184 179862 351236 179868
rect 350080 177812 350132 177818
rect 350080 177754 350132 177760
rect 349988 177744 350040 177750
rect 349988 177686 350040 177692
rect 349802 177576 349858 177585
rect 352576 177546 352604 352650
rect 352668 177614 352696 352854
rect 352748 352844 352800 352850
rect 352748 352786 352800 352792
rect 352760 178906 352788 352786
rect 352840 350056 352892 350062
rect 352840 349998 352892 350004
rect 352748 178900 352800 178906
rect 352748 178842 352800 178848
rect 352656 177608 352708 177614
rect 352656 177550 352708 177556
rect 349802 177511 349858 177520
rect 352564 177540 352616 177546
rect 352564 177482 352616 177488
rect 352852 177478 352880 349998
rect 353298 349752 353354 349761
rect 353298 349687 353354 349696
rect 353312 347177 353340 349687
rect 353298 347168 353354 347177
rect 353298 347103 353354 347112
rect 352932 198008 352984 198014
rect 352932 197950 352984 197956
rect 352944 184210 352972 197950
rect 352932 184204 352984 184210
rect 352932 184146 352984 184152
rect 352840 177472 352892 177478
rect 352840 177414 352892 177420
rect 347320 176656 347372 176662
rect 347320 176598 347372 176604
rect 341614 176559 341670 176568
rect 347044 176588 347096 176594
rect 347044 176530 347096 176536
rect 349988 169176 350040 169182
rect 349988 169118 350040 169124
rect 349804 169108 349856 169114
rect 349804 169050 349856 169056
rect 339130 151192 339186 151201
rect 339130 151127 339186 151136
rect 349816 118454 349844 169050
rect 349896 169040 349948 169046
rect 349896 168982 349948 168988
rect 349804 118448 349856 118454
rect 349804 118390 349856 118396
rect 349908 118250 349936 168982
rect 350000 118318 350028 169118
rect 353956 147665 353984 386951
rect 355060 340338 355088 390116
rect 355968 387048 356020 387054
rect 355968 386990 356020 386996
rect 355980 385098 356008 386990
rect 355888 385070 356008 385098
rect 355888 383654 355916 385070
rect 355968 384940 356020 384946
rect 355968 384882 356020 384888
rect 355980 384033 356008 384882
rect 355966 384024 356022 384033
rect 355966 383959 356022 383968
rect 355888 383626 356008 383654
rect 355324 361004 355376 361010
rect 355324 360946 355376 360952
rect 355048 340332 355100 340338
rect 355048 340274 355100 340280
rect 355336 180062 355364 360946
rect 355416 355428 355468 355434
rect 355416 355370 355468 355376
rect 355324 180056 355376 180062
rect 355324 179998 355376 180004
rect 355428 179382 355456 355370
rect 355508 352640 355560 352646
rect 355508 352582 355560 352588
rect 355416 179376 355468 179382
rect 355416 179318 355468 179324
rect 355520 177721 355548 352582
rect 355600 352572 355652 352578
rect 355600 352514 355652 352520
rect 355612 177954 355640 352514
rect 355692 244928 355744 244934
rect 355692 244870 355744 244876
rect 355704 181801 355732 244870
rect 355690 181792 355746 181801
rect 355690 181727 355746 181736
rect 355704 180794 355732 181727
rect 355704 180766 355916 180794
rect 355600 177948 355652 177954
rect 355600 177890 355652 177896
rect 355506 177712 355562 177721
rect 355506 177647 355562 177656
rect 355888 173233 355916 180766
rect 355874 173224 355930 173233
rect 355874 173159 355930 173168
rect 355980 151814 356008 383626
rect 356704 366580 356756 366586
rect 356704 366522 356756 366528
rect 356716 343126 356744 366522
rect 356704 343120 356756 343126
rect 356704 343062 356756 343068
rect 356808 342242 356836 390116
rect 357346 387288 357402 387297
rect 357268 387246 357346 387274
rect 357268 383654 357296 387246
rect 357346 387223 357402 387232
rect 357348 384872 357400 384878
rect 357348 384814 357400 384820
rect 357360 383897 357388 384814
rect 357346 383888 357402 383897
rect 357346 383823 357402 383832
rect 357268 383626 357388 383654
rect 357254 347848 357310 347857
rect 357254 347783 357310 347792
rect 356796 342236 356848 342242
rect 356796 342178 356848 342184
rect 357268 299441 357296 347783
rect 357360 299538 357388 383626
rect 358266 373144 358322 373153
rect 358266 373079 358322 373088
rect 358084 366512 358136 366518
rect 358084 366454 358136 366460
rect 357348 299532 357400 299538
rect 357348 299474 357400 299480
rect 357254 299432 357310 299441
rect 357310 299390 357480 299418
rect 357254 299367 357310 299376
rect 357348 299328 357400 299334
rect 357348 299270 357400 299276
rect 355888 151786 356008 151814
rect 352562 147656 352618 147665
rect 352562 147591 352618 147600
rect 353942 147656 353998 147665
rect 353942 147591 353998 147600
rect 350078 147112 350134 147121
rect 350078 147047 350134 147056
rect 350092 120018 350120 147047
rect 350080 120012 350132 120018
rect 350080 119954 350132 119960
rect 349988 118312 350040 118318
rect 349988 118254 350040 118260
rect 349896 118244 349948 118250
rect 349896 118186 349948 118192
rect 352576 115569 352604 147591
rect 355416 146804 355468 146810
rect 355416 146746 355468 146752
rect 352656 146736 352708 146742
rect 352656 146678 352708 146684
rect 355322 146704 355378 146713
rect 352668 116958 352696 146678
rect 355322 146639 355378 146648
rect 352746 146568 352802 146577
rect 352746 146503 352802 146512
rect 352656 116952 352708 116958
rect 352656 116894 352708 116900
rect 352760 115705 352788 146503
rect 352930 146432 352986 146441
rect 352930 146367 352986 146376
rect 352746 115696 352802 115705
rect 352746 115631 352802 115640
rect 352562 115560 352618 115569
rect 352562 115495 352618 115504
rect 352944 115433 352972 146367
rect 355336 115841 355364 146639
rect 355428 117094 355456 146746
rect 355600 146464 355652 146470
rect 355600 146406 355652 146412
rect 355506 144392 355562 144401
rect 355506 144327 355562 144336
rect 355416 117088 355468 117094
rect 355520 117065 355548 144327
rect 355612 120630 355640 146406
rect 355888 146334 355916 151786
rect 355966 147384 356022 147393
rect 355966 147319 356022 147328
rect 355980 146946 356008 147319
rect 355968 146940 356020 146946
rect 355968 146882 356020 146888
rect 357360 146577 357388 299270
rect 357452 171134 357480 299390
rect 357532 288380 357584 288386
rect 357532 288322 357584 288328
rect 357544 287881 357572 288322
rect 357530 287872 357586 287881
rect 357530 287807 357586 287816
rect 357532 282872 357584 282878
rect 357532 282814 357584 282820
rect 357544 282305 357572 282814
rect 357530 282296 357586 282305
rect 357530 282231 357586 282240
rect 357532 277364 357584 277370
rect 357532 277306 357584 277312
rect 357544 276865 357572 277306
rect 357530 276856 357586 276865
rect 357530 276791 357586 276800
rect 357532 273216 357584 273222
rect 357532 273158 357584 273164
rect 357544 272649 357572 273158
rect 357530 272640 357586 272649
rect 357530 272575 357586 272584
rect 357532 271856 357584 271862
rect 357532 271798 357584 271804
rect 357544 271425 357572 271798
rect 357530 271416 357586 271425
rect 357530 271351 357586 271360
rect 357532 270496 357584 270502
rect 357532 270438 357584 270444
rect 357544 270201 357572 270438
rect 357530 270192 357586 270201
rect 357530 270127 357586 270136
rect 357532 262200 357584 262206
rect 357532 262142 357584 262148
rect 357544 261633 357572 262142
rect 357530 261624 357586 261633
rect 357530 261559 357586 261568
rect 357532 256692 357584 256698
rect 357532 256634 357584 256640
rect 357544 256193 357572 256634
rect 357530 256184 357586 256193
rect 357530 256119 357586 256128
rect 357532 255264 357584 255270
rect 357532 255206 357584 255212
rect 357544 254969 357572 255206
rect 357530 254960 357586 254969
rect 357530 254895 357586 254904
rect 357532 251184 357584 251190
rect 357532 251126 357584 251132
rect 357544 250753 357572 251126
rect 357530 250744 357586 250753
rect 357530 250679 357586 250688
rect 357532 247036 357584 247042
rect 357532 246978 357584 246984
rect 357544 246945 357572 246978
rect 357530 246936 357586 246945
rect 357530 246871 357586 246880
rect 357532 245608 357584 245614
rect 357532 245550 357584 245556
rect 357544 245177 357572 245550
rect 357530 245168 357586 245177
rect 357530 245103 357586 245112
rect 357532 244248 357584 244254
rect 357532 244190 357584 244196
rect 357544 243953 357572 244190
rect 357530 243944 357586 243953
rect 357530 243879 357586 243888
rect 357532 240100 357584 240106
rect 357532 240042 357584 240048
rect 357544 239737 357572 240042
rect 357530 239728 357586 239737
rect 357530 239663 357586 239672
rect 357532 235952 357584 235958
rect 357532 235894 357584 235900
rect 357544 235521 357572 235894
rect 357530 235512 357586 235521
rect 357530 235447 357586 235456
rect 357532 231804 357584 231810
rect 357532 231746 357584 231752
rect 357544 231305 357572 231746
rect 357530 231296 357586 231305
rect 357530 231231 357586 231240
rect 357716 226296 357768 226302
rect 357530 226264 357586 226273
rect 357716 226238 357768 226244
rect 357530 226199 357532 226208
rect 357584 226199 357586 226208
rect 357532 226170 357584 226176
rect 357728 225729 357756 226238
rect 357714 225720 357770 225729
rect 357714 225655 357770 225664
rect 357532 224936 357584 224942
rect 357532 224878 357584 224884
rect 357544 224505 357572 224878
rect 357530 224496 357586 224505
rect 357530 224431 357586 224440
rect 357532 223576 357584 223582
rect 357532 223518 357584 223524
rect 357544 223281 357572 223518
rect 357530 223272 357586 223281
rect 357530 223207 357586 223216
rect 357716 222148 357768 222154
rect 357716 222090 357768 222096
rect 357532 222080 357584 222086
rect 357530 222048 357532 222057
rect 357584 222048 357586 222057
rect 357530 221983 357586 221992
rect 357728 221513 357756 222090
rect 357714 221504 357770 221513
rect 357714 221439 357770 221448
rect 357532 218000 357584 218006
rect 357532 217942 357584 217948
rect 357544 217841 357572 217942
rect 357530 217832 357586 217841
rect 357530 217767 357586 217776
rect 357532 216640 357584 216646
rect 357530 216608 357532 216617
rect 357584 216608 357586 216617
rect 357530 216543 357586 216552
rect 357532 215280 357584 215286
rect 357532 215222 357584 215228
rect 357544 214849 357572 215222
rect 357530 214840 357586 214849
rect 357530 214775 357586 214784
rect 357532 212492 357584 212498
rect 357532 212434 357584 212440
rect 357544 212401 357572 212434
rect 357530 212392 357586 212401
rect 357530 212327 357586 212336
rect 357530 211168 357586 211177
rect 357530 211103 357532 211112
rect 357584 211103 357586 211112
rect 357532 211074 357584 211080
rect 357532 209772 357584 209778
rect 357532 209714 357584 209720
rect 357544 209409 357572 209714
rect 357530 209400 357586 209409
rect 357530 209335 357586 209344
rect 357532 208344 357584 208350
rect 357532 208286 357584 208292
rect 357544 208049 357572 208286
rect 357530 208040 357586 208049
rect 357530 207975 357586 207984
rect 357532 206984 357584 206990
rect 357532 206926 357584 206932
rect 357544 206825 357572 206926
rect 357530 206816 357586 206825
rect 357530 206751 357586 206760
rect 357532 206712 357584 206718
rect 357532 206654 357584 206660
rect 357544 206281 357572 206654
rect 357530 206272 357586 206281
rect 357530 206207 357586 206216
rect 357532 205624 357584 205630
rect 357532 205566 357584 205572
rect 357544 205057 357572 205566
rect 357530 205048 357586 205057
rect 357530 204983 357586 204992
rect 357532 204264 357584 204270
rect 357532 204206 357584 204212
rect 357544 203833 357572 204206
rect 357530 203824 357586 203833
rect 357530 203759 357586 203768
rect 357532 201476 357584 201482
rect 357532 201418 357584 201424
rect 357544 201385 357572 201418
rect 357530 201376 357586 201385
rect 357530 201311 357586 201320
rect 357532 201272 357584 201278
rect 357532 201214 357584 201220
rect 357544 200841 357572 201214
rect 357530 200832 357586 200841
rect 357530 200767 357586 200776
rect 357532 195968 357584 195974
rect 357530 195936 357532 195945
rect 357584 195936 357586 195945
rect 357530 195871 357586 195880
rect 358096 179994 358124 366454
rect 358176 347064 358228 347070
rect 358176 347006 358228 347012
rect 358084 179988 358136 179994
rect 358084 179930 358136 179936
rect 358188 177993 358216 347006
rect 358280 298761 358308 373079
rect 358360 367804 358412 367810
rect 358360 367746 358412 367752
rect 358372 343194 358400 367746
rect 358450 356008 358506 356017
rect 358450 355943 358506 355952
rect 358360 343188 358412 343194
rect 358360 343130 358412 343136
rect 358360 339448 358412 339454
rect 358360 339390 358412 339396
rect 358266 298752 358322 298761
rect 358266 298687 358322 298696
rect 358372 293865 358400 339390
rect 358464 325553 358492 355943
rect 358556 342990 358584 390116
rect 359648 388476 359700 388482
rect 359648 388418 359700 388424
rect 359660 387598 359688 388418
rect 359648 387592 359700 387598
rect 359648 387534 359700 387540
rect 359660 386753 359688 387534
rect 360014 387424 360070 387433
rect 360014 387359 360070 387368
rect 359740 387184 359792 387190
rect 359740 387126 359792 387132
rect 359830 387152 359886 387161
rect 359646 386744 359702 386753
rect 359646 386679 359702 386688
rect 359372 369164 359424 369170
rect 359372 369106 359424 369112
rect 358726 351928 358782 351937
rect 358726 351863 358782 351872
rect 358544 342984 358596 342990
rect 358544 342926 358596 342932
rect 358634 338736 358690 338745
rect 358634 338671 358690 338680
rect 358542 336016 358598 336025
rect 358542 335951 358598 335960
rect 358450 325544 358506 325553
rect 358450 325479 358506 325488
rect 358556 317257 358584 335951
rect 358648 323785 358676 338671
rect 358634 323776 358690 323785
rect 358634 323711 358690 323720
rect 358542 317248 358598 317257
rect 358542 317183 358598 317192
rect 358358 293856 358414 293865
rect 358358 293791 358414 293800
rect 358268 189780 358320 189786
rect 358268 189722 358320 189728
rect 358280 178702 358308 189722
rect 358636 181484 358688 181490
rect 358636 181426 358688 181432
rect 358268 178696 358320 178702
rect 358268 178638 358320 178644
rect 358648 178090 358676 181426
rect 358636 178084 358688 178090
rect 358636 178026 358688 178032
rect 358174 177984 358230 177993
rect 358174 177919 358230 177928
rect 358740 172553 358768 351863
rect 359384 343058 359412 369106
rect 359464 363792 359516 363798
rect 359464 363734 359516 363740
rect 359372 343052 359424 343058
rect 359372 342994 359424 343000
rect 359476 177342 359504 363734
rect 359556 360936 359608 360942
rect 359556 360878 359608 360884
rect 359568 180577 359596 360878
rect 359648 349988 359700 349994
rect 359648 349930 359700 349936
rect 359554 180568 359610 180577
rect 359554 180503 359610 180512
rect 359660 178022 359688 349930
rect 359752 340270 359780 387126
rect 359830 387087 359886 387096
rect 359844 347041 359872 387087
rect 360028 386617 360056 387359
rect 360200 387252 360252 387258
rect 360200 387194 360252 387200
rect 360108 387116 360160 387122
rect 360108 387058 360160 387064
rect 360014 386608 360070 386617
rect 360120 386578 360148 387058
rect 360014 386543 360070 386552
rect 360108 386572 360160 386578
rect 359924 351484 359976 351490
rect 359924 351426 359976 351432
rect 359830 347032 359886 347041
rect 359830 346967 359886 346976
rect 359740 340264 359792 340270
rect 359740 340206 359792 340212
rect 359740 184204 359792 184210
rect 359740 184146 359792 184152
rect 359752 178634 359780 184146
rect 359936 180169 359964 351426
rect 359922 180160 359978 180169
rect 359922 180095 359978 180104
rect 359740 178628 359792 178634
rect 359740 178570 359792 178576
rect 359648 178016 359700 178022
rect 359648 177958 359700 177964
rect 359464 177336 359516 177342
rect 359464 177278 359516 177284
rect 358726 172544 358782 172553
rect 358726 172479 358782 172488
rect 357452 171106 357572 171134
rect 357544 147121 357572 171106
rect 358740 161474 358768 172479
rect 360028 171737 360056 386543
rect 360108 386514 360160 386520
rect 360014 171728 360070 171737
rect 360014 171663 360070 171672
rect 360120 169318 360148 386514
rect 360212 386510 360240 387194
rect 360200 386504 360252 386510
rect 360198 386472 360200 386481
rect 360252 386472 360254 386481
rect 360198 386407 360254 386416
rect 360304 345030 360332 390116
rect 360476 389836 360528 389842
rect 360476 389778 360528 389784
rect 360384 387116 360436 387122
rect 360384 387058 360436 387064
rect 360396 346390 360424 387058
rect 360488 387054 360516 389778
rect 360476 387048 360528 387054
rect 360476 386990 360528 386996
rect 362052 386889 362080 390116
rect 363800 386889 363828 390116
rect 362038 386880 362094 386889
rect 362038 386815 362094 386824
rect 363786 386880 363842 386889
rect 363786 386815 363842 386824
rect 365548 359417 365576 390116
rect 367296 362817 367324 390116
rect 369044 384169 369072 390116
rect 369030 384160 369086 384169
rect 369030 384095 369086 384104
rect 370792 368121 370820 390116
rect 370778 368112 370834 368121
rect 370778 368047 370834 368056
rect 367282 362808 367338 362817
rect 367282 362743 367338 362752
rect 365534 359408 365590 359417
rect 365534 359343 365590 359352
rect 372540 355201 372568 390116
rect 372526 355192 372582 355201
rect 372526 355127 372582 355136
rect 374288 353705 374316 390116
rect 376036 377913 376064 390116
rect 376022 377904 376078 377913
rect 376022 377839 376078 377848
rect 377784 362681 377812 390116
rect 379532 384985 379560 390116
rect 379518 384976 379574 384985
rect 379518 384911 379574 384920
rect 381280 373969 381308 390116
rect 383028 376689 383056 390116
rect 383014 376680 383070 376689
rect 383014 376615 383070 376624
rect 381266 373960 381322 373969
rect 381266 373895 381322 373904
rect 384776 365537 384804 390116
rect 386524 377777 386552 390116
rect 386510 377768 386566 377777
rect 386510 377703 386566 377712
rect 384762 365528 384818 365537
rect 384762 365463 384818 365472
rect 377770 362672 377826 362681
rect 377770 362607 377826 362616
rect 374274 353696 374330 353705
rect 374274 353631 374330 353640
rect 388272 352889 388300 390116
rect 390020 380769 390048 390116
rect 390006 380760 390062 380769
rect 390006 380695 390062 380704
rect 391768 372201 391796 390116
rect 391754 372192 391810 372201
rect 391754 372127 391810 372136
rect 393516 369209 393544 390116
rect 394608 386572 394660 386578
rect 394608 386514 394660 386520
rect 394620 386374 394648 386514
rect 394608 386368 394660 386374
rect 394608 386310 394660 386316
rect 395264 378593 395292 390116
rect 395988 386504 396040 386510
rect 395988 386446 396040 386452
rect 396000 386306 396028 386446
rect 395988 386300 396040 386306
rect 395988 386242 396040 386248
rect 395250 378584 395306 378593
rect 395250 378519 395306 378528
rect 393502 369200 393558 369209
rect 393502 369135 393558 369144
rect 397012 364041 397040 390116
rect 398104 389904 398156 389910
rect 398104 389846 398156 389852
rect 398116 388890 398144 389846
rect 398104 388884 398156 388890
rect 398104 388826 398156 388832
rect 398760 381449 398788 390116
rect 400312 388884 400364 388890
rect 400312 388826 400364 388832
rect 398930 388784 398986 388793
rect 398930 388719 398986 388728
rect 398840 388544 398892 388550
rect 398840 388486 398892 388492
rect 398852 387841 398880 388486
rect 398838 387832 398894 387841
rect 398838 387767 398894 387776
rect 398944 387025 398972 388719
rect 400218 388240 400274 388249
rect 400218 388175 400274 388184
rect 400232 387297 400260 388175
rect 400324 387977 400352 388826
rect 400310 387968 400366 387977
rect 400310 387903 400366 387912
rect 400218 387288 400274 387297
rect 400218 387223 400274 387232
rect 398930 387016 398986 387025
rect 398930 386951 398986 386960
rect 398746 381440 398802 381449
rect 398746 381375 398802 381384
rect 400508 374921 400536 390116
rect 400494 374912 400550 374921
rect 400494 374847 400550 374856
rect 396998 364032 397054 364041
rect 396998 363967 397054 363976
rect 402256 361321 402284 390116
rect 404004 387190 404032 390116
rect 403992 387184 404044 387190
rect 403992 387126 404044 387132
rect 403622 387016 403678 387025
rect 403622 386951 403678 386960
rect 402242 361312 402298 361321
rect 402242 361247 402298 361256
rect 402244 358080 402296 358086
rect 402244 358022 402296 358028
rect 402256 353258 402284 358022
rect 403636 357785 403664 386951
rect 404266 386608 404322 386617
rect 404266 386543 404322 386552
rect 404280 386209 404308 386543
rect 404266 386200 404322 386209
rect 404266 386135 404322 386144
rect 405752 370705 405780 390116
rect 405738 370696 405794 370705
rect 405738 370631 405794 370640
rect 403622 357776 403678 357785
rect 403622 357711 403678 357720
rect 407500 355881 407528 390116
rect 408500 360936 408552 360942
rect 408500 360878 408552 360884
rect 408512 358086 408540 360878
rect 408500 358080 408552 358086
rect 408500 358022 408552 358028
rect 407486 355872 407542 355881
rect 407486 355807 407542 355816
rect 409248 353841 409276 390116
rect 410996 366489 411024 390116
rect 412744 367849 412772 390116
rect 414492 377505 414520 390116
rect 416240 383217 416268 390116
rect 417988 387161 418016 390116
rect 417974 387152 418030 387161
rect 419736 387122 419764 390116
rect 417974 387087 418030 387096
rect 419724 387116 419776 387122
rect 419724 387058 419776 387064
rect 416226 383208 416282 383217
rect 416226 383143 416282 383152
rect 414478 377496 414534 377505
rect 414478 377431 414534 377440
rect 412730 367840 412786 367849
rect 412730 367775 412786 367784
rect 410982 366480 411038 366489
rect 410982 366415 411038 366424
rect 420920 365084 420972 365090
rect 420920 365026 420972 365032
rect 420932 360942 420960 365026
rect 420920 360936 420972 360942
rect 420920 360878 420972 360884
rect 421484 357921 421512 390116
rect 421562 359408 421618 359417
rect 421562 359343 421618 359352
rect 421470 357912 421526 357921
rect 421470 357847 421526 357856
rect 409234 353832 409290 353841
rect 409234 353767 409290 353776
rect 402244 353252 402296 353258
rect 402244 353194 402296 353200
rect 388258 352880 388314 352889
rect 388258 352815 388314 352824
rect 401966 352744 402022 352753
rect 401966 352679 402022 352688
rect 373998 351928 374054 351937
rect 373998 351863 374054 351872
rect 374012 349860 374040 351863
rect 401980 349860 402008 352679
rect 421576 352617 421604 359343
rect 423232 358601 423260 390116
rect 424980 359281 425008 390116
rect 426728 360097 426756 390116
rect 426714 360088 426770 360097
rect 426714 360023 426770 360032
rect 428476 359961 428504 390116
rect 428462 359952 428518 359961
rect 428462 359887 428518 359896
rect 430224 359582 430252 390116
rect 431222 386064 431278 386073
rect 431222 385999 431278 386008
rect 430212 359576 430264 359582
rect 430212 359518 430264 359524
rect 424966 359272 425022 359281
rect 424966 359207 425022 359216
rect 423218 358592 423274 358601
rect 423218 358527 423274 358536
rect 421562 352608 421618 352617
rect 421562 352543 421618 352552
rect 431236 352073 431264 385999
rect 431972 359825 432000 390116
rect 431958 359816 432014 359825
rect 431958 359751 432014 359760
rect 433720 359689 433748 390116
rect 435468 369170 435496 390116
rect 436744 377460 436796 377466
rect 436744 377402 436796 377408
rect 435456 369164 435508 369170
rect 435456 369106 435508 369112
rect 436756 365090 436784 377402
rect 436744 365084 436796 365090
rect 436744 365026 436796 365032
rect 433706 359680 433762 359689
rect 433706 359615 433762 359624
rect 437216 356561 437244 390116
rect 438964 357377 438992 390116
rect 438950 357368 439006 357377
rect 438950 357303 439006 357312
rect 440712 357241 440740 390116
rect 440698 357232 440754 357241
rect 440698 357167 440754 357176
rect 442460 357105 442488 390116
rect 442446 357096 442502 357105
rect 442446 357031 442502 357040
rect 444208 356969 444236 390116
rect 445668 382968 445720 382974
rect 445668 382910 445720 382916
rect 445680 377466 445708 382910
rect 445668 377460 445720 377466
rect 445668 377402 445720 377408
rect 444194 356960 444250 356969
rect 444194 356895 444250 356904
rect 445956 356833 445984 390116
rect 445942 356824 445998 356833
rect 445942 356759 445998 356768
rect 447704 356697 447732 390116
rect 449452 356862 449480 390116
rect 449440 356856 449492 356862
rect 449440 356798 449492 356804
rect 451200 356794 451228 390116
rect 452948 366586 452976 390116
rect 454696 380633 454724 390116
rect 454682 380624 454738 380633
rect 454682 380559 454738 380568
rect 452936 366580 452988 366586
rect 452936 366522 452988 366528
rect 456444 365129 456472 390116
rect 458192 385937 458220 390116
rect 458178 385928 458234 385937
rect 458178 385863 458234 385872
rect 456430 365120 456486 365129
rect 456430 365055 456486 365064
rect 459940 363905 459968 390116
rect 461688 382129 461716 390116
rect 461674 382120 461730 382129
rect 461674 382055 461730 382064
rect 459926 363896 459982 363905
rect 459926 363831 459982 363840
rect 451188 356788 451240 356794
rect 451188 356730 451240 356736
rect 447690 356688 447746 356697
rect 447690 356623 447746 356632
rect 437202 356552 437258 356561
rect 437202 356487 437258 356496
rect 460938 356008 460994 356017
rect 460938 355943 460994 355952
rect 452660 355428 452712 355434
rect 452660 355370 452712 355376
rect 452672 354006 452700 355370
rect 452660 354000 452712 354006
rect 452660 353942 452712 353948
rect 457902 352608 457958 352617
rect 457902 352543 457958 352552
rect 429934 352064 429990 352073
rect 429934 351999 429990 352008
rect 431222 352064 431278 352073
rect 431222 351999 431278 352008
rect 429948 349860 429976 351999
rect 457916 349860 457944 352543
rect 460952 350554 460980 355943
rect 463436 355745 463464 390116
rect 465184 387025 465212 390116
rect 465170 387016 465226 387025
rect 465170 386951 465226 386960
rect 466368 385688 466420 385694
rect 466368 385630 466420 385636
rect 466380 382974 466408 385630
rect 466368 382968 466420 382974
rect 466368 382910 466420 382916
rect 466932 358329 466960 390116
rect 467838 360224 467894 360233
rect 467838 360159 467894 360168
rect 466918 358320 466974 358329
rect 466918 358255 466974 358264
rect 467852 356017 467880 360159
rect 468680 358193 468708 390116
rect 468666 358184 468722 358193
rect 468666 358119 468722 358128
rect 470428 358057 470456 390116
rect 471242 383208 471298 383217
rect 471242 383143 471298 383152
rect 470414 358048 470470 358057
rect 470414 357983 470470 357992
rect 467838 356008 467894 356017
rect 467838 355943 467894 355952
rect 463422 355736 463478 355745
rect 463422 355671 463478 355680
rect 471256 352617 471284 383143
rect 472176 358630 472204 390116
rect 473266 362128 473322 362137
rect 473266 362063 473322 362072
rect 473280 360233 473308 362063
rect 473266 360224 473322 360233
rect 473266 360159 473322 360168
rect 472164 358624 472216 358630
rect 472164 358566 472216 358572
rect 473924 358562 473952 390116
rect 473912 358556 473964 358562
rect 473912 358498 473964 358504
rect 475672 358494 475700 390116
rect 476394 367024 476450 367033
rect 476394 366959 476450 366968
rect 476408 362137 476436 366959
rect 476394 362128 476450 362137
rect 476394 362063 476450 362072
rect 475660 358488 475712 358494
rect 475660 358430 475712 358436
rect 477420 358426 477448 390116
rect 478878 369880 478934 369889
rect 478878 369815 478934 369824
rect 478892 367033 478920 369815
rect 479168 367810 479196 390116
rect 480916 387705 480944 390116
rect 480902 387696 480958 387705
rect 480902 387631 480958 387640
rect 479156 367804 479208 367810
rect 479156 367746 479208 367752
rect 478878 367024 478934 367033
rect 478878 366959 478934 366968
rect 477500 363792 477552 363798
rect 477500 363734 477552 363740
rect 477408 358420 477460 358426
rect 477408 358362 477460 358368
rect 477512 357678 477540 363734
rect 479522 362944 479578 362953
rect 479522 362879 479578 362888
rect 474648 357672 474700 357678
rect 474648 357614 474700 357620
rect 477500 357672 477552 357678
rect 477500 357614 477552 357620
rect 474660 355434 474688 357614
rect 474648 355428 474700 355434
rect 474648 355370 474700 355376
rect 471242 352608 471298 352617
rect 471242 352543 471298 352552
rect 479536 350713 479564 362879
rect 480916 359417 480944 387631
rect 482282 372736 482338 372745
rect 482282 372671 482338 372680
rect 482296 363225 482324 372671
rect 482282 363216 482338 363225
rect 482282 363151 482338 363160
rect 482664 359553 482692 390116
rect 484412 387161 484440 390116
rect 485780 389972 485832 389978
rect 485780 389914 485832 389920
rect 484398 387152 484454 387161
rect 484398 387087 484454 387096
rect 485792 385694 485820 389914
rect 486160 387297 486188 390116
rect 486146 387288 486202 387297
rect 486146 387223 486202 387232
rect 485870 387016 485926 387025
rect 485870 386951 485926 386960
rect 485780 385688 485832 385694
rect 485780 385630 485832 385636
rect 485410 376680 485466 376689
rect 485410 376615 485466 376624
rect 485424 371793 485452 376615
rect 485778 375864 485834 375873
rect 485778 375799 485834 375808
rect 485792 372745 485820 375799
rect 485778 372736 485834 372745
rect 485778 372671 485834 372680
rect 482834 371784 482890 371793
rect 482834 371719 482890 371728
rect 485410 371784 485466 371793
rect 485410 371719 485466 371728
rect 482848 369889 482876 371719
rect 482834 369880 482890 369889
rect 482834 369815 482890 369824
rect 482650 359544 482706 359553
rect 482650 359479 482706 359488
rect 480902 359408 480958 359417
rect 480902 359343 480958 359352
rect 476118 350704 476174 350713
rect 476118 350639 476174 350648
rect 479522 350704 479578 350713
rect 479522 350639 479578 350648
rect 460860 350526 460980 350554
rect 460860 349897 460888 350526
rect 460846 349888 460902 349897
rect 460846 349823 460902 349832
rect 476132 349761 476160 350639
rect 485884 349860 485912 386951
rect 487908 384441 487936 390116
rect 487894 384432 487950 384441
rect 487894 384367 487950 384376
rect 489656 384305 489684 390116
rect 491298 385928 491354 385937
rect 491298 385863 491354 385872
rect 489642 384296 489698 384305
rect 489642 384231 489698 384240
rect 491312 383654 491340 385863
rect 491404 385014 491432 390116
rect 498212 389910 498240 390594
rect 498200 389904 498252 389910
rect 498200 389846 498252 389852
rect 491942 387424 491998 387433
rect 491942 387359 491998 387368
rect 491392 385008 491444 385014
rect 491392 384950 491444 384956
rect 491220 383626 491340 383654
rect 490930 381032 490986 381041
rect 490930 380967 490986 380976
rect 487342 378584 487398 378593
rect 487342 378519 487398 378528
rect 487250 378040 487306 378049
rect 487250 377975 487306 377984
rect 485964 376644 486016 376650
rect 485964 376586 486016 376592
rect 485976 375465 486004 376586
rect 487264 375873 487292 377975
rect 487356 376689 487384 378519
rect 490944 378049 490972 380967
rect 491220 378593 491248 383626
rect 491956 381041 491984 387359
rect 498304 386594 498332 390623
rect 499500 387433 499528 390646
rect 499486 387424 499542 387433
rect 499486 387359 499542 387368
rect 498120 386566 498332 386594
rect 498120 385937 498148 386566
rect 498200 386436 498252 386442
rect 498200 386378 498252 386384
rect 498106 385928 498162 385937
rect 498106 385863 498162 385872
rect 498212 384402 498240 386378
rect 498200 384396 498252 384402
rect 498200 384338 498252 384344
rect 497462 384296 497518 384305
rect 497462 384231 497518 384240
rect 491942 381032 491998 381041
rect 491942 380967 491998 380976
rect 491206 378584 491262 378593
rect 491206 378519 491262 378528
rect 490930 378040 490986 378049
rect 490930 377975 490986 377984
rect 487342 376680 487398 376689
rect 487342 376615 487398 376624
rect 487250 375864 487306 375873
rect 487250 375799 487306 375808
rect 485962 375456 486018 375465
rect 485962 375391 486018 375400
rect 495440 368824 495492 368830
rect 495440 368766 495492 368772
rect 495452 366518 495480 368766
rect 487804 366512 487856 366518
rect 487804 366454 487856 366460
rect 495440 366512 495492 366518
rect 495440 366454 495492 366460
rect 487816 363798 487844 366454
rect 487804 363792 487856 363798
rect 487804 363734 487856 363740
rect 497476 352753 497504 384231
rect 498844 383716 498896 383722
rect 498844 383658 498896 383664
rect 498856 368830 498884 383658
rect 499684 373994 499712 402946
rect 499948 388544 500000 388550
rect 499948 388486 500000 388492
rect 499960 388113 499988 388486
rect 499946 388104 500002 388113
rect 499946 388039 500002 388048
rect 499762 387152 499818 387161
rect 499762 387087 499818 387096
rect 499592 373966 499712 373994
rect 498844 368824 498896 368830
rect 498844 368766 498896 368772
rect 497462 352744 497518 352753
rect 497462 352679 497518 352688
rect 476118 349752 476174 349761
rect 476118 349687 476174 349696
rect 360384 346384 360436 346390
rect 360384 346326 360436 346332
rect 360474 345808 360530 345817
rect 360474 345743 360530 345752
rect 360292 345024 360344 345030
rect 360292 344966 360344 344972
rect 360488 171134 360516 345743
rect 379624 180674 379914 180690
rect 379612 180668 379914 180674
rect 379664 180662 379914 180668
rect 488198 180674 488488 180690
rect 488198 180668 488500 180674
rect 488198 180662 488448 180668
rect 379612 180610 379664 180616
rect 488448 180610 488500 180616
rect 380808 180600 380860 180606
rect 492496 180600 492548 180606
rect 387982 180568 388038 180577
rect 380860 180548 380926 180554
rect 380808 180542 380926 180548
rect 380820 180526 380926 180542
rect 384592 180538 384974 180554
rect 384580 180532 384974 180538
rect 384632 180526 384974 180532
rect 387982 180503 388038 180512
rect 478050 180568 478106 180577
rect 489210 180538 489592 180554
rect 492246 180548 492496 180554
rect 492246 180542 492548 180548
rect 489210 180532 489604 180538
rect 489210 180526 489552 180532
rect 478050 180503 478106 180512
rect 384580 180474 384632 180480
rect 492246 180526 492536 180542
rect 489552 180474 489604 180480
rect 382556 180464 382608 180470
rect 477408 180464 477460 180470
rect 392030 180432 392086 180441
rect 382608 180412 382950 180418
rect 382556 180406 382950 180412
rect 382568 180390 382950 180406
rect 383764 180402 383962 180418
rect 383752 180396 383962 180402
rect 383804 180390 383962 180396
rect 392030 180367 392086 180376
rect 461858 180432 461914 180441
rect 477066 180412 477408 180418
rect 477066 180406 477460 180412
rect 477066 180390 477448 180406
rect 479090 180402 479472 180418
rect 479090 180396 479484 180402
rect 479090 180390 479432 180396
rect 461858 180367 461914 180376
rect 383752 180338 383804 180344
rect 479432 180338 479484 180344
rect 381636 180328 381688 180334
rect 475384 180328 475436 180334
rect 405186 180296 405242 180305
rect 381688 180276 381938 180282
rect 381636 180270 381938 180276
rect 381648 180254 381938 180270
rect 385696 180266 385986 180282
rect 385684 180260 385986 180266
rect 385736 180254 385986 180260
rect 454774 180296 454830 180305
rect 448730 180266 449112 180282
rect 448730 180260 449124 180266
rect 448730 180254 449072 180260
rect 405186 180231 405242 180240
rect 385684 180202 385736 180208
rect 475042 180276 475384 180282
rect 475042 180270 475436 180276
rect 475042 180254 475424 180270
rect 454774 180231 454830 180240
rect 449072 180202 449124 180208
rect 386604 180192 386656 180198
rect 365732 177886 365760 180132
rect 366376 180118 366758 180146
rect 366376 178022 366404 180118
rect 367008 179920 367060 179926
rect 367008 179862 367060 179868
rect 366364 178016 366416 178022
rect 366364 177958 366416 177964
rect 367020 177886 367048 179862
rect 365720 177880 365772 177886
rect 365720 177822 365772 177828
rect 367008 177880 367060 177886
rect 367008 177822 367060 177828
rect 367756 177410 367784 180132
rect 368768 177682 368796 180132
rect 369504 180118 369794 180146
rect 369504 179994 369532 180118
rect 369492 179988 369544 179994
rect 369492 179930 369544 179936
rect 369124 178696 369176 178702
rect 369124 178638 369176 178644
rect 368756 177676 368808 177682
rect 368756 177618 368808 177624
rect 369136 177410 369164 178638
rect 369860 178628 369912 178634
rect 369860 178570 369912 178576
rect 369872 177682 369900 178570
rect 370792 177954 370820 180132
rect 370780 177948 370832 177954
rect 370780 177890 370832 177896
rect 371804 177857 371832 180132
rect 372816 177993 372844 180132
rect 373828 178498 373856 180132
rect 373816 178492 373868 178498
rect 373816 178434 373868 178440
rect 372802 177984 372858 177993
rect 372802 177919 372858 177928
rect 371790 177848 371846 177857
rect 371790 177783 371846 177792
rect 374840 177721 374868 180132
rect 375576 180118 375866 180146
rect 375576 180062 375604 180118
rect 375564 180056 375616 180062
rect 375564 179998 375616 180004
rect 376864 177886 376892 180132
rect 377600 180130 377890 180146
rect 449808 180192 449860 180198
rect 421378 180160 421434 180169
rect 386656 180140 386998 180146
rect 386604 180134 386998 180140
rect 377588 180124 377890 180130
rect 377640 180118 377890 180124
rect 377588 180066 377640 180072
rect 376852 177880 376904 177886
rect 376852 177822 376904 177828
rect 374826 177712 374882 177721
rect 369860 177676 369912 177682
rect 374826 177647 374882 177656
rect 369860 177618 369912 177624
rect 367744 177404 367796 177410
rect 367744 177346 367796 177352
rect 369124 177404 369176 177410
rect 369124 177346 369176 177352
rect 378888 177274 378916 180132
rect 386616 180118 386998 180134
rect 389008 177342 389036 180132
rect 390020 178838 390048 180132
rect 390008 178832 390060 178838
rect 390008 178774 390060 178780
rect 388996 177336 389048 177342
rect 388996 177278 389048 177284
rect 378876 177268 378928 177274
rect 378876 177210 378928 177216
rect 391032 176633 391060 180132
rect 391018 176624 391074 176633
rect 393056 176594 393084 180132
rect 394068 177206 394096 180132
rect 395080 178770 395108 180132
rect 396092 179042 396120 180132
rect 396080 179036 396132 179042
rect 396080 178978 396132 178984
rect 395068 178764 395120 178770
rect 395068 178706 395120 178712
rect 394056 177200 394108 177206
rect 394056 177142 394108 177148
rect 397104 177138 397132 180132
rect 398116 178974 398144 180132
rect 398104 178968 398156 178974
rect 398104 178910 398156 178916
rect 399128 177478 399156 180132
rect 400140 177546 400168 180132
rect 401152 177614 401180 180132
rect 402164 179178 402192 180132
rect 402152 179172 402204 179178
rect 402152 179114 402204 179120
rect 403176 177750 403204 180132
rect 404188 177818 404216 180132
rect 406212 178906 406240 180132
rect 407224 179110 407252 180132
rect 407762 179888 407818 179897
rect 407762 179823 407818 179832
rect 407212 179104 407264 179110
rect 407212 179046 407264 179052
rect 406200 178900 406252 178906
rect 406200 178842 406252 178848
rect 404176 177812 404228 177818
rect 404176 177754 404228 177760
rect 403164 177744 403216 177750
rect 403164 177686 403216 177692
rect 401140 177608 401192 177614
rect 401140 177550 401192 177556
rect 400128 177540 400180 177546
rect 400128 177482 400180 177488
rect 399116 177472 399168 177478
rect 399116 177414 399168 177420
rect 397092 177132 397144 177138
rect 397092 177074 397144 177080
rect 391018 176559 391074 176568
rect 393044 176588 393096 176594
rect 393044 176530 393096 176536
rect 371056 175976 371108 175982
rect 371056 175918 371108 175924
rect 365718 173224 365774 173233
rect 365718 173159 365774 173168
rect 365732 171134 365760 173159
rect 360488 171106 361528 171134
rect 365732 171106 365944 171134
rect 360108 169312 360160 169318
rect 360108 169254 360160 169260
rect 358096 161446 358768 161474
rect 357530 147112 357586 147121
rect 357530 147047 357586 147056
rect 357346 146568 357402 146577
rect 357346 146503 357402 146512
rect 355876 146328 355928 146334
rect 355876 146270 355928 146276
rect 355888 142154 355916 146270
rect 355888 142126 356008 142154
rect 355600 120624 355652 120630
rect 355600 120566 355652 120572
rect 355416 117030 355468 117036
rect 355506 117056 355562 117065
rect 355506 116991 355562 117000
rect 355322 115832 355378 115841
rect 355980 115802 356008 142126
rect 358096 118697 358124 161446
rect 358728 147008 358780 147014
rect 358726 146976 358728 146985
rect 358780 146976 358782 146985
rect 358726 146911 358782 146920
rect 358176 146668 358228 146674
rect 358176 146610 358228 146616
rect 358082 118688 358138 118697
rect 358082 118623 358138 118632
rect 358188 117026 358216 146610
rect 358268 146600 358320 146606
rect 358268 146542 358320 146548
rect 358280 117298 358308 146542
rect 359556 146532 359608 146538
rect 359556 146474 359608 146480
rect 359464 146396 359516 146402
rect 359464 146338 359516 146344
rect 358542 144528 358598 144537
rect 358360 144492 358412 144498
rect 358542 144463 358598 144472
rect 358360 144434 358412 144440
rect 358268 117292 358320 117298
rect 358268 117234 358320 117240
rect 358372 117230 358400 144434
rect 358452 144288 358504 144294
rect 358452 144230 358504 144236
rect 358360 117224 358412 117230
rect 358360 117166 358412 117172
rect 358464 117162 358492 144230
rect 358556 119746 358584 144463
rect 358636 144424 358688 144430
rect 358636 144366 358688 144372
rect 358648 120086 358676 144366
rect 358636 120080 358688 120086
rect 358636 120022 358688 120028
rect 358544 119740 358596 119746
rect 358544 119682 358596 119688
rect 359476 118046 359504 146338
rect 359568 118522 359596 146474
rect 361500 144922 361528 171106
rect 364982 169008 365038 169017
rect 364982 168943 365038 168952
rect 363602 166288 363658 166297
rect 363602 166223 363658 166232
rect 363616 147014 363644 166223
rect 363604 147008 363656 147014
rect 363604 146950 363656 146956
rect 362868 146804 362920 146810
rect 362868 146746 362920 146752
rect 362880 146470 362908 146746
rect 362776 146464 362828 146470
rect 362776 146406 362828 146412
rect 362868 146464 362920 146470
rect 362868 146406 362920 146412
rect 362788 146334 362816 146406
rect 362684 146328 362736 146334
rect 362684 146270 362736 146276
rect 362776 146328 362828 146334
rect 362776 146270 362828 146276
rect 360764 144908 361528 144922
rect 362696 144908 362724 146270
rect 363616 144922 363644 146950
rect 364996 146946 365024 168943
rect 364984 146940 365036 146946
rect 364984 146882 365036 146888
rect 364996 144922 365024 146882
rect 365916 146742 365944 171106
rect 369858 167648 369914 167657
rect 369858 167583 369914 167592
rect 368664 164892 368716 164898
rect 368664 164834 368716 164840
rect 367466 147112 367522 147121
rect 367466 147047 367522 147056
rect 365904 146736 365956 146742
rect 365904 146678 365956 146684
rect 365916 144922 365944 146678
rect 360764 144894 361514 144908
rect 363616 144894 363906 144922
rect 364996 144894 365102 144922
rect 365916 144894 366298 144922
rect 367480 144908 367508 147047
rect 368676 144908 368704 164834
rect 369872 144908 369900 167583
rect 371068 144908 371096 175918
rect 407118 172544 407174 172553
rect 407118 172479 407174 172488
rect 402978 171728 403034 171737
rect 402978 171663 403034 171672
rect 372252 170400 372304 170406
rect 372252 170342 372304 170348
rect 372264 144908 372292 170342
rect 393780 169312 393832 169318
rect 393780 169254 393832 169260
rect 377036 169244 377088 169250
rect 377036 169186 377088 169192
rect 373448 160744 373500 160750
rect 373448 160686 373500 160692
rect 373460 144908 373488 160686
rect 375838 151192 375894 151201
rect 375838 151127 375894 151136
rect 374644 149728 374696 149734
rect 374644 149670 374696 149676
rect 374656 144908 374684 149670
rect 375852 144908 375880 151127
rect 377048 144908 377076 169186
rect 384212 162172 384264 162178
rect 384212 162114 384264 162120
rect 383014 148608 383070 148617
rect 383014 148543 383070 148552
rect 379426 148472 379482 148481
rect 379426 148407 379482 148416
rect 381820 148436 381872 148442
rect 378230 148336 378286 148345
rect 378230 148271 378286 148280
rect 378244 144908 378272 148271
rect 379440 144908 379468 148407
rect 381820 148378 381872 148384
rect 380624 148368 380676 148374
rect 380624 148310 380676 148316
rect 380636 144908 380664 148310
rect 381832 144908 381860 148378
rect 383028 144908 383056 148543
rect 384224 144908 384252 162114
rect 388996 146668 389048 146674
rect 388996 146610 389048 146616
rect 389008 144908 389036 146610
rect 390192 146600 390244 146606
rect 390192 146542 390244 146548
rect 390204 144908 390232 146542
rect 392584 146532 392636 146538
rect 392584 146474 392636 146480
rect 391388 146464 391440 146470
rect 391388 146406 391440 146412
rect 391400 144908 391428 146406
rect 392596 144908 392624 146474
rect 393792 144908 393820 169254
rect 394974 169144 395030 169153
rect 394974 169079 395030 169088
rect 394988 144908 395016 169079
rect 400954 147248 401010 147257
rect 400954 147183 401010 147192
rect 399758 146704 399814 146713
rect 399758 146639 399814 146648
rect 397368 146396 397420 146402
rect 397368 146338 397420 146344
rect 397380 144908 397408 146338
rect 398564 146328 398616 146334
rect 398564 146270 398616 146276
rect 398576 144908 398604 146270
rect 399772 144908 399800 146639
rect 400968 144908 400996 147183
rect 402150 146568 402206 146577
rect 402150 146503 402206 146512
rect 402164 144908 402192 146503
rect 402992 146441 403020 171663
rect 402978 146432 403034 146441
rect 402978 146367 403034 146376
rect 402992 144922 403020 146367
rect 402992 144894 403374 144922
rect 359648 144356 359700 144362
rect 359648 144298 359700 144304
rect 359556 118516 359608 118522
rect 359556 118458 359608 118464
rect 359660 118386 359688 144298
rect 360764 122834 360792 144894
rect 386432 144498 386630 144514
rect 386420 144492 386630 144498
rect 386472 144486 386630 144492
rect 386420 144434 386472 144440
rect 385132 144424 385184 144430
rect 396170 144392 396226 144401
rect 385184 144372 385434 144378
rect 385132 144366 385434 144372
rect 385144 144350 385434 144366
rect 387720 144350 387826 144378
rect 387720 144294 387748 144350
rect 396170 144327 396226 144336
rect 387708 144288 387760 144294
rect 387708 144230 387760 144236
rect 360672 122806 360792 122834
rect 359648 118380 359700 118386
rect 359648 118322 359700 118328
rect 359464 118040 359516 118046
rect 359464 117982 359516 117988
rect 360672 117978 360700 122806
rect 360660 117972 360712 117978
rect 360660 117914 360712 117920
rect 358452 117156 358504 117162
rect 358452 117098 358504 117104
rect 358176 117020 358228 117026
rect 358176 116962 358228 116968
rect 355322 115767 355378 115776
rect 355968 115796 356020 115802
rect 355968 115738 356020 115744
rect 358084 115796 358136 115802
rect 358084 115738 358136 115744
rect 352930 115424 352986 115433
rect 352930 115359 352986 115368
rect 358096 86970 358124 115738
rect 360672 89010 360700 117914
rect 407132 105777 407160 172479
rect 407210 144800 407266 144809
rect 407210 144735 407266 144744
rect 407224 139233 407252 144735
rect 407776 144362 407804 179823
rect 408236 179246 408264 180132
rect 409248 179314 409276 180132
rect 410260 179353 410288 180132
rect 410246 179344 410302 179353
rect 409236 179308 409288 179314
rect 410246 179279 410302 179288
rect 409236 179250 409288 179256
rect 408224 179240 408276 179246
rect 408224 179182 408276 179188
rect 411272 179081 411300 180132
rect 411258 179072 411314 179081
rect 411258 179007 411314 179016
rect 412284 177410 412312 180132
rect 413296 177585 413324 180132
rect 414308 178945 414336 180132
rect 415320 179353 415348 180132
rect 415306 179344 415362 179353
rect 415306 179279 415362 179288
rect 414294 178936 414350 178945
rect 414294 178871 414350 178880
rect 413282 177576 413338 177585
rect 413282 177511 413338 177520
rect 412272 177404 412324 177410
rect 412272 177346 412324 177352
rect 416332 175234 416360 180132
rect 417344 176662 417372 180132
rect 417332 176656 417384 176662
rect 417332 176598 417384 176604
rect 418356 175273 418384 180132
rect 419368 177682 419396 180132
rect 419356 177676 419408 177682
rect 419356 177618 419408 177624
rect 420380 176633 420408 180132
rect 441618 180160 441674 180169
rect 421378 180095 421434 180104
rect 420366 176624 420422 176633
rect 420366 176559 420422 176568
rect 418342 175264 418398 175273
rect 416320 175228 416372 175234
rect 418342 175199 418398 175208
rect 416320 175170 416372 175176
rect 422404 175137 422432 180132
rect 423416 179382 423444 180132
rect 423404 179376 423456 179382
rect 423404 179318 423456 179324
rect 424428 176089 424456 180132
rect 424414 176080 424470 176089
rect 424414 176015 424470 176024
rect 422390 175128 422446 175137
rect 422390 175063 422446 175072
rect 425440 175001 425468 180132
rect 426452 176662 426480 180132
rect 427464 178022 427492 180132
rect 427452 178016 427504 178022
rect 427452 177958 427504 177964
rect 426440 176656 426492 176662
rect 426440 176598 426492 176604
rect 425426 174992 425482 175001
rect 425426 174927 425482 174936
rect 428476 174865 428504 180132
rect 429488 176458 429516 180132
rect 429476 176452 429528 176458
rect 429476 176394 429528 176400
rect 430500 175166 430528 180132
rect 430488 175160 430540 175166
rect 430488 175102 430540 175108
rect 428462 174856 428518 174865
rect 428462 174791 428518 174800
rect 431512 174593 431540 180132
rect 432524 174729 432552 180132
rect 433536 176361 433564 180132
rect 433522 176352 433578 176361
rect 434548 176322 434576 180132
rect 433522 176287 433578 176296
rect 434536 176316 434588 176322
rect 434536 176258 434588 176264
rect 435560 176225 435588 180132
rect 435546 176216 435602 176225
rect 435546 176151 435602 176160
rect 436572 175030 436600 180132
rect 437584 176497 437612 180132
rect 438596 177313 438624 180132
rect 438582 177304 438638 177313
rect 438582 177239 438638 177248
rect 437570 176488 437626 176497
rect 437570 176423 437626 176432
rect 436560 175024 436612 175030
rect 436560 174966 436612 174972
rect 432510 174720 432566 174729
rect 432510 174655 432566 174664
rect 431498 174584 431554 174593
rect 431498 174519 431554 174528
rect 439608 174457 439636 180132
rect 440620 176390 440648 180132
rect 449742 180140 449808 180146
rect 449742 180134 449860 180140
rect 441618 180095 441674 180104
rect 442644 178634 442672 180132
rect 443656 178906 443684 180132
rect 444668 178974 444696 180132
rect 444656 178968 444708 178974
rect 444656 178910 444708 178916
rect 443644 178900 443696 178906
rect 443644 178842 443696 178848
rect 442632 178628 442684 178634
rect 442632 178570 442684 178576
rect 445680 176594 445708 180132
rect 446692 178770 446720 180132
rect 446680 178764 446732 178770
rect 446680 178706 446732 178712
rect 445668 176588 445720 176594
rect 445668 176530 445720 176536
rect 440608 176384 440660 176390
rect 440608 176326 440660 176332
rect 447704 175098 447732 180132
rect 449742 180118 449848 180134
rect 447692 175092 447744 175098
rect 447692 175034 447744 175040
rect 450740 174962 450768 180132
rect 451752 179382 451780 180132
rect 451740 179376 451792 179382
rect 451740 179318 451792 179324
rect 452764 176526 452792 180132
rect 453776 177274 453804 180132
rect 455800 179314 455828 180132
rect 455788 179308 455840 179314
rect 455788 179250 455840 179256
rect 456812 178809 456840 180132
rect 457824 178945 457852 180132
rect 458836 179246 458864 180132
rect 458824 179240 458876 179246
rect 458824 179182 458876 179188
rect 459848 179178 459876 180132
rect 459836 179172 459888 179178
rect 459836 179114 459888 179120
rect 460860 179110 460888 180132
rect 460848 179104 460900 179110
rect 462884 179081 462912 180132
rect 460848 179046 460900 179052
rect 462870 179072 462926 179081
rect 463896 179042 463924 180132
rect 462870 179007 462926 179016
rect 463884 179036 463936 179042
rect 463884 178978 463936 178984
rect 457810 178936 457866 178945
rect 457810 178871 457866 178880
rect 456798 178800 456854 178809
rect 456798 178735 456854 178744
rect 464908 178702 464936 180132
rect 465920 178838 465948 180132
rect 465908 178832 465960 178838
rect 465908 178774 465960 178780
rect 464896 178696 464948 178702
rect 464896 178638 464948 178644
rect 466932 177886 466960 180132
rect 467944 177954 467972 180132
rect 467932 177948 467984 177954
rect 467932 177890 467984 177896
rect 466920 177880 466972 177886
rect 466920 177822 466972 177828
rect 468956 177818 468984 180132
rect 468944 177812 468996 177818
rect 468944 177754 468996 177760
rect 469968 177410 469996 180132
rect 469956 177404 470008 177410
rect 469956 177346 470008 177352
rect 470980 177342 471008 180132
rect 471992 177857 472020 180132
rect 473004 178022 473032 180132
rect 474016 179761 474044 180132
rect 476054 180130 476160 180146
rect 480102 180130 480208 180146
rect 476054 180124 476172 180130
rect 476054 180118 476120 180124
rect 480102 180124 480220 180130
rect 480102 180118 480168 180124
rect 476120 180066 476172 180072
rect 480168 180066 480220 180072
rect 474002 179752 474058 179761
rect 474002 179687 474058 179696
rect 472992 178016 473044 178022
rect 472992 177958 473044 177964
rect 471978 177848 472034 177857
rect 471978 177783 472034 177792
rect 481100 177585 481128 180132
rect 482112 177614 482140 180132
rect 483124 177750 483152 180132
rect 483112 177744 483164 177750
rect 483112 177686 483164 177692
rect 482100 177608 482152 177614
rect 481086 177576 481142 177585
rect 482100 177550 482152 177556
rect 481086 177511 481142 177520
rect 484136 177478 484164 180132
rect 485148 177546 485176 180132
rect 486160 177682 486188 180132
rect 487172 177721 487200 180132
rect 490208 177993 490236 180132
rect 491128 180118 491234 180146
rect 491128 180062 491156 180118
rect 491116 180056 491168 180062
rect 491116 179998 491168 180004
rect 490194 177984 490250 177993
rect 490194 177919 490250 177928
rect 487158 177712 487214 177721
rect 486148 177676 486200 177682
rect 487158 177647 487214 177656
rect 486148 177618 486200 177624
rect 485136 177540 485188 177546
rect 485136 177482 485188 177488
rect 484124 177472 484176 177478
rect 493244 177449 493272 180132
rect 484124 177414 484176 177420
rect 493230 177440 493286 177449
rect 493230 177375 493286 177384
rect 470968 177336 471020 177342
rect 470968 177278 471020 177284
rect 453764 177268 453816 177274
rect 453764 177210 453816 177216
rect 494256 177206 494284 180132
rect 499592 178022 499620 373966
rect 499672 363724 499724 363730
rect 499672 363666 499724 363672
rect 499684 202745 499712 363666
rect 499670 202736 499726 202745
rect 499670 202671 499726 202680
rect 499776 179897 499804 387087
rect 499762 179888 499818 179897
rect 499762 179823 499818 179832
rect 499580 178016 499632 178022
rect 499580 177958 499632 177964
rect 494244 177200 494296 177206
rect 494244 177142 494296 177148
rect 452752 176520 452804 176526
rect 452752 176462 452804 176468
rect 450728 174956 450780 174962
rect 450728 174898 450780 174904
rect 439594 174448 439650 174457
rect 439594 174383 439650 174392
rect 500236 159769 500264 441934
rect 500328 390658 500356 513266
rect 500512 512650 500540 524386
rect 500960 521892 501012 521898
rect 500960 521834 501012 521840
rect 500592 521824 500644 521830
rect 500592 521766 500644 521772
rect 500866 521792 500922 521801
rect 500500 512644 500552 512650
rect 500500 512586 500552 512592
rect 500604 511873 500632 521766
rect 500866 521727 500922 521736
rect 500776 520940 500828 520946
rect 500776 520882 500828 520888
rect 500684 520872 500736 520878
rect 500684 520814 500736 520820
rect 500696 520266 500724 520814
rect 500684 520260 500736 520266
rect 500684 520202 500736 520208
rect 500788 519330 500816 520882
rect 500880 519897 500908 521727
rect 500866 519888 500922 519897
rect 500866 519823 500922 519832
rect 500866 519344 500922 519353
rect 500788 519302 500866 519330
rect 500866 519279 500922 519288
rect 500972 513330 501000 521834
rect 500960 513324 501012 513330
rect 500960 513266 501012 513272
rect 500590 511864 500646 511873
rect 500590 511799 500646 511808
rect 500408 511284 500460 511290
rect 500408 511226 500460 511232
rect 500316 390652 500368 390658
rect 500316 390594 500368 390600
rect 500420 390046 500448 511226
rect 500590 488336 500646 488345
rect 500590 488271 500646 488280
rect 500500 486124 500552 486130
rect 500500 486066 500552 486072
rect 500512 482361 500540 486066
rect 500498 482352 500554 482361
rect 500498 482287 500554 482296
rect 500498 474600 500554 474609
rect 500498 474535 500554 474544
rect 500408 390040 500460 390046
rect 500408 389982 500460 389988
rect 500512 388929 500540 474535
rect 500604 391921 500632 488271
rect 500866 451208 500922 451217
rect 500866 451143 500922 451152
rect 500880 441998 500908 451143
rect 500868 441992 500920 441998
rect 500868 441934 500920 441940
rect 501064 438841 501092 538426
rect 501156 442921 501184 541583
rect 501236 521348 501288 521354
rect 501236 521290 501288 521296
rect 501248 519858 501276 521290
rect 501328 521212 501380 521218
rect 501328 521154 501380 521160
rect 501340 519858 501368 521154
rect 501236 519852 501288 519858
rect 501236 519794 501288 519800
rect 501328 519852 501380 519858
rect 501328 519794 501380 519800
rect 501248 519722 501368 519738
rect 501248 519716 501380 519722
rect 501248 519710 501328 519716
rect 501142 442912 501198 442921
rect 501142 442847 501198 442856
rect 501248 441561 501276 519710
rect 501328 519658 501380 519664
rect 501328 519580 501380 519586
rect 501328 519522 501380 519528
rect 501340 443193 501368 519522
rect 501432 479913 501460 559671
rect 501602 554568 501658 554577
rect 501602 554503 501658 554512
rect 501510 523288 501566 523297
rect 501510 523223 501566 523232
rect 501418 479904 501474 479913
rect 501418 479839 501474 479848
rect 501524 443737 501552 523223
rect 501616 483993 501644 554503
rect 501800 526726 501828 600100
rect 503180 598913 503208 600100
rect 503166 598904 503222 598913
rect 503166 598839 503222 598848
rect 504560 598097 504588 600100
rect 504822 600063 504878 600072
rect 504546 598088 504602 598097
rect 504546 598023 504602 598032
rect 504836 586514 504864 600063
rect 505098 599584 505154 599593
rect 505098 599519 505154 599528
rect 504744 586486 504864 586514
rect 503996 558272 504048 558278
rect 503996 558214 504048 558220
rect 502338 552528 502394 552537
rect 502338 552463 502394 552472
rect 502062 551032 502118 551041
rect 502062 550967 502118 550976
rect 501880 529576 501932 529582
rect 501880 529518 501932 529524
rect 501788 526720 501840 526726
rect 501788 526662 501840 526668
rect 501696 526244 501748 526250
rect 501696 526186 501748 526192
rect 501708 519586 501736 526186
rect 501788 521280 501840 521286
rect 501788 521222 501840 521228
rect 501696 519580 501748 519586
rect 501696 519522 501748 519528
rect 501800 519194 501828 521222
rect 501892 519654 501920 529518
rect 501970 522200 502026 522209
rect 501970 522135 502026 522144
rect 501880 519648 501932 519654
rect 501880 519590 501932 519596
rect 501878 519208 501934 519217
rect 501800 519166 501878 519194
rect 501878 519143 501934 519152
rect 501984 509234 502012 522135
rect 501708 509206 502012 509234
rect 501602 483984 501658 483993
rect 501602 483919 501658 483928
rect 501604 483676 501656 483682
rect 501604 483618 501656 483624
rect 501510 443728 501566 443737
rect 501510 443663 501566 443672
rect 501326 443184 501382 443193
rect 501326 443119 501382 443128
rect 501234 441552 501290 441561
rect 501234 441487 501290 441496
rect 501050 438832 501106 438841
rect 501050 438767 501106 438776
rect 500682 404968 500738 404977
rect 500682 404903 500738 404912
rect 500590 391912 500646 391921
rect 500590 391847 500646 391856
rect 500696 389065 500724 404903
rect 500682 389056 500738 389065
rect 500682 388991 500738 389000
rect 500498 388920 500554 388929
rect 500498 388855 500554 388864
rect 500958 387288 501014 387297
rect 500958 387223 501014 387232
rect 500972 181393 501000 387223
rect 501144 366376 501196 366382
rect 501144 366318 501196 366324
rect 501050 360904 501106 360913
rect 501050 360839 501106 360848
rect 501064 190369 501092 360839
rect 501156 208321 501184 366318
rect 501236 349920 501288 349926
rect 501236 349862 501288 349868
rect 501142 208312 501198 208321
rect 501142 208247 501198 208256
rect 501248 196761 501276 349862
rect 501234 196752 501290 196761
rect 501234 196687 501290 196696
rect 501050 190360 501106 190369
rect 501050 190295 501106 190304
rect 500958 181384 501014 181393
rect 500958 181319 501014 181328
rect 501616 178634 501644 483618
rect 501708 474609 501736 509206
rect 501694 474600 501750 474609
rect 501694 474535 501750 474544
rect 501696 457496 501748 457502
rect 501696 457438 501748 457444
rect 501708 390250 501736 457438
rect 502076 442649 502104 550967
rect 502156 528080 502208 528086
rect 502156 528022 502208 528028
rect 502168 519722 502196 528022
rect 502246 520296 502302 520305
rect 502246 520231 502302 520240
rect 502260 519926 502288 520231
rect 502248 519920 502300 519926
rect 502248 519862 502300 519868
rect 502248 519784 502300 519790
rect 502248 519726 502300 519732
rect 502156 519716 502208 519722
rect 502156 519658 502208 519664
rect 502154 519072 502210 519081
rect 502260 519058 502288 519726
rect 502210 519030 502288 519058
rect 502154 519007 502210 519016
rect 502246 512000 502302 512009
rect 502246 511935 502302 511944
rect 502260 485874 502288 511935
rect 502352 499574 502380 552463
rect 503534 551168 503590 551177
rect 503534 551103 503590 551112
rect 502522 547768 502578 547777
rect 502522 547703 502578 547712
rect 502352 499546 502472 499574
rect 502260 485846 502380 485874
rect 502352 485450 502380 485846
rect 502340 485444 502392 485450
rect 502340 485386 502392 485392
rect 502444 485330 502472 499546
rect 502260 485302 502472 485330
rect 502260 485058 502288 485302
rect 502432 485240 502484 485246
rect 502432 485182 502484 485188
rect 502260 485030 502380 485058
rect 502352 482089 502380 485030
rect 502338 482080 502394 482089
rect 502338 482015 502394 482024
rect 502338 481400 502394 481409
rect 502338 481335 502394 481344
rect 502062 442640 502118 442649
rect 502062 442575 502118 442584
rect 501880 440360 501932 440366
rect 501880 440302 501932 440308
rect 501788 440292 501840 440298
rect 501788 440234 501840 440240
rect 501696 390244 501748 390250
rect 501696 390186 501748 390192
rect 501800 383722 501828 440234
rect 501892 389978 501920 440302
rect 502352 422294 502380 481335
rect 502444 440298 502472 485182
rect 502536 483449 502564 547703
rect 502614 543688 502670 543697
rect 502614 543623 502670 543632
rect 502628 483721 502656 543623
rect 502706 538656 502762 538665
rect 502706 538591 502762 538600
rect 502720 484537 502748 538591
rect 502798 534576 502854 534585
rect 502798 534511 502854 534520
rect 502706 484528 502762 484537
rect 502706 484463 502762 484472
rect 502706 483984 502762 483993
rect 502706 483919 502762 483928
rect 502614 483712 502670 483721
rect 502614 483647 502670 483656
rect 502522 483440 502578 483449
rect 502522 483375 502578 483384
rect 502720 480254 502748 483919
rect 502812 482905 502840 534511
rect 502892 528284 502944 528290
rect 502892 528226 502944 528232
rect 502798 482896 502854 482905
rect 502798 482831 502854 482840
rect 502904 482633 502932 528226
rect 503074 525464 503130 525473
rect 503074 525399 503130 525408
rect 503088 486441 503116 525399
rect 503258 523424 503314 523433
rect 503258 523359 503314 523368
rect 503166 520296 503222 520305
rect 503166 520231 503222 520240
rect 503074 486432 503130 486441
rect 503074 486367 503130 486376
rect 503180 485897 503208 520231
rect 503166 485888 503222 485897
rect 503166 485823 503222 485832
rect 502984 485104 503036 485110
rect 502984 485046 503036 485052
rect 502890 482624 502946 482633
rect 502890 482559 502946 482568
rect 502996 480894 503024 485046
rect 503168 482316 503220 482322
rect 503168 482258 503220 482264
rect 503076 481772 503128 481778
rect 503076 481714 503128 481720
rect 502984 480888 503036 480894
rect 502984 480830 503036 480836
rect 502720 480226 503024 480254
rect 502892 470552 502944 470558
rect 502892 470494 502944 470500
rect 502904 469305 502932 470494
rect 502890 469296 502946 469305
rect 502890 469231 502946 469240
rect 502892 469192 502944 469198
rect 502892 469134 502944 469140
rect 502800 469124 502852 469130
rect 502800 469066 502852 469072
rect 502812 468217 502840 469066
rect 502904 468489 502932 469134
rect 502890 468480 502946 468489
rect 502890 468415 502946 468424
rect 502798 468208 502854 468217
rect 502798 468143 502854 468152
rect 502708 467832 502760 467838
rect 502708 467774 502760 467780
rect 502720 466857 502748 467774
rect 502800 467764 502852 467770
rect 502800 467706 502852 467712
rect 502706 466848 502762 466857
rect 502706 466783 502762 466792
rect 502812 466585 502840 467706
rect 502892 467696 502944 467702
rect 502892 467638 502944 467644
rect 502904 467401 502932 467638
rect 502890 467392 502946 467401
rect 502890 467327 502946 467336
rect 502798 466576 502854 466585
rect 502798 466511 502854 466520
rect 502708 466404 502760 466410
rect 502708 466346 502760 466352
rect 502616 466336 502668 466342
rect 502616 466278 502668 466284
rect 502628 465497 502656 466278
rect 502720 466041 502748 466346
rect 502890 466304 502946 466313
rect 502800 466268 502852 466274
rect 502890 466239 502946 466248
rect 502800 466210 502852 466216
rect 502706 466032 502762 466041
rect 502706 465967 502762 465976
rect 502812 465769 502840 466210
rect 502904 466206 502932 466239
rect 502892 466200 502944 466206
rect 502892 466142 502944 466148
rect 502798 465760 502854 465769
rect 502798 465695 502854 465704
rect 502614 465488 502670 465497
rect 502614 465423 502670 465432
rect 502892 465044 502944 465050
rect 502892 464986 502944 464992
rect 502904 464137 502932 464986
rect 502890 464128 502946 464137
rect 502890 464063 502946 464072
rect 502616 463684 502668 463690
rect 502616 463626 502668 463632
rect 502628 462505 502656 463626
rect 502708 463616 502760 463622
rect 502708 463558 502760 463564
rect 502720 463321 502748 463558
rect 502800 463548 502852 463554
rect 502800 463490 502852 463496
rect 502706 463312 502762 463321
rect 502706 463247 502762 463256
rect 502812 462777 502840 463490
rect 502892 463480 502944 463486
rect 502892 463422 502944 463428
rect 502904 463049 502932 463422
rect 502890 463040 502946 463049
rect 502890 462975 502946 462984
rect 502798 462768 502854 462777
rect 502798 462703 502854 462712
rect 502614 462496 502670 462505
rect 502614 462431 502670 462440
rect 502524 462324 502576 462330
rect 502524 462266 502576 462272
rect 502536 461961 502564 462266
rect 502892 462256 502944 462262
rect 502890 462224 502892 462233
rect 502944 462224 502946 462233
rect 502616 462188 502668 462194
rect 502890 462159 502946 462168
rect 502616 462130 502668 462136
rect 502522 461952 502578 461961
rect 502522 461887 502578 461896
rect 502628 461417 502656 462130
rect 502892 462120 502944 462126
rect 502892 462062 502944 462068
rect 502800 462052 502852 462058
rect 502800 461994 502852 462000
rect 502614 461408 502670 461417
rect 502614 461343 502670 461352
rect 502812 461145 502840 461994
rect 502904 461689 502932 462062
rect 502890 461680 502946 461689
rect 502890 461615 502946 461624
rect 502798 461136 502854 461145
rect 502798 461071 502854 461080
rect 502800 460896 502852 460902
rect 502800 460838 502852 460844
rect 502812 460601 502840 460838
rect 502892 460828 502944 460834
rect 502892 460770 502944 460776
rect 502798 460592 502854 460601
rect 502798 460527 502854 460536
rect 502904 460329 502932 460770
rect 502890 460320 502946 460329
rect 502890 460255 502946 460264
rect 502616 459536 502668 459542
rect 502616 459478 502668 459484
rect 502628 458969 502656 459478
rect 502892 459468 502944 459474
rect 502892 459410 502944 459416
rect 502800 459400 502852 459406
rect 502800 459342 502852 459348
rect 502708 459332 502760 459338
rect 502708 459274 502760 459280
rect 502614 458960 502670 458969
rect 502614 458895 502670 458904
rect 502720 458425 502748 459274
rect 502812 458697 502840 459342
rect 502904 459241 502932 459410
rect 502890 459232 502946 459241
rect 502890 459167 502946 459176
rect 502798 458688 502854 458697
rect 502798 458623 502854 458632
rect 502706 458416 502762 458425
rect 502706 458351 502762 458360
rect 502800 458176 502852 458182
rect 502800 458118 502852 458124
rect 502890 458144 502946 458153
rect 502616 458108 502668 458114
rect 502616 458050 502668 458056
rect 502628 457065 502656 458050
rect 502708 458040 502760 458046
rect 502708 457982 502760 457988
rect 502720 457337 502748 457982
rect 502812 457881 502840 458118
rect 502890 458079 502946 458088
rect 502904 457978 502932 458079
rect 502892 457972 502944 457978
rect 502892 457914 502944 457920
rect 502798 457872 502854 457881
rect 502798 457807 502854 457816
rect 502706 457328 502762 457337
rect 502706 457263 502762 457272
rect 502614 457056 502670 457065
rect 502614 456991 502670 457000
rect 502890 456784 502946 456793
rect 502616 456748 502668 456754
rect 502890 456719 502946 456728
rect 502616 456690 502668 456696
rect 502628 455705 502656 456690
rect 502904 456686 502932 456719
rect 502892 456680 502944 456686
rect 502892 456622 502944 456628
rect 502800 456612 502852 456618
rect 502800 456554 502852 456560
rect 502812 455977 502840 456554
rect 502892 456544 502944 456550
rect 502890 456512 502892 456521
rect 502944 456512 502946 456521
rect 502890 456447 502946 456456
rect 502798 455968 502854 455977
rect 502798 455903 502854 455912
rect 502614 455696 502670 455705
rect 502614 455631 502670 455640
rect 502798 455424 502854 455433
rect 502708 455388 502760 455394
rect 502798 455359 502854 455368
rect 502708 455330 502760 455336
rect 502524 455320 502576 455326
rect 502524 455262 502576 455268
rect 502536 454073 502564 455262
rect 502616 455252 502668 455258
rect 502616 455194 502668 455200
rect 502628 454345 502656 455194
rect 502720 454889 502748 455330
rect 502812 455190 502840 455359
rect 502800 455184 502852 455190
rect 502800 455126 502852 455132
rect 502890 455152 502946 455161
rect 502890 455087 502892 455096
rect 502944 455087 502946 455096
rect 502892 455058 502944 455064
rect 502706 454880 502762 454889
rect 502706 454815 502762 454824
rect 502614 454336 502670 454345
rect 502614 454271 502670 454280
rect 502522 454064 502578 454073
rect 502522 453999 502578 454008
rect 502892 453960 502944 453966
rect 502892 453902 502944 453908
rect 502708 453892 502760 453898
rect 502708 453834 502760 453840
rect 502720 452713 502748 453834
rect 502800 453824 502852 453830
rect 502904 453801 502932 453902
rect 502800 453766 502852 453772
rect 502890 453792 502946 453801
rect 502812 453257 502840 453766
rect 502890 453727 502946 453736
rect 502798 453248 502854 453257
rect 502798 453183 502854 453192
rect 502706 452704 502762 452713
rect 502706 452639 502762 452648
rect 502708 452600 502760 452606
rect 502708 452542 502760 452548
rect 502616 452532 502668 452538
rect 502616 452474 502668 452480
rect 502628 451625 502656 452474
rect 502720 452169 502748 452542
rect 502892 452464 502944 452470
rect 502890 452432 502892 452441
rect 502944 452432 502946 452441
rect 502800 452396 502852 452402
rect 502890 452367 502946 452376
rect 502800 452338 502852 452344
rect 502706 452160 502762 452169
rect 502706 452095 502762 452104
rect 502812 451897 502840 452338
rect 502798 451888 502854 451897
rect 502798 451823 502854 451832
rect 502614 451616 502670 451625
rect 502614 451551 502670 451560
rect 502616 451240 502668 451246
rect 502616 451182 502668 451188
rect 502628 449993 502656 451182
rect 502708 451172 502760 451178
rect 502708 451114 502760 451120
rect 502720 450537 502748 451114
rect 502892 451036 502944 451042
rect 502892 450978 502944 450984
rect 502706 450528 502762 450537
rect 502706 450463 502762 450472
rect 502904 450265 502932 450978
rect 502890 450256 502946 450265
rect 502890 450191 502946 450200
rect 502614 449984 502670 449993
rect 502614 449919 502670 449928
rect 502708 449812 502760 449818
rect 502708 449754 502760 449760
rect 502720 448905 502748 449754
rect 502800 449744 502852 449750
rect 502800 449686 502852 449692
rect 502706 448896 502762 448905
rect 502706 448831 502762 448840
rect 502812 448633 502840 449686
rect 502892 449676 502944 449682
rect 502892 449618 502944 449624
rect 502904 449177 502932 449618
rect 502890 449168 502946 449177
rect 502890 449103 502946 449112
rect 502798 448624 502854 448633
rect 502798 448559 502854 448568
rect 502708 448520 502760 448526
rect 502708 448462 502760 448468
rect 502616 448452 502668 448458
rect 502616 448394 502668 448400
rect 502628 447545 502656 448394
rect 502720 447817 502748 448462
rect 502892 448316 502944 448322
rect 502892 448258 502944 448264
rect 502904 448089 502932 448258
rect 502890 448080 502946 448089
rect 502890 448015 502946 448024
rect 502706 447808 502762 447817
rect 502706 447743 502762 447752
rect 502614 447536 502670 447545
rect 502614 447471 502670 447480
rect 502432 440292 502484 440298
rect 502432 440234 502484 440240
rect 502892 436824 502944 436830
rect 502892 436766 502944 436772
rect 502800 434716 502852 434722
rect 502800 434658 502852 434664
rect 502812 434217 502840 434658
rect 502798 434208 502854 434217
rect 502798 434143 502854 434152
rect 502616 433288 502668 433294
rect 502616 433230 502668 433236
rect 502628 432857 502656 433230
rect 502614 432848 502670 432857
rect 502614 432783 502670 432792
rect 502524 431452 502576 431458
rect 502524 431394 502576 431400
rect 502536 430953 502564 431394
rect 502708 431316 502760 431322
rect 502708 431258 502760 431264
rect 502522 430944 502578 430953
rect 502522 430879 502578 430888
rect 502720 430681 502748 431258
rect 502706 430672 502762 430681
rect 502706 430607 502762 430616
rect 502616 430568 502668 430574
rect 502616 430510 502668 430516
rect 502628 430137 502656 430510
rect 502614 430128 502670 430137
rect 502614 430063 502670 430072
rect 502524 429140 502576 429146
rect 502524 429082 502576 429088
rect 502536 428233 502564 429082
rect 502522 428224 502578 428233
rect 502522 428159 502578 428168
rect 502706 427680 502762 427689
rect 502706 427615 502762 427624
rect 502720 427514 502748 427615
rect 502800 427576 502852 427582
rect 502800 427518 502852 427524
rect 502708 427508 502760 427514
rect 502708 427450 502760 427456
rect 502812 427417 502840 427518
rect 502798 427408 502854 427417
rect 502798 427343 502854 427352
rect 502904 425513 502932 436766
rect 502890 425504 502946 425513
rect 502890 425439 502946 425448
rect 502614 423328 502670 423337
rect 502614 423263 502670 423272
rect 502430 423056 502486 423065
rect 502430 422991 502486 423000
rect 501984 422266 502380 422294
rect 501984 390697 502012 422266
rect 501970 390688 502026 390697
rect 501970 390623 502026 390632
rect 501880 389972 501932 389978
rect 501880 389914 501932 389920
rect 502444 384305 502472 422991
rect 502522 422784 502578 422793
rect 502522 422719 502578 422728
rect 502536 386073 502564 422719
rect 502628 387025 502656 423263
rect 502706 422512 502762 422521
rect 502706 422447 502762 422456
rect 502614 387016 502670 387025
rect 502614 386951 502670 386960
rect 502522 386064 502578 386073
rect 502522 385999 502578 386008
rect 502430 384296 502486 384305
rect 502430 384231 502486 384240
rect 501788 383716 501840 383722
rect 501788 383658 501840 383664
rect 502720 383217 502748 422447
rect 502706 383208 502762 383217
rect 502706 383143 502762 383152
rect 502340 366444 502392 366450
rect 502340 366386 502392 366392
rect 502352 214713 502380 366386
rect 502432 365016 502484 365022
rect 502432 364958 502484 364964
rect 502444 220833 502472 364958
rect 502524 359508 502576 359514
rect 502524 359450 502576 359456
rect 502536 232937 502564 359450
rect 502708 356720 502760 356726
rect 502708 356662 502760 356668
rect 502616 349852 502668 349858
rect 502616 349794 502668 349800
rect 502522 232928 502578 232937
rect 502522 232863 502578 232872
rect 502628 226273 502656 349794
rect 502720 238377 502748 356662
rect 502800 251184 502852 251190
rect 502800 251126 502852 251132
rect 502812 250617 502840 251126
rect 502798 250608 502854 250617
rect 502798 250543 502854 250552
rect 502706 238368 502762 238377
rect 502706 238303 502762 238312
rect 502614 226264 502670 226273
rect 502614 226199 502670 226208
rect 502430 220824 502486 220833
rect 502430 220759 502486 220768
rect 502338 214704 502394 214713
rect 502338 214639 502394 214648
rect 501604 178628 501656 178634
rect 501604 178570 501656 178576
rect 502996 177410 503024 480226
rect 502984 177404 503036 177410
rect 502984 177346 503036 177352
rect 503088 177342 503116 481714
rect 503180 179994 503208 482258
rect 503272 481001 503300 523359
rect 503548 489914 503576 551103
rect 503720 546712 503772 546718
rect 503720 546654 503772 546660
rect 503732 546553 503760 546654
rect 503718 546544 503774 546553
rect 503718 546479 503774 546488
rect 503812 543176 503864 543182
rect 503812 543118 503864 543124
rect 503720 523388 503772 523394
rect 503720 523330 503772 523336
rect 503732 523161 503760 523330
rect 503718 523152 503774 523161
rect 503718 523087 503774 523096
rect 503720 519648 503772 519654
rect 503718 519616 503720 519625
rect 503772 519616 503774 519625
rect 503718 519551 503774 519560
rect 503364 489886 503576 489914
rect 503364 481817 503392 489886
rect 503628 488504 503680 488510
rect 503628 488446 503680 488452
rect 503640 487529 503668 488446
rect 503626 487520 503682 487529
rect 503626 487455 503682 487464
rect 503626 484392 503682 484401
rect 503626 484327 503682 484336
rect 503536 482996 503588 483002
rect 503536 482938 503588 482944
rect 503444 482384 503496 482390
rect 503444 482326 503496 482332
rect 503350 481808 503406 481817
rect 503350 481743 503406 481752
rect 503258 480992 503314 481001
rect 503258 480927 503314 480936
rect 503260 480888 503312 480894
rect 503260 480830 503312 480836
rect 503272 480254 503300 480830
rect 503272 480226 503392 480254
rect 503260 478916 503312 478922
rect 503260 478858 503312 478864
rect 503272 351490 503300 478858
rect 503364 390318 503392 480226
rect 503456 436830 503484 482326
rect 503548 481409 503576 482938
rect 503534 481400 503590 481409
rect 503534 481335 503590 481344
rect 503536 478168 503588 478174
rect 503536 478110 503588 478116
rect 503548 440366 503576 478110
rect 503640 451217 503668 484327
rect 503626 451208 503682 451217
rect 503626 451143 503682 451152
rect 503628 451104 503680 451110
rect 503626 451072 503628 451081
rect 503680 451072 503682 451081
rect 503626 451007 503682 451016
rect 503628 450968 503680 450974
rect 503628 450910 503680 450916
rect 503640 450809 503668 450910
rect 503626 450800 503682 450809
rect 503626 450735 503682 450744
rect 503628 449880 503680 449886
rect 503628 449822 503680 449828
rect 503640 449721 503668 449822
rect 503626 449712 503682 449721
rect 503626 449647 503682 449656
rect 503628 449608 503680 449614
rect 503628 449550 503680 449556
rect 503640 449449 503668 449550
rect 503626 449440 503682 449449
rect 503626 449375 503682 449384
rect 503628 448384 503680 448390
rect 503626 448352 503628 448361
rect 503680 448352 503682 448361
rect 503626 448287 503682 448296
rect 503628 445732 503680 445738
rect 503628 445674 503680 445680
rect 503640 445369 503668 445674
rect 503626 445360 503682 445369
rect 503626 445295 503682 445304
rect 503628 442944 503680 442950
rect 503628 442886 503680 442892
rect 503640 441833 503668 442886
rect 503626 441824 503682 441833
rect 503626 441759 503682 441768
rect 503628 441176 503680 441182
rect 503628 441118 503680 441124
rect 503640 440745 503668 441118
rect 503626 440736 503682 440745
rect 503626 440671 503682 440680
rect 503536 440360 503588 440366
rect 503536 440302 503588 440308
rect 503628 440224 503680 440230
rect 503626 440192 503628 440201
rect 503680 440192 503682 440201
rect 503626 440127 503682 440136
rect 503628 440088 503680 440094
rect 503628 440030 503680 440036
rect 503640 439929 503668 440030
rect 503626 439920 503682 439929
rect 503626 439855 503682 439864
rect 503536 438864 503588 438870
rect 503536 438806 503588 438812
rect 503548 437753 503576 438806
rect 503628 438796 503680 438802
rect 503628 438738 503680 438744
rect 503640 438025 503668 438738
rect 503626 438016 503682 438025
rect 503626 437951 503682 437960
rect 503534 437744 503590 437753
rect 503534 437679 503590 437688
rect 503628 437436 503680 437442
rect 503628 437378 503680 437384
rect 503640 437209 503668 437378
rect 503626 437200 503682 437209
rect 503626 437135 503682 437144
rect 503628 437096 503680 437102
rect 503628 437038 503680 437044
rect 503640 436937 503668 437038
rect 503626 436928 503682 436937
rect 503626 436863 503682 436872
rect 503444 436824 503496 436830
rect 503444 436766 503496 436772
rect 503628 436076 503680 436082
rect 503628 436018 503680 436024
rect 503444 436008 503496 436014
rect 503444 435950 503496 435956
rect 503456 434761 503484 435950
rect 503640 435577 503668 436018
rect 503626 435568 503682 435577
rect 503626 435503 503682 435512
rect 503442 434752 503498 434761
rect 503442 434687 503498 434696
rect 503536 434648 503588 434654
rect 503536 434590 503588 434596
rect 503444 434512 503496 434518
rect 503444 434454 503496 434460
rect 503456 433401 503484 434454
rect 503548 433945 503576 434590
rect 503628 434580 503680 434586
rect 503628 434522 503680 434528
rect 503640 434489 503668 434522
rect 503626 434480 503682 434489
rect 503626 434415 503682 434424
rect 503534 433936 503590 433945
rect 503534 433871 503590 433880
rect 503442 433392 503498 433401
rect 503442 433327 503498 433336
rect 503444 433220 503496 433226
rect 503444 433162 503496 433168
rect 503456 433129 503484 433162
rect 503536 433152 503588 433158
rect 503442 433120 503498 433129
rect 503536 433094 503588 433100
rect 503442 433055 503498 433064
rect 503444 433016 503496 433022
rect 503444 432958 503496 432964
rect 503456 432041 503484 432958
rect 503548 432585 503576 433094
rect 503628 433084 503680 433090
rect 503628 433026 503680 433032
rect 503534 432576 503590 432585
rect 503534 432511 503590 432520
rect 503640 432313 503668 433026
rect 503626 432304 503682 432313
rect 503626 432239 503682 432248
rect 503442 432032 503498 432041
rect 503442 431967 503498 431976
rect 503824 431954 503852 543118
rect 503904 542564 503956 542570
rect 503904 542506 503956 542512
rect 503916 433673 503944 542506
rect 504008 452985 504036 558214
rect 504454 554432 504510 554441
rect 504454 554367 504510 554376
rect 504178 536208 504234 536217
rect 504178 536143 504234 536152
rect 504086 533352 504142 533361
rect 504086 533287 504142 533296
rect 503994 452976 504050 452985
rect 503994 452911 504050 452920
rect 504100 439113 504128 533287
rect 504192 444009 504220 536143
rect 504272 520804 504324 520810
rect 504272 520746 504324 520752
rect 504178 444000 504234 444009
rect 504178 443935 504234 443944
rect 504086 439104 504142 439113
rect 504086 439039 504142 439048
rect 504284 438569 504312 520746
rect 504364 520600 504416 520606
rect 504364 520542 504416 520548
rect 504270 438560 504326 438569
rect 504270 438495 504326 438504
rect 504376 438297 504404 520542
rect 504468 479641 504496 554367
rect 504638 552800 504694 552809
rect 504638 552735 504694 552744
rect 504546 542328 504602 542337
rect 504546 542263 504602 542272
rect 504560 483177 504588 542263
rect 504652 520577 504680 552735
rect 504638 520568 504694 520577
rect 504638 520503 504694 520512
rect 504546 483168 504602 483177
rect 504546 483103 504602 483112
rect 504454 479632 504510 479641
rect 504454 479567 504510 479576
rect 504362 438288 504418 438297
rect 504362 438223 504418 438232
rect 503902 433664 503958 433673
rect 503902 433599 503958 433608
rect 503444 431928 503496 431934
rect 503444 431870 503496 431876
rect 503732 431926 503852 431954
rect 503456 431225 503484 431870
rect 503628 431792 503680 431798
rect 503626 431760 503628 431769
rect 503680 431760 503682 431769
rect 503536 431724 503588 431730
rect 503626 431695 503682 431704
rect 503536 431666 503588 431672
rect 503548 431497 503576 431666
rect 503534 431488 503590 431497
rect 503534 431423 503590 431432
rect 503442 431216 503498 431225
rect 503442 431151 503498 431160
rect 503628 430500 503680 430506
rect 503628 430442 503680 430448
rect 503444 430432 503496 430438
rect 503640 430409 503668 430442
rect 503444 430374 503496 430380
rect 503626 430400 503682 430409
rect 503456 429321 503484 430374
rect 503536 430364 503588 430370
rect 503626 430335 503682 430344
rect 503536 430306 503588 430312
rect 503548 429593 503576 430306
rect 503626 429992 503682 430001
rect 503732 429978 503760 431926
rect 503682 429950 503760 429978
rect 503626 429927 503682 429936
rect 503534 429584 503590 429593
rect 503534 429519 503590 429528
rect 503442 429312 503498 429321
rect 503442 429247 503498 429256
rect 503628 429072 503680 429078
rect 503626 429040 503628 429049
rect 503680 429040 503682 429049
rect 503626 428975 503682 428984
rect 503628 428868 503680 428874
rect 503628 428810 503680 428816
rect 503640 428777 503668 428810
rect 503626 428768 503682 428777
rect 503626 428703 503682 428712
rect 503628 428664 503680 428670
rect 503628 428606 503680 428612
rect 503640 428505 503668 428606
rect 503626 428496 503682 428505
rect 503626 428431 503682 428440
rect 503628 428392 503680 428398
rect 503628 428334 503680 428340
rect 503640 427961 503668 428334
rect 503626 427952 503682 427961
rect 503626 427887 503682 427896
rect 503444 427780 503496 427786
rect 503444 427722 503496 427728
rect 503456 426873 503484 427722
rect 503536 427712 503588 427718
rect 503536 427654 503588 427660
rect 503442 426864 503498 426873
rect 503442 426799 503498 426808
rect 503548 426601 503576 427654
rect 503628 427644 503680 427650
rect 503628 427586 503680 427592
rect 503640 427145 503668 427586
rect 503626 427136 503682 427145
rect 503626 427071 503682 427080
rect 503534 426592 503590 426601
rect 503534 426527 503590 426536
rect 503444 426420 503496 426426
rect 503444 426362 503496 426368
rect 503456 425785 503484 426362
rect 503628 426352 503680 426358
rect 503626 426320 503628 426329
rect 503680 426320 503682 426329
rect 503536 426284 503588 426290
rect 503626 426255 503682 426264
rect 503536 426226 503588 426232
rect 503442 425776 503498 425785
rect 503442 425711 503498 425720
rect 503548 425241 503576 426226
rect 503534 425232 503590 425241
rect 503534 425167 503590 425176
rect 503628 425060 503680 425066
rect 503628 425002 503680 425008
rect 503444 424992 503496 424998
rect 503640 424969 503668 425002
rect 503444 424934 503496 424940
rect 503626 424960 503682 424969
rect 503456 423881 503484 424934
rect 503536 424924 503588 424930
rect 503626 424895 503682 424904
rect 503536 424866 503588 424872
rect 503548 424153 503576 424866
rect 503628 424856 503680 424862
rect 503628 424798 503680 424804
rect 503640 424425 503668 424798
rect 503626 424416 503682 424425
rect 503626 424351 503682 424360
rect 503534 424144 503590 424153
rect 503534 424079 503590 424088
rect 503442 423872 503498 423881
rect 503442 423807 503498 423816
rect 503628 423632 503680 423638
rect 503626 423600 503628 423609
rect 503680 423600 503682 423609
rect 503626 423535 503682 423544
rect 503352 390312 503404 390318
rect 503352 390254 503404 390260
rect 504744 373697 504772 586486
rect 505112 387705 505140 599519
rect 505940 598097 505968 600100
rect 507320 598097 507348 600100
rect 505926 598088 505982 598097
rect 505926 598023 505982 598032
rect 507306 598088 507362 598097
rect 507306 598023 507362 598032
rect 507860 555484 507912 555490
rect 507860 555426 507912 555432
rect 507872 554849 507900 555426
rect 507858 554840 507914 554849
rect 507858 554775 507914 554784
rect 507400 551472 507452 551478
rect 507400 551414 507452 551420
rect 506572 550044 506624 550050
rect 506572 549986 506624 549992
rect 505376 548752 505428 548758
rect 505376 548694 505428 548700
rect 505192 524816 505244 524822
rect 505192 524758 505244 524764
rect 505098 387696 505154 387705
rect 505098 387631 505154 387640
rect 504730 373688 504786 373697
rect 504730 373623 504786 373632
rect 505100 363656 505152 363662
rect 505100 363598 505152 363604
rect 503904 362228 503956 362234
rect 503904 362170 503956 362176
rect 503812 360868 503864 360874
rect 503812 360810 503864 360816
rect 503260 351484 503312 351490
rect 503260 351426 503312 351432
rect 503720 351212 503772 351218
rect 503720 351154 503772 351160
rect 503628 346384 503680 346390
rect 503628 346326 503680 346332
rect 503640 346089 503668 346326
rect 503626 346080 503682 346089
rect 503626 346015 503682 346024
rect 503628 340876 503680 340882
rect 503628 340818 503680 340824
rect 503640 340377 503668 340818
rect 503626 340368 503682 340377
rect 503626 340303 503682 340312
rect 503628 333940 503680 333946
rect 503628 333882 503680 333888
rect 503640 333849 503668 333882
rect 503626 333840 503682 333849
rect 503626 333775 503682 333784
rect 503628 328432 503680 328438
rect 503628 328374 503680 328380
rect 503640 328137 503668 328374
rect 503626 328128 503682 328137
rect 503626 328063 503682 328072
rect 503628 322924 503680 322930
rect 503628 322866 503680 322872
rect 503640 322425 503668 322866
rect 503626 322416 503682 322425
rect 503626 322351 503682 322360
rect 503628 304972 503680 304978
rect 503628 304914 503680 304920
rect 503640 304473 503668 304914
rect 503626 304464 503682 304473
rect 503626 304399 503682 304408
rect 503628 298104 503680 298110
rect 503628 298046 503680 298052
rect 503640 297945 503668 298046
rect 503626 297936 503682 297945
rect 503626 297871 503682 297880
rect 503628 292528 503680 292534
rect 503628 292470 503680 292476
rect 503640 292233 503668 292470
rect 503626 292224 503682 292233
rect 503626 292159 503682 292168
rect 503628 287020 503680 287026
rect 503628 286962 503680 286968
rect 503640 286521 503668 286962
rect 503626 286512 503682 286521
rect 503626 286447 503682 286456
rect 503628 274644 503680 274650
rect 503628 274586 503680 274592
rect 503640 274281 503668 274586
rect 503626 274272 503682 274281
rect 503626 274207 503682 274216
rect 503626 184920 503682 184929
rect 503732 184906 503760 351154
rect 503824 244361 503852 360810
rect 503916 256737 503944 362170
rect 503902 256728 503958 256737
rect 503902 256663 503958 256672
rect 505112 251190 505140 363598
rect 505100 251184 505152 251190
rect 505100 251126 505152 251132
rect 503810 244352 503866 244361
rect 503810 244287 503866 244296
rect 503682 184878 503760 184906
rect 503626 184855 503682 184864
rect 503168 179988 503220 179994
rect 503168 179930 503220 179936
rect 503076 177336 503128 177342
rect 503076 177278 503128 177284
rect 505204 175234 505232 524758
rect 505284 522708 505336 522714
rect 505284 522650 505336 522656
rect 505296 176458 505324 522650
rect 505388 431458 505416 548694
rect 506480 548004 506532 548010
rect 506480 547946 506532 547952
rect 506492 547913 506520 547946
rect 506478 547904 506534 547913
rect 506478 547839 506534 547848
rect 506478 541104 506534 541113
rect 506478 541039 506480 541048
rect 506532 541039 506534 541048
rect 506480 541010 506532 541016
rect 505560 537668 505612 537674
rect 505560 537610 505612 537616
rect 505468 533452 505520 533458
rect 505468 533394 505520 533400
rect 505376 431452 505428 431458
rect 505376 431394 505428 431400
rect 505480 429146 505508 533394
rect 505572 433294 505600 537610
rect 505744 534812 505796 534818
rect 505744 534754 505796 534760
rect 505652 533588 505704 533594
rect 505652 533530 505704 533536
rect 505560 433288 505612 433294
rect 505560 433230 505612 433236
rect 505664 430574 505692 533530
rect 505756 431322 505784 534754
rect 505928 528692 505980 528698
rect 505928 528634 505980 528640
rect 505836 523660 505888 523666
rect 505836 523602 505888 523608
rect 505848 483002 505876 523602
rect 505940 520946 505968 528634
rect 505928 520940 505980 520946
rect 505928 520882 505980 520888
rect 506020 520192 506072 520198
rect 506020 520134 506072 520140
rect 505928 520124 505980 520130
rect 505928 520066 505980 520072
rect 505940 484401 505968 520066
rect 506032 519761 506060 520134
rect 506018 519752 506074 519761
rect 506018 519687 506074 519696
rect 505926 484392 505982 484401
rect 505926 484327 505982 484336
rect 505836 482996 505888 483002
rect 505836 482938 505888 482944
rect 505834 480312 505890 480321
rect 505834 480247 505890 480256
rect 505744 431316 505796 431322
rect 505744 431258 505796 431264
rect 505652 430568 505704 430574
rect 505652 430510 505704 430516
rect 505468 429140 505520 429146
rect 505468 429082 505520 429088
rect 505374 394632 505430 394641
rect 505374 394567 505430 394576
rect 505388 390425 505416 394567
rect 505374 390416 505430 390425
rect 505374 390351 505430 390360
rect 505848 388958 505876 480247
rect 506584 434722 506612 549986
rect 506664 544536 506716 544542
rect 506664 544478 506716 544484
rect 506572 434716 506624 434722
rect 506572 434658 506624 434664
rect 506676 433022 506704 544478
rect 506756 541272 506808 541278
rect 506756 541214 506808 541220
rect 506768 433158 506796 541214
rect 507030 540016 507086 540025
rect 507030 539951 507086 539960
rect 506848 538960 506900 538966
rect 506848 538902 506900 538908
rect 506860 433226 506888 538902
rect 506940 534880 506992 534886
rect 506940 534822 506992 534828
rect 506952 436014 506980 534822
rect 507044 445097 507072 539951
rect 507306 530496 507362 530505
rect 507306 530431 507362 530440
rect 507122 525056 507178 525065
rect 507122 524991 507178 525000
rect 507136 445913 507164 524991
rect 507216 524544 507268 524550
rect 507216 524486 507268 524492
rect 507228 450974 507256 524486
rect 507320 472297 507348 530431
rect 507306 472288 507362 472297
rect 507306 472223 507362 472232
rect 507216 450968 507268 450974
rect 507216 450910 507268 450916
rect 507122 445904 507178 445913
rect 507122 445839 507178 445848
rect 507030 445088 507086 445097
rect 507030 445023 507086 445032
rect 506940 436008 506992 436014
rect 506940 435950 506992 435956
rect 506848 433220 506900 433226
rect 506848 433162 506900 433168
rect 506756 433152 506808 433158
rect 506756 433094 506808 433100
rect 507412 433090 507440 551414
rect 508044 551336 508096 551342
rect 508044 551278 508096 551284
rect 507860 531616 507912 531622
rect 507860 531558 507912 531564
rect 507400 433084 507452 433090
rect 507400 433026 507452 433032
rect 506664 433016 506716 433022
rect 506664 432958 506716 432964
rect 505836 388952 505888 388958
rect 505836 388894 505888 388900
rect 507872 177818 507900 531558
rect 507952 520260 508004 520266
rect 507952 520202 508004 520208
rect 507964 519761 507992 520202
rect 507950 519752 508006 519761
rect 507950 519687 508006 519696
rect 507950 519072 508006 519081
rect 507950 519007 508006 519016
rect 507964 381721 507992 519007
rect 508056 428670 508084 551278
rect 508136 547256 508188 547262
rect 508136 547198 508188 547204
rect 508044 428664 508096 428670
rect 508044 428606 508096 428612
rect 508148 427582 508176 547198
rect 508228 540388 508280 540394
rect 508228 540330 508280 540336
rect 508240 428398 508268 540330
rect 508410 539064 508466 539073
rect 508410 538999 508466 539008
rect 508320 536104 508372 536110
rect 508320 536046 508372 536052
rect 508228 428392 508280 428398
rect 508228 428334 508280 428340
rect 508136 427576 508188 427582
rect 508136 427518 508188 427524
rect 508332 427514 508360 536046
rect 508424 447273 508452 538999
rect 508504 528012 508556 528018
rect 508504 527954 508556 527960
rect 508410 447264 508466 447273
rect 508410 447199 508466 447208
rect 508516 441182 508544 527954
rect 508596 521756 508648 521762
rect 508596 521698 508648 521704
rect 508608 482458 508636 521698
rect 508596 482452 508648 482458
rect 508596 482394 508648 482400
rect 508504 441176 508556 441182
rect 508504 441118 508556 441124
rect 508320 427508 508372 427514
rect 508320 427450 508372 427456
rect 508502 407824 508558 407833
rect 508502 407759 508558 407768
rect 508516 394641 508544 407759
rect 508502 394632 508558 394641
rect 508502 394567 508558 394576
rect 507950 381712 508006 381721
rect 507950 381647 508006 381656
rect 508700 354113 508728 600100
rect 509976 556232 510028 556238
rect 509976 556174 510028 556180
rect 509698 552936 509754 552945
rect 509698 552871 509754 552880
rect 509606 551304 509662 551313
rect 509606 551239 509662 551248
rect 509238 550760 509294 550769
rect 509238 550695 509294 550704
rect 509252 550662 509280 550695
rect 509240 550656 509292 550662
rect 509240 550598 509292 550604
rect 509240 520124 509292 520130
rect 509240 520066 509292 520072
rect 508686 354104 508742 354113
rect 508686 354039 508742 354048
rect 507860 177812 507912 177818
rect 507860 177754 507912 177760
rect 505284 176452 505336 176458
rect 505284 176394 505336 176400
rect 509252 176322 509280 520066
rect 509516 519648 509568 519654
rect 509516 519590 509568 519596
rect 509422 519208 509478 519217
rect 509422 519143 509478 519152
rect 509332 512644 509384 512650
rect 509332 512586 509384 512592
rect 509344 177886 509372 512586
rect 509436 382945 509464 519143
rect 509528 388482 509556 519590
rect 509620 441017 509648 551239
rect 509712 477193 509740 552871
rect 509792 533044 509844 533050
rect 509792 532986 509844 532992
rect 509804 532817 509832 532986
rect 509790 532808 509846 532817
rect 509790 532743 509846 532752
rect 509792 529304 509844 529310
rect 509792 529246 509844 529252
rect 509698 477184 509754 477193
rect 509698 477119 509754 477128
rect 509804 455122 509832 529246
rect 509884 524612 509936 524618
rect 509884 524554 509936 524560
rect 509896 481778 509924 524554
rect 509988 513505 510016 556174
rect 509974 513496 510030 513505
rect 509974 513431 510030 513440
rect 509884 481772 509936 481778
rect 509884 481714 509936 481720
rect 509792 455116 509844 455122
rect 509792 455058 509844 455064
rect 509606 441008 509662 441017
rect 509606 440943 509662 440952
rect 509516 388476 509568 388482
rect 509516 388418 509568 388424
rect 509422 382936 509478 382945
rect 509422 382871 509478 382880
rect 510080 351354 510108 600100
rect 510160 554804 510212 554810
rect 510160 554746 510212 554752
rect 510172 523666 510200 554746
rect 510252 528760 510304 528766
rect 510252 528702 510304 528708
rect 510160 523660 510212 523666
rect 510160 523602 510212 523608
rect 510264 521626 510292 528702
rect 510252 521620 510304 521626
rect 510252 521562 510304 521568
rect 510356 518894 510384 600170
rect 524052 600160 524104 600166
rect 524052 600102 524104 600108
rect 510804 550112 510856 550118
rect 510804 550054 510856 550060
rect 510620 525972 510672 525978
rect 510620 525914 510672 525920
rect 510632 520010 510660 525914
rect 510540 519982 510660 520010
rect 510540 519194 510568 519982
rect 510620 519920 510672 519926
rect 510620 519862 510672 519868
rect 510632 519353 510660 519862
rect 510710 519752 510766 519761
rect 510710 519687 510766 519696
rect 510618 519344 510674 519353
rect 510618 519279 510674 519288
rect 510540 519166 510660 519194
rect 510356 518866 510568 518894
rect 510540 511970 510568 518866
rect 510528 511964 510580 511970
rect 510528 511906 510580 511912
rect 510540 511290 510568 511906
rect 510528 511284 510580 511290
rect 510528 511226 510580 511232
rect 510068 351348 510120 351354
rect 510068 351290 510120 351296
rect 510632 177954 510660 519166
rect 510724 389881 510752 519687
rect 510816 440094 510844 550054
rect 510894 548720 510950 548729
rect 510894 548655 510950 548664
rect 510908 440473 510936 548655
rect 510986 547224 511042 547233
rect 510986 547159 511042 547168
rect 511000 441289 511028 547159
rect 511172 542632 511224 542638
rect 511172 542574 511224 542580
rect 511080 529440 511132 529446
rect 511080 529382 511132 529388
rect 510986 441280 511042 441289
rect 510986 441215 511042 441224
rect 510894 440464 510950 440473
rect 510894 440399 510950 440408
rect 510804 440088 510856 440094
rect 510804 440030 510856 440036
rect 511092 437102 511120 529382
rect 511184 488510 511212 542574
rect 511264 523660 511316 523666
rect 511264 523602 511316 523608
rect 511172 488504 511224 488510
rect 511172 488446 511224 488452
rect 511276 478922 511304 523602
rect 511460 510066 511488 600100
rect 512840 598330 512868 600100
rect 512828 598324 512880 598330
rect 512828 598266 512880 598272
rect 514220 598262 514248 600100
rect 515600 598874 515628 600100
rect 515588 598868 515640 598874
rect 515588 598810 515640 598816
rect 514208 598256 514260 598262
rect 514208 598198 514260 598204
rect 514852 559564 514904 559570
rect 514852 559506 514904 559512
rect 511998 559056 512054 559065
rect 511998 558991 512000 559000
rect 512052 558991 512054 559000
rect 512000 558962 512052 558968
rect 512184 558204 512236 558210
rect 512184 558146 512236 558152
rect 512090 545320 512146 545329
rect 512090 545255 512146 545264
rect 511540 537056 511592 537062
rect 511540 536998 511592 537004
rect 511552 519761 511580 536998
rect 512000 527400 512052 527406
rect 512000 527342 512052 527348
rect 512012 527241 512040 527342
rect 511998 527232 512054 527241
rect 511998 527167 512054 527176
rect 512000 525632 512052 525638
rect 512000 525574 512052 525580
rect 512012 524521 512040 525574
rect 511998 524512 512054 524521
rect 511998 524447 512054 524456
rect 511630 520568 511686 520577
rect 511630 520503 511686 520512
rect 511538 519752 511594 519761
rect 511538 519687 511594 519696
rect 511644 518894 511672 520503
rect 511552 518866 511672 518894
rect 511448 510060 511500 510066
rect 511448 510002 511500 510008
rect 511552 507226 511580 518866
rect 511632 510060 511684 510066
rect 511632 510002 511684 510008
rect 511368 507198 511580 507226
rect 511368 485353 511396 507198
rect 511644 502334 511672 510002
rect 511460 502306 511672 502334
rect 511354 485344 511410 485353
rect 511354 485279 511410 485288
rect 511354 481400 511410 481409
rect 511354 481335 511410 481344
rect 511264 478916 511316 478922
rect 511264 478858 511316 478864
rect 511080 437096 511132 437102
rect 511080 437038 511132 437044
rect 510710 389872 510766 389881
rect 510710 389807 510766 389816
rect 510620 177948 510672 177954
rect 510620 177890 510672 177896
rect 509332 177880 509384 177886
rect 509332 177822 509384 177828
rect 509240 176316 509292 176322
rect 509240 176258 509292 176264
rect 505192 175228 505244 175234
rect 505192 175170 505244 175176
rect 511368 175030 511396 481335
rect 511460 373998 511488 502306
rect 512104 439385 512132 545255
rect 512196 455190 512224 558146
rect 513564 553444 513616 553450
rect 513564 553386 513616 553392
rect 512920 552084 512972 552090
rect 512920 552026 512972 552032
rect 512274 544776 512330 544785
rect 512274 544711 512330 544720
rect 512184 455184 512236 455190
rect 512184 455126 512236 455132
rect 512288 446729 512316 544711
rect 512458 540288 512514 540297
rect 512458 540223 512514 540232
rect 512366 532672 512422 532681
rect 512366 532607 512422 532616
rect 512274 446720 512330 446729
rect 512274 446655 512330 446664
rect 512090 439376 512146 439385
rect 512090 439311 512146 439320
rect 512380 437481 512408 532607
rect 512472 445641 512500 540223
rect 512550 537568 512606 537577
rect 512550 537503 512606 537512
rect 512564 447001 512592 537503
rect 512734 534848 512790 534857
rect 512734 534783 512790 534792
rect 512642 519072 512698 519081
rect 512642 519007 512698 519016
rect 512656 486169 512684 519007
rect 512642 486160 512698 486169
rect 512642 486095 512698 486104
rect 512642 480856 512698 480865
rect 512642 480791 512698 480800
rect 512550 446992 512606 447001
rect 512550 446927 512606 446936
rect 512458 445632 512514 445641
rect 512458 445567 512514 445576
rect 512366 437472 512422 437481
rect 512366 437407 512422 437416
rect 511448 373992 511500 373998
rect 511448 373934 511500 373940
rect 511356 175024 511408 175030
rect 511356 174966 511408 174972
rect 512656 174962 512684 480791
rect 512748 446457 512776 534783
rect 512828 531412 512880 531418
rect 512828 531354 512880 531360
rect 512840 451042 512868 531354
rect 512828 451036 512880 451042
rect 512828 450978 512880 450984
rect 512734 446448 512790 446457
rect 512734 446383 512790 446392
rect 512932 440230 512960 552026
rect 513380 522640 513432 522646
rect 513380 522582 513432 522588
rect 512920 440224 512972 440230
rect 512920 440166 512972 440172
rect 513392 176662 513420 522582
rect 513472 521620 513524 521626
rect 513472 521562 513524 521568
rect 513484 180130 513512 521562
rect 513576 448322 513604 553386
rect 513840 534744 513892 534750
rect 513840 534686 513892 534692
rect 513748 533384 513800 533390
rect 513748 533326 513800 533332
rect 513656 526516 513708 526522
rect 513656 526458 513708 526464
rect 513564 448316 513616 448322
rect 513564 448258 513616 448264
rect 513668 424862 513696 526458
rect 513760 451110 513788 533326
rect 513852 452402 513880 534686
rect 513932 533112 513984 533118
rect 513932 533054 513984 533060
rect 513944 456550 513972 533054
rect 514760 532840 514812 532846
rect 514758 532808 514760 532817
rect 514812 532808 514814 532817
rect 514758 532743 514814 532752
rect 514022 529136 514078 529145
rect 514022 529071 514078 529080
rect 514036 457609 514064 529071
rect 514760 527332 514812 527338
rect 514760 527274 514812 527280
rect 514772 527241 514800 527274
rect 514758 527232 514814 527241
rect 514758 527167 514814 527176
rect 514206 525872 514262 525881
rect 514206 525807 514262 525816
rect 514114 519888 514170 519897
rect 514114 519823 514170 519832
rect 514128 476105 514156 519823
rect 514220 485625 514248 525807
rect 514760 521552 514812 521558
rect 514760 521494 514812 521500
rect 514772 520305 514800 521494
rect 514758 520296 514814 520305
rect 514758 520231 514814 520240
rect 514666 514720 514722 514729
rect 514666 514655 514722 514664
rect 514680 505345 514708 514655
rect 514666 505336 514722 505345
rect 514666 505271 514722 505280
rect 514206 485616 514262 485625
rect 514206 485551 514262 485560
rect 514114 476096 514170 476105
rect 514114 476031 514170 476040
rect 514022 457600 514078 457609
rect 514022 457535 514078 457544
rect 513932 456544 513984 456550
rect 513932 456486 513984 456492
rect 514864 453898 514892 559506
rect 515402 558376 515458 558385
rect 515402 558311 515458 558320
rect 514944 549908 514996 549914
rect 514944 549850 514996 549856
rect 514852 453892 514904 453898
rect 514852 453834 514904 453840
rect 514956 452470 514984 549850
rect 515128 544400 515180 544406
rect 515128 544342 515180 544348
rect 515036 520736 515088 520742
rect 515036 520678 515088 520684
rect 514944 452464 514996 452470
rect 514944 452406 514996 452412
rect 513840 452396 513892 452402
rect 513840 452338 513892 452344
rect 513748 451104 513800 451110
rect 513748 451046 513800 451052
rect 515048 426290 515076 520678
rect 515140 452538 515168 544342
rect 515312 540320 515364 540326
rect 515312 540262 515364 540268
rect 515220 526108 515272 526114
rect 515220 526050 515272 526056
rect 515128 452532 515180 452538
rect 515128 452474 515180 452480
rect 515232 437442 515260 526050
rect 515324 452606 515352 540262
rect 515416 471481 515444 558311
rect 515494 555520 515550 555529
rect 515494 555455 515550 555464
rect 515402 471472 515458 471481
rect 515402 471407 515458 471416
rect 515508 471209 515536 555455
rect 516600 541204 516652 541210
rect 516600 541146 516652 541152
rect 516508 541000 516560 541006
rect 516508 540942 516560 540948
rect 516140 538348 516192 538354
rect 516140 538290 516192 538296
rect 515678 534984 515734 534993
rect 515678 534919 515734 534928
rect 515588 523932 515640 523938
rect 515588 523874 515640 523880
rect 515600 482390 515628 523874
rect 515588 482384 515640 482390
rect 515588 482326 515640 482332
rect 515494 471200 515550 471209
rect 515494 471135 515550 471144
rect 515312 452600 515364 452606
rect 515312 452542 515364 452548
rect 515220 437436 515272 437442
rect 515220 437378 515272 437384
rect 515036 426284 515088 426290
rect 515036 426226 515088 426232
rect 515692 426057 515720 534919
rect 515678 426048 515734 426057
rect 515678 425983 515734 425992
rect 513656 424856 513708 424862
rect 513656 424798 513708 424804
rect 513472 180124 513524 180130
rect 513472 180066 513524 180072
rect 513380 176656 513432 176662
rect 513380 176598 513432 176604
rect 516152 176390 516180 538290
rect 516232 530120 516284 530126
rect 516232 530062 516284 530068
rect 516244 177614 516272 530062
rect 516324 525836 516376 525842
rect 516324 525778 516376 525784
rect 516336 274650 516364 525778
rect 516416 520328 516468 520334
rect 516416 520270 516468 520276
rect 516428 298110 516456 520270
rect 516520 333946 516548 540942
rect 516612 448390 516640 541146
rect 516690 530904 516746 530913
rect 516690 530839 516746 530848
rect 516704 456249 516732 530839
rect 516876 523252 516928 523258
rect 516876 523194 516928 523200
rect 516784 522504 516836 522510
rect 516784 522446 516836 522452
rect 516796 463486 516824 522446
rect 516888 482322 516916 523194
rect 516876 482316 516928 482322
rect 516876 482258 516928 482264
rect 516784 463480 516836 463486
rect 516784 463422 516836 463428
rect 516690 456240 516746 456249
rect 516690 456175 516746 456184
rect 516600 448384 516652 448390
rect 516600 448326 516652 448332
rect 516980 364993 517008 600100
rect 518360 598806 518388 600100
rect 519740 598942 519768 600100
rect 519728 598936 519780 598942
rect 519728 598878 519780 598884
rect 518348 598800 518400 598806
rect 518348 598742 518400 598748
rect 521120 597582 521148 600100
rect 518164 597576 518216 597582
rect 518164 597518 518216 597524
rect 521108 597576 521160 597582
rect 521108 597518 521160 597524
rect 517704 542496 517756 542502
rect 517704 542438 517756 542444
rect 517060 534132 517112 534138
rect 517060 534074 517112 534080
rect 517072 521257 517100 534074
rect 517612 531684 517664 531690
rect 517612 531626 517664 531632
rect 517520 527876 517572 527882
rect 517520 527818 517572 527824
rect 517532 527241 517560 527818
rect 517518 527232 517574 527241
rect 517518 527167 517574 527176
rect 517520 526720 517572 526726
rect 517520 526662 517572 526668
rect 517532 522306 517560 526662
rect 517520 522300 517572 522306
rect 517520 522242 517572 522248
rect 517520 522028 517572 522034
rect 517520 521970 517572 521976
rect 517532 521801 517560 521970
rect 517518 521792 517574 521801
rect 517518 521727 517574 521736
rect 517058 521248 517114 521257
rect 517058 521183 517114 521192
rect 516966 364984 517022 364993
rect 516966 364919 517022 364928
rect 516508 333940 516560 333946
rect 516508 333882 516560 333888
rect 516416 298104 516468 298110
rect 516416 298046 516468 298052
rect 516324 274644 516376 274650
rect 516324 274586 516376 274592
rect 516232 177608 516284 177614
rect 516232 177550 516284 177556
rect 517624 177478 517652 531626
rect 517716 483682 517744 542438
rect 517796 542428 517848 542434
rect 517796 542370 517848 542376
rect 517704 483676 517756 483682
rect 517704 483618 517756 483624
rect 517704 482452 517756 482458
rect 517704 482394 517756 482400
rect 517612 177472 517664 177478
rect 517612 177414 517664 177420
rect 516140 176384 516192 176390
rect 516140 176326 516192 176332
rect 517716 175166 517744 482394
rect 517808 328438 517836 542370
rect 517980 541748 518032 541754
rect 517980 541690 518032 541696
rect 517886 536072 517942 536081
rect 517886 536007 517942 536016
rect 517900 424697 517928 536007
rect 517992 449614 518020 541690
rect 518070 523152 518126 523161
rect 518070 523087 518126 523096
rect 518084 523054 518112 523087
rect 518072 523048 518124 523054
rect 518072 522990 518124 522996
rect 518072 522844 518124 522850
rect 518072 522786 518124 522792
rect 518084 457978 518112 522786
rect 518072 457972 518124 457978
rect 518072 457914 518124 457920
rect 517980 449608 518032 449614
rect 517980 449550 518032 449556
rect 517886 424688 517942 424697
rect 517886 424623 517942 424632
rect 518176 379001 518204 597518
rect 520740 558952 520792 558958
rect 520740 558894 520792 558900
rect 519360 552696 519412 552702
rect 519360 552638 519412 552644
rect 518900 550792 518952 550798
rect 518900 550734 518952 550740
rect 518440 537124 518492 537130
rect 518440 537066 518492 537072
rect 518254 533760 518310 533769
rect 518254 533695 518310 533704
rect 518268 526561 518296 533695
rect 518254 526552 518310 526561
rect 518254 526487 518310 526496
rect 518346 521520 518402 521529
rect 518346 521455 518402 521464
rect 518256 521144 518308 521150
rect 518256 521086 518308 521092
rect 518268 463554 518296 521086
rect 518360 469577 518388 521455
rect 518346 469568 518402 469577
rect 518346 469503 518402 469512
rect 518256 463548 518308 463554
rect 518256 463490 518308 463496
rect 518162 378992 518218 379001
rect 518162 378927 518218 378936
rect 517796 328432 517848 328438
rect 517796 328374 517848 328380
rect 518452 177750 518480 537066
rect 518440 177744 518492 177750
rect 518440 177686 518492 177692
rect 518912 177206 518940 550734
rect 519176 535492 519228 535498
rect 519176 535434 519228 535440
rect 519084 532976 519136 532982
rect 519084 532918 519136 532924
rect 518990 532808 519046 532817
rect 518990 532743 518992 532752
rect 519044 532743 519046 532752
rect 518992 532714 519044 532720
rect 519096 528554 519124 532918
rect 519004 528526 519124 528554
rect 519004 177546 519032 528526
rect 519084 525904 519136 525910
rect 519084 525846 519136 525852
rect 519096 178906 519124 525846
rect 519188 292534 519216 535434
rect 519268 524476 519320 524482
rect 519268 524418 519320 524424
rect 519280 304978 519308 524418
rect 519372 427650 519400 552638
rect 520648 547936 520700 547942
rect 520648 547878 520700 547884
rect 520556 546508 520608 546514
rect 520556 546450 520608 546456
rect 519450 543144 519506 543153
rect 519450 543079 519506 543088
rect 519464 444281 519492 543079
rect 520464 536852 520516 536858
rect 520464 536794 520516 536800
rect 520280 535696 520332 535702
rect 520280 535638 520332 535644
rect 519542 526416 519598 526425
rect 519542 526351 519598 526360
rect 519556 446185 519584 526351
rect 519636 525428 519688 525434
rect 519636 525370 519688 525376
rect 519648 453966 519676 525370
rect 519726 523560 519782 523569
rect 519726 523495 519782 523504
rect 519740 464409 519768 523495
rect 519726 464400 519782 464409
rect 519726 464335 519782 464344
rect 519636 453960 519688 453966
rect 519636 453902 519688 453908
rect 519542 446176 519598 446185
rect 519542 446111 519598 446120
rect 519450 444272 519506 444281
rect 519450 444207 519506 444216
rect 519360 427644 519412 427650
rect 519360 427586 519412 427592
rect 519268 304972 519320 304978
rect 519268 304914 519320 304920
rect 519176 292528 519228 292534
rect 519176 292470 519228 292476
rect 519084 178900 519136 178906
rect 519084 178842 519136 178848
rect 520292 177682 520320 535638
rect 520372 520940 520424 520946
rect 520372 520882 520424 520888
rect 520384 178974 520412 520882
rect 520476 287026 520504 536794
rect 520568 322930 520596 546450
rect 520660 340882 520688 547878
rect 520752 451178 520780 558894
rect 521936 558340 521988 558346
rect 521936 558282 521988 558288
rect 521660 539776 521712 539782
rect 521658 539744 521660 539753
rect 521712 539744 521714 539753
rect 521658 539679 521714 539688
rect 521660 539640 521712 539646
rect 521658 539608 521660 539617
rect 521712 539608 521714 539617
rect 521658 539543 521714 539552
rect 521106 535120 521162 535129
rect 521106 535055 521162 535064
rect 520924 528352 520976 528358
rect 520924 528294 520976 528300
rect 520830 522744 520886 522753
rect 520830 522679 520886 522688
rect 520740 451172 520792 451178
rect 520740 451114 520792 451120
rect 520844 435849 520872 522679
rect 520936 465050 520964 528294
rect 521016 522436 521068 522442
rect 521016 522378 521068 522384
rect 520924 465044 520976 465050
rect 520924 464986 520976 464992
rect 521028 462058 521056 522378
rect 521120 485081 521148 535055
rect 521660 531752 521712 531758
rect 521660 531694 521712 531700
rect 521672 531457 521700 531694
rect 521658 531448 521714 531457
rect 521658 531383 521714 531392
rect 521752 530324 521804 530330
rect 521752 530266 521804 530272
rect 521106 485072 521162 485081
rect 521106 485007 521162 485016
rect 521016 462052 521068 462058
rect 521016 461994 521068 462000
rect 520830 435840 520886 435849
rect 520830 435775 520886 435784
rect 520648 340876 520700 340882
rect 520648 340818 520700 340824
rect 520556 322924 520608 322930
rect 520556 322866 520608 322872
rect 520464 287020 520516 287026
rect 520464 286962 520516 286968
rect 520372 178968 520424 178974
rect 520372 178910 520424 178916
rect 521764 178770 521792 530266
rect 521844 520532 521896 520538
rect 521844 520474 521896 520480
rect 521856 180470 521884 520474
rect 521948 431798 521976 558282
rect 522302 539336 522358 539345
rect 522302 539271 522358 539280
rect 522026 538792 522082 538801
rect 522026 538727 522082 538736
rect 522040 439657 522068 538727
rect 522120 523456 522172 523462
rect 522120 523398 522172 523404
rect 522132 455258 522160 523398
rect 522212 522572 522264 522578
rect 522212 522514 522264 522520
rect 522224 459338 522252 522514
rect 522316 475561 522344 539271
rect 522396 526448 522448 526454
rect 522396 526390 522448 526396
rect 522302 475552 522358 475561
rect 522302 475487 522358 475496
rect 522408 469130 522436 526390
rect 522396 469124 522448 469130
rect 522396 469066 522448 469072
rect 522212 459332 522264 459338
rect 522212 459274 522264 459280
rect 522120 455252 522172 455258
rect 522120 455194 522172 455200
rect 522026 439648 522082 439657
rect 522026 439583 522082 439592
rect 521936 431792 521988 431798
rect 521936 431734 521988 431740
rect 522500 363769 522528 600100
rect 523040 554940 523092 554946
rect 523040 554882 523092 554888
rect 523052 554849 523080 554882
rect 523038 554840 523094 554849
rect 523038 554775 523094 554784
rect 523132 553512 523184 553518
rect 523132 553454 523184 553460
rect 522580 545148 522632 545154
rect 522580 545090 522632 545096
rect 522486 363760 522542 363769
rect 522486 363695 522542 363704
rect 522592 180674 522620 545090
rect 523040 527264 523092 527270
rect 523038 527232 523040 527241
rect 523092 527232 523094 527241
rect 523038 527167 523094 527176
rect 522580 180668 522632 180674
rect 522580 180610 522632 180616
rect 523144 180538 523172 553454
rect 523500 548616 523552 548622
rect 523500 548558 523552 548564
rect 523408 543788 523460 543794
rect 523408 543730 523460 543736
rect 523316 527944 523368 527950
rect 523316 527886 523368 527892
rect 523224 521688 523276 521694
rect 523224 521630 523276 521636
rect 523132 180532 523184 180538
rect 523132 180474 523184 180480
rect 521844 180464 521896 180470
rect 521844 180406 521896 180412
rect 523236 180334 523264 521630
rect 523328 455326 523356 527886
rect 523316 455320 523368 455326
rect 523316 455262 523368 455268
rect 523420 346390 523448 543730
rect 523512 431730 523540 548558
rect 523682 525736 523738 525745
rect 523682 525671 523738 525680
rect 523590 522472 523646 522481
rect 523590 522407 523646 522416
rect 523604 436665 523632 522407
rect 523696 463593 523724 525671
rect 523774 523696 523830 523705
rect 523774 523631 523830 523640
rect 523788 468081 523816 523631
rect 523774 468072 523830 468081
rect 523774 468007 523830 468016
rect 523682 463584 523738 463593
rect 523682 463519 523738 463528
rect 523590 436656 523646 436665
rect 523590 436591 523646 436600
rect 523500 431724 523552 431730
rect 523500 431666 523552 431672
rect 523880 379137 523908 600100
rect 523958 467936 524014 467945
rect 523958 467871 524014 467880
rect 523866 379128 523922 379137
rect 523866 379063 523922 379072
rect 523408 346384 523460 346390
rect 523408 346326 523460 346332
rect 523224 180328 523276 180334
rect 523224 180270 523276 180276
rect 521752 178764 521804 178770
rect 521752 178706 521804 178712
rect 520280 177676 520332 177682
rect 520280 177618 520332 177624
rect 518992 177540 519044 177546
rect 518992 177482 519044 177488
rect 518900 177200 518952 177206
rect 518900 177142 518952 177148
rect 517704 175160 517756 175166
rect 517704 175102 517756 175108
rect 523972 175098 524000 467871
rect 524064 190454 524092 600102
rect 524696 557660 524748 557666
rect 524696 557602 524748 557608
rect 524420 549364 524472 549370
rect 524420 549306 524472 549312
rect 524064 190426 524368 190454
rect 523960 175092 524012 175098
rect 523960 175034 524012 175040
rect 512644 174956 512696 174962
rect 512644 174898 512696 174904
rect 524340 167006 524368 190426
rect 524432 180062 524460 549306
rect 524512 541136 524564 541142
rect 524512 541078 524564 541084
rect 524524 180266 524552 541078
rect 524604 536240 524656 536246
rect 524604 536182 524656 536188
rect 524616 423638 524644 536182
rect 524708 449682 524736 557602
rect 525154 529408 525210 529417
rect 525154 529343 525210 529352
rect 524972 528216 525024 528222
rect 524972 528158 525024 528164
rect 524786 522336 524842 522345
rect 524786 522271 524842 522280
rect 524696 449676 524748 449682
rect 524696 449618 524748 449624
rect 524800 436393 524828 522271
rect 524880 521008 524932 521014
rect 524880 520950 524932 520956
rect 524892 438802 524920 520950
rect 524984 463622 525012 528158
rect 525064 525292 525116 525298
rect 525064 525234 525116 525240
rect 524972 463616 525024 463622
rect 524972 463558 525024 463564
rect 525076 462126 525104 525234
rect 525168 486985 525196 529343
rect 525154 486976 525210 486985
rect 525154 486911 525210 486920
rect 525064 462120 525116 462126
rect 525064 462062 525116 462068
rect 524880 438796 524932 438802
rect 524880 438738 524932 438744
rect 524786 436384 524842 436393
rect 524786 436319 524842 436328
rect 524604 423632 524656 423638
rect 524604 423574 524656 423580
rect 525260 361185 525288 600100
rect 525892 600092 525944 600098
rect 525892 600034 525944 600040
rect 525800 531548 525852 531554
rect 525800 531490 525852 531496
rect 525812 531457 525840 531490
rect 525798 531448 525854 531457
rect 525798 531383 525854 531392
rect 525800 524748 525852 524754
rect 525800 524690 525852 524696
rect 525812 523410 525840 524690
rect 525720 523382 525840 523410
rect 525720 523002 525748 523382
rect 525800 523320 525852 523326
rect 525800 523262 525852 523268
rect 525812 523161 525840 523262
rect 525798 523152 525854 523161
rect 525798 523087 525854 523096
rect 525720 522974 525840 523002
rect 525246 361176 525302 361185
rect 525246 361111 525302 361120
rect 525812 180606 525840 522974
rect 525904 389842 525932 600034
rect 525984 560992 526036 560998
rect 525984 560934 526036 560940
rect 525996 430438 526024 560934
rect 526260 550724 526312 550730
rect 526260 550666 526312 550672
rect 526076 548684 526128 548690
rect 526076 548626 526128 548632
rect 526088 434586 526116 548626
rect 526168 543924 526220 543930
rect 526168 543866 526220 543872
rect 526180 438870 526208 543866
rect 526272 451246 526300 550666
rect 526442 530768 526498 530777
rect 526442 530703 526498 530712
rect 526352 525088 526404 525094
rect 526352 525030 526404 525036
rect 526364 458046 526392 525030
rect 526456 467673 526484 530703
rect 526536 522368 526588 522374
rect 526536 522310 526588 522316
rect 526442 467664 526498 467673
rect 526442 467599 526498 467608
rect 526548 462194 526576 522310
rect 526536 462188 526588 462194
rect 526536 462130 526588 462136
rect 526352 458040 526404 458046
rect 526352 457982 526404 457988
rect 526260 451240 526312 451246
rect 526260 451182 526312 451188
rect 526168 438864 526220 438870
rect 526168 438806 526220 438812
rect 526076 434580 526128 434586
rect 526076 434522 526128 434528
rect 525984 430432 526036 430438
rect 525984 430374 526036 430380
rect 525892 389836 525944 389842
rect 525892 389778 525944 389784
rect 526640 355473 526668 600100
rect 527272 598324 527324 598330
rect 527272 598266 527324 598272
rect 527180 534268 527232 534274
rect 527180 534210 527232 534216
rect 526626 355464 526682 355473
rect 526626 355399 526682 355408
rect 525800 180600 525852 180606
rect 525800 180542 525852 180548
rect 527192 180402 527220 534210
rect 527284 382158 527312 598266
rect 527364 547188 527416 547194
rect 527364 547130 527416 547136
rect 527376 427718 527404 547130
rect 527456 541680 527508 541686
rect 527456 541622 527508 541628
rect 527364 427712 527416 427718
rect 527364 427654 527416 427660
rect 527468 426358 527496 541622
rect 527640 536920 527692 536926
rect 527640 536862 527692 536868
rect 527548 529372 527600 529378
rect 527548 529314 527600 529320
rect 527456 426352 527508 426358
rect 527456 426294 527508 426300
rect 527560 424930 527588 529314
rect 527652 449750 527680 536862
rect 527730 528184 527786 528193
rect 527730 528119 527786 528128
rect 527744 463865 527772 528119
rect 527916 526652 527968 526658
rect 527916 526594 527968 526600
rect 527824 525360 527876 525366
rect 527824 525302 527876 525308
rect 527730 463856 527786 463865
rect 527730 463791 527786 463800
rect 527836 463690 527864 525302
rect 527928 467702 527956 526594
rect 527916 467696 527968 467702
rect 527916 467638 527968 467644
rect 527824 463684 527876 463690
rect 527824 463626 527876 463632
rect 527640 449744 527692 449750
rect 527640 449686 527692 449692
rect 527548 424924 527600 424930
rect 527548 424866 527600 424872
rect 527272 382152 527324 382158
rect 527272 382094 527324 382100
rect 528020 376417 528048 600100
rect 528742 599992 528798 600001
rect 528742 599927 528798 599936
rect 529204 599956 529256 599962
rect 528650 598496 528706 598505
rect 528650 598431 528706 598440
rect 528560 523116 528612 523122
rect 528560 523058 528612 523064
rect 528006 376408 528062 376417
rect 528006 376343 528062 376352
rect 527180 180396 527232 180402
rect 527180 180338 527232 180344
rect 524512 180260 524564 180266
rect 524512 180202 524564 180208
rect 524420 180056 524472 180062
rect 524420 179998 524472 180004
rect 528572 176526 528600 523058
rect 528664 376281 528692 598431
rect 528756 390153 528784 599927
rect 529204 599898 529256 599904
rect 528928 545896 528980 545902
rect 528928 545838 528980 545844
rect 528836 545828 528888 545834
rect 528836 545770 528888 545776
rect 528848 427786 528876 545770
rect 528940 430506 528968 545838
rect 529020 528148 529072 528154
rect 529020 528090 529072 528096
rect 529032 459406 529060 528090
rect 529112 525156 529164 525162
rect 529112 525098 529164 525104
rect 529124 462262 529152 525098
rect 529112 462256 529164 462262
rect 529112 462198 529164 462204
rect 529020 459400 529072 459406
rect 529020 459342 529072 459348
rect 528928 430500 528980 430506
rect 528928 430442 528980 430448
rect 528836 427780 528888 427786
rect 528836 427722 528888 427728
rect 528742 390144 528798 390153
rect 528742 390079 528798 390088
rect 528650 376272 528706 376281
rect 528650 376207 528706 376216
rect 529216 206310 529244 599898
rect 529296 525224 529348 525230
rect 529296 525166 529348 525172
rect 529308 462330 529336 525166
rect 529296 462324 529348 462330
rect 529296 462266 529348 462272
rect 529400 374649 529428 600100
rect 530584 599888 530636 599894
rect 530584 599830 530636 599836
rect 529848 598868 529900 598874
rect 529848 598810 529900 598816
rect 529860 597961 529888 598810
rect 529846 597952 529902 597961
rect 529846 597887 529902 597896
rect 529938 560416 529994 560425
rect 529938 560351 529994 560360
rect 529846 531448 529902 531457
rect 529846 531383 529848 531392
rect 529900 531383 529902 531392
rect 529848 531354 529900 531360
rect 529952 429078 529980 560351
rect 530032 552764 530084 552770
rect 530032 552706 530084 552712
rect 530044 434518 530072 552706
rect 530216 544468 530268 544474
rect 530216 544410 530268 544416
rect 530124 540252 530176 540258
rect 530124 540194 530176 540200
rect 530032 434512 530084 434518
rect 530032 434454 530084 434460
rect 529940 429072 529992 429078
rect 529940 429014 529992 429020
rect 530136 428874 530164 540194
rect 530228 434654 530256 544410
rect 530400 536444 530452 536450
rect 530400 536386 530452 536392
rect 530308 521076 530360 521082
rect 530308 521018 530360 521024
rect 530216 434648 530268 434654
rect 530216 434590 530268 434596
rect 530124 428868 530176 428874
rect 530124 428810 530176 428816
rect 530320 426426 530348 521018
rect 530412 456618 530440 536386
rect 530492 523864 530544 523870
rect 530492 523806 530544 523812
rect 530504 459474 530532 523806
rect 530492 459468 530544 459474
rect 530492 459410 530544 459416
rect 530400 456612 530452 456618
rect 530400 456554 530452 456560
rect 530308 426420 530360 426426
rect 530308 426362 530360 426368
rect 529940 384396 529992 384402
rect 529940 384338 529992 384344
rect 529952 382294 529980 384338
rect 529940 382288 529992 382294
rect 529940 382230 529992 382236
rect 529386 374640 529442 374649
rect 529386 374575 529442 374584
rect 529938 356008 529994 356017
rect 529938 355943 529994 355952
rect 529952 355570 529980 355943
rect 529940 355564 529992 355570
rect 529940 355506 529992 355512
rect 530596 244934 530624 599830
rect 530676 530868 530728 530874
rect 530676 530810 530728 530816
rect 530688 467770 530716 530810
rect 530676 467764 530728 467770
rect 530676 467706 530728 467712
rect 530780 376718 530808 600100
rect 531412 599820 531464 599826
rect 531412 599762 531464 599768
rect 531320 598800 531372 598806
rect 531320 598742 531372 598748
rect 531228 598188 531280 598194
rect 531228 598130 531280 598136
rect 531240 521665 531268 598130
rect 531332 597825 531360 598742
rect 531318 597816 531374 597825
rect 531318 597751 531374 597760
rect 531320 546644 531372 546650
rect 531320 546586 531372 546592
rect 531226 521656 531282 521665
rect 531226 521591 531282 521600
rect 531228 382288 531280 382294
rect 531228 382230 531280 382236
rect 530768 376712 530820 376718
rect 530768 376654 530820 376660
rect 531240 353258 531268 382230
rect 531228 353252 531280 353258
rect 531228 353194 531280 353200
rect 530584 244928 530636 244934
rect 530584 244870 530636 244876
rect 529204 206304 529256 206310
rect 529204 206246 529256 206252
rect 528560 176520 528612 176526
rect 528560 176462 528612 176468
rect 529216 169017 529244 206246
rect 530596 181801 530624 244870
rect 530582 181792 530638 181801
rect 530582 181727 530638 181736
rect 531332 176594 531360 546586
rect 531424 347857 531452 599762
rect 531502 598360 531558 598369
rect 531502 598295 531558 598304
rect 531516 377369 531544 598295
rect 531688 530800 531740 530806
rect 531688 530742 531740 530748
rect 531596 529508 531648 529514
rect 531596 529450 531648 529456
rect 531608 455394 531636 529450
rect 531700 459542 531728 530742
rect 531870 528320 531926 528329
rect 531870 528255 531926 528264
rect 531778 527912 531834 527921
rect 531778 527847 531834 527856
rect 531792 464681 531820 527847
rect 531884 464953 531912 528255
rect 531962 527096 532018 527105
rect 531962 527031 532018 527040
rect 531976 469033 532004 527031
rect 532054 524104 532110 524113
rect 532054 524039 532110 524048
rect 532068 486713 532096 524039
rect 532054 486704 532110 486713
rect 532054 486639 532110 486648
rect 531962 469024 532018 469033
rect 531962 468959 532018 468968
rect 531870 464944 531926 464953
rect 531870 464879 531926 464888
rect 531778 464672 531834 464681
rect 531778 464607 531834 464616
rect 531688 459536 531740 459542
rect 531688 459478 531740 459484
rect 531596 455388 531648 455394
rect 531596 455330 531648 455336
rect 531502 377360 531558 377369
rect 531502 377295 531558 377304
rect 532160 355337 532188 600100
rect 532882 599856 532938 599865
rect 532882 599791 532938 599800
rect 532792 599752 532844 599758
rect 532792 599694 532844 599700
rect 532698 598768 532754 598777
rect 532698 598703 532754 598712
rect 532712 376009 532740 598703
rect 532804 382294 532832 599694
rect 532896 404977 532924 599791
rect 532976 598936 533028 598942
rect 532976 598878 533028 598884
rect 532988 598369 533016 598878
rect 532974 598360 533030 598369
rect 532974 598295 533030 598304
rect 533540 598097 533568 600100
rect 534078 598632 534134 598641
rect 534078 598567 534134 598576
rect 533526 598088 533582 598097
rect 533526 598023 533582 598032
rect 532976 543040 533028 543046
rect 532976 542982 533028 542988
rect 532988 430370 533016 542982
rect 533066 533896 533122 533905
rect 533066 533831 533122 533840
rect 533080 460873 533108 533831
rect 533434 533216 533490 533225
rect 533434 533151 533490 533160
rect 533252 531004 533304 531010
rect 533252 530946 533304 530952
rect 533160 523728 533212 523734
rect 533160 523670 533212 523676
rect 533066 460864 533122 460873
rect 533066 460799 533122 460808
rect 533172 456686 533200 523670
rect 533264 466274 533292 530946
rect 533344 530936 533396 530942
rect 533344 530878 533396 530884
rect 533252 466268 533304 466274
rect 533252 466210 533304 466216
rect 533356 466206 533384 530878
rect 533448 468761 533476 533151
rect 533526 530632 533582 530641
rect 533526 530567 533582 530576
rect 533434 468752 533490 468761
rect 533434 468687 533490 468696
rect 533540 467129 533568 530567
rect 533526 467120 533582 467129
rect 533526 467055 533582 467064
rect 533344 466200 533396 466206
rect 533344 466142 533396 466148
rect 533160 456680 533212 456686
rect 533160 456622 533212 456628
rect 532976 430364 533028 430370
rect 532976 430306 533028 430312
rect 533342 427136 533398 427145
rect 533342 427071 533398 427080
rect 533356 407833 533384 427071
rect 533342 407824 533398 407833
rect 533342 407759 533398 407768
rect 532882 404968 532938 404977
rect 532882 404903 532938 404912
rect 532792 382288 532844 382294
rect 532792 382230 532844 382236
rect 534092 376145 534120 598567
rect 534920 598097 534948 600100
rect 535736 599684 535788 599690
rect 535736 599626 535788 599632
rect 535458 598904 535514 598913
rect 535458 598839 535514 598848
rect 534906 598088 534962 598097
rect 534906 598023 534962 598032
rect 534170 597816 534226 597825
rect 534170 597751 534226 597760
rect 534184 378865 534212 597751
rect 534262 559872 534318 559881
rect 534262 559807 534318 559816
rect 534276 480729 534304 559807
rect 535368 535560 535420 535566
rect 535366 535528 535368 535537
rect 535420 535528 535422 535537
rect 535366 535463 535422 535472
rect 534354 533488 534410 533497
rect 534354 533423 534410 533432
rect 534262 480720 534318 480729
rect 534262 480655 534318 480664
rect 534368 459785 534396 533423
rect 534908 531072 534960 531078
rect 534908 531014 534960 531020
rect 534724 530732 534776 530738
rect 534724 530674 534776 530680
rect 534540 530664 534592 530670
rect 534540 530606 534592 530612
rect 534448 526584 534500 526590
rect 534448 526526 534500 526532
rect 534354 459776 534410 459785
rect 534354 459711 534410 459720
rect 534460 458182 534488 526526
rect 534552 466342 534580 530606
rect 534632 530596 534684 530602
rect 534632 530538 534684 530544
rect 534644 466410 534672 530538
rect 534736 467838 534764 530674
rect 534814 527776 534870 527785
rect 534814 527711 534870 527720
rect 534724 467832 534776 467838
rect 534724 467774 534776 467780
rect 534632 466404 534684 466410
rect 534632 466346 534684 466352
rect 534540 466336 534592 466342
rect 534540 466278 534592 466284
rect 534828 465225 534856 527711
rect 534920 469198 534948 531014
rect 534908 469192 534960 469198
rect 534908 469134 534960 469140
rect 534998 468480 535054 468489
rect 534998 468415 535054 468424
rect 534814 465216 534870 465225
rect 534814 465151 534870 465160
rect 534448 458176 534500 458182
rect 534448 458118 534500 458124
rect 535012 444825 535040 468415
rect 534998 444816 535054 444825
rect 534998 444751 535054 444760
rect 534170 378856 534226 378865
rect 534170 378791 534226 378800
rect 534078 376136 534134 376145
rect 534078 376071 534134 376080
rect 532698 376000 532754 376009
rect 532698 375935 532754 375944
rect 535472 373289 535500 598839
rect 535552 598256 535604 598262
rect 535552 598198 535604 598204
rect 535564 382226 535592 598198
rect 535642 597680 535698 597689
rect 535642 597615 535698 597624
rect 535552 382220 535604 382226
rect 535552 382162 535604 382168
rect 535656 381585 535684 597615
rect 535748 458182 535776 599626
rect 536300 598194 536328 600100
rect 536930 598360 536986 598369
rect 536930 598295 536986 598304
rect 536288 598188 536340 598194
rect 536288 598130 536340 598136
rect 536104 597576 536156 597582
rect 536104 597518 536156 597524
rect 535828 536308 535880 536314
rect 535828 536250 535880 536256
rect 535736 458176 535788 458182
rect 535736 458118 535788 458124
rect 535748 457502 535776 458118
rect 535736 457496 535788 457502
rect 535736 457438 535788 457444
rect 535840 424998 535868 536250
rect 535918 534032 535974 534041
rect 535918 533967 535974 533976
rect 535932 459513 535960 533967
rect 536012 529236 536064 529242
rect 536012 529178 536064 529184
rect 535918 459504 535974 459513
rect 535918 459439 535974 459448
rect 536024 456754 536052 529178
rect 536012 456748 536064 456754
rect 536012 456690 536064 456696
rect 535828 424992 535880 424998
rect 535828 424934 535880 424940
rect 535642 381576 535698 381585
rect 535642 381511 535698 381520
rect 535458 373280 535514 373289
rect 535458 373215 535514 373224
rect 532698 356008 532754 356017
rect 532698 355943 532754 355952
rect 534078 356008 534134 356017
rect 534078 355943 534134 355952
rect 532712 355910 532740 355943
rect 532700 355904 532752 355910
rect 532700 355846 532752 355852
rect 534092 355842 534120 355943
rect 534080 355836 534132 355842
rect 534080 355778 534132 355784
rect 536116 355366 536144 597518
rect 536288 541884 536340 541890
rect 536288 541826 536340 541832
rect 536194 533624 536250 533633
rect 536194 533559 536250 533568
rect 536208 460057 536236 533559
rect 536300 470558 536328 541826
rect 536840 538280 536892 538286
rect 536840 538222 536892 538228
rect 536288 470552 536340 470558
rect 536288 470494 536340 470500
rect 536378 460184 536434 460193
rect 536378 460119 536434 460128
rect 536194 460048 536250 460057
rect 536194 459983 536250 459992
rect 536392 427145 536420 460119
rect 536378 427136 536434 427145
rect 536378 427071 536434 427080
rect 536104 355360 536156 355366
rect 532146 355328 532202 355337
rect 536104 355302 536156 355308
rect 532146 355263 532202 355272
rect 531410 347848 531466 347857
rect 531410 347783 531466 347792
rect 531424 345014 531452 347783
rect 531424 344986 532004 345014
rect 531976 299470 532004 344986
rect 531964 299464 532016 299470
rect 531964 299406 532016 299412
rect 536852 180198 536880 538222
rect 536944 378729 536972 598295
rect 537312 596174 537340 600471
rect 537576 600296 537628 600302
rect 537576 600238 537628 600244
rect 537312 596146 537524 596174
rect 537024 557592 537076 557598
rect 537024 557534 537076 557540
rect 537036 449818 537064 557534
rect 537116 549296 537168 549302
rect 537116 549238 537168 549244
rect 537128 449886 537156 549238
rect 537300 536376 537352 536382
rect 537300 536318 537352 536324
rect 537208 520464 537260 520470
rect 537208 520406 537260 520412
rect 537116 449880 537168 449886
rect 537116 449822 537168 449828
rect 537024 449812 537076 449818
rect 537024 449754 537076 449760
rect 537220 425066 537248 520406
rect 537312 458114 537340 536318
rect 537300 458108 537352 458114
rect 537300 458050 537352 458056
rect 537208 425060 537260 425066
rect 537208 425002 537260 425008
rect 537496 386345 537524 596146
rect 537588 389094 537616 600238
rect 537576 389088 537628 389094
rect 537576 389030 537628 389036
rect 537482 386336 537538 386345
rect 537482 386271 537538 386280
rect 536930 378720 536986 378729
rect 536930 378655 536986 378664
rect 537680 376038 537708 600100
rect 538310 598224 538366 598233
rect 538310 598159 538366 598168
rect 537760 563712 537812 563718
rect 537760 563654 537812 563660
rect 537772 389162 537800 563654
rect 538220 532908 538272 532914
rect 538220 532850 538272 532856
rect 537760 389156 537812 389162
rect 537760 389098 537812 389104
rect 537668 376032 537720 376038
rect 537668 375974 537720 375980
rect 536840 180192 536892 180198
rect 536840 180134 536892 180140
rect 538232 178702 538260 532850
rect 538324 388521 538352 598159
rect 539060 597582 539088 600100
rect 539048 597576 539100 597582
rect 539048 597518 539100 597524
rect 538404 546100 538456 546106
rect 538404 546042 538456 546048
rect 538416 445738 538444 546042
rect 538496 545760 538548 545766
rect 538496 545702 538548 545708
rect 538508 448458 538536 545702
rect 538588 531140 538640 531146
rect 538588 531082 538640 531088
rect 538600 460834 538628 531082
rect 538680 522300 538732 522306
rect 538680 522242 538732 522248
rect 538692 478174 538720 522242
rect 538680 478168 538732 478174
rect 538680 478110 538732 478116
rect 538588 460828 538640 460834
rect 538588 460770 538640 460776
rect 538496 448452 538548 448458
rect 538496 448394 538548 448400
rect 538404 445732 538456 445738
rect 538404 445674 538456 445680
rect 538310 388512 538366 388521
rect 538310 388447 538366 388456
rect 539244 387666 539272 600986
rect 539520 473249 539548 601015
rect 539506 473240 539562 473249
rect 539506 473175 539562 473184
rect 539232 387660 539284 387666
rect 539232 387602 539284 387608
rect 539612 353190 539640 640455
rect 539966 637800 540022 637809
rect 539966 637735 540022 637744
rect 539690 634672 539746 634681
rect 539690 634607 539746 634616
rect 539600 353184 539652 353190
rect 539600 353126 539652 353132
rect 539704 351121 539732 634607
rect 539782 625016 539838 625025
rect 539782 624951 539838 624960
rect 539690 351112 539746 351121
rect 539690 351047 539746 351056
rect 539796 350334 539824 624951
rect 539876 543856 539928 543862
rect 539876 543798 539928 543804
rect 539784 350328 539836 350334
rect 539784 350270 539836 350276
rect 539888 179382 539916 543798
rect 539980 376106 540008 637735
rect 540256 637537 540284 655415
rect 540242 637528 540298 637537
rect 540242 637463 540298 637472
rect 540242 632224 540298 632233
rect 540242 632159 540298 632168
rect 540150 628144 540206 628153
rect 540150 628079 540206 628088
rect 540058 622432 540114 622441
rect 540058 622367 540114 622376
rect 539968 376100 540020 376106
rect 539968 376042 540020 376048
rect 540072 362409 540100 622367
rect 540164 371929 540192 628079
rect 540256 385665 540284 632159
rect 540348 604518 540376 656882
rect 540428 655648 540480 655654
rect 540428 655590 540480 655596
rect 540440 617574 540468 655590
rect 540428 617568 540480 617574
rect 540428 617510 540480 617516
rect 540336 604512 540388 604518
rect 540336 604454 540388 604460
rect 540440 600302 540468 617510
rect 540992 601050 541020 657358
rect 541070 657319 541126 657328
rect 540980 601044 541032 601050
rect 540980 600986 541032 600992
rect 541084 600545 541112 657319
rect 543740 655580 543792 655586
rect 543740 655522 543792 655528
rect 543554 651264 543610 651273
rect 543554 651199 543610 651208
rect 543568 650078 543596 651199
rect 543556 650072 543608 650078
rect 543556 650014 543608 650020
rect 541162 645824 541218 645833
rect 541162 645759 541218 645768
rect 541070 600536 541126 600545
rect 541070 600471 541126 600480
rect 540428 600296 540480 600302
rect 540428 600238 540480 600244
rect 540336 546576 540388 546582
rect 540336 546518 540388 546524
rect 540348 448526 540376 546518
rect 541072 530052 541124 530058
rect 541072 529994 541124 530000
rect 540980 529984 541032 529990
rect 540980 529926 541032 529932
rect 540426 476232 540482 476241
rect 540426 476167 540482 476176
rect 540440 468489 540468 476167
rect 540426 468480 540482 468489
rect 540426 468415 540482 468424
rect 540336 448520 540388 448526
rect 540336 448462 540388 448468
rect 540242 385656 540298 385665
rect 540242 385591 540298 385600
rect 540150 371920 540206 371929
rect 540150 371855 540206 371864
rect 540058 362400 540114 362409
rect 540058 362335 540114 362344
rect 539876 179376 539928 179382
rect 539876 179318 539928 179324
rect 538220 178696 538272 178702
rect 538220 178638 538272 178644
rect 540992 177274 541020 529926
rect 541084 178838 541112 529994
rect 541176 351422 541204 645759
rect 541254 644464 541310 644473
rect 541254 644399 541310 644408
rect 541268 378894 541296 644399
rect 541346 641744 541402 641753
rect 541346 641679 541402 641688
rect 541256 378888 541308 378894
rect 541256 378830 541308 378836
rect 541360 378826 541388 641679
rect 542358 639024 542414 639033
rect 542358 638959 542414 638968
rect 541440 604512 541492 604518
rect 541440 604454 541492 604460
rect 541452 485110 541480 604454
rect 541532 546032 541584 546038
rect 541532 545974 541584 545980
rect 541440 485104 541492 485110
rect 541440 485046 541492 485052
rect 541544 436082 541572 545974
rect 541624 523796 541676 523802
rect 541624 523738 541676 523744
rect 541636 453830 541664 523738
rect 541624 453824 541676 453830
rect 541624 453766 541676 453772
rect 541532 436076 541584 436082
rect 541532 436018 541584 436024
rect 541348 378820 541400 378826
rect 541348 378762 541400 378768
rect 542372 371385 542400 638959
rect 542726 637528 542782 637537
rect 542726 637463 542782 637472
rect 542450 636304 542506 636313
rect 542450 636239 542506 636248
rect 542464 382265 542492 636239
rect 542542 633584 542598 633593
rect 542542 633519 542598 633528
rect 542556 383081 542584 633519
rect 542634 630864 542690 630873
rect 542634 630799 542690 630808
rect 542648 385801 542676 630799
rect 542740 630057 542768 637463
rect 542726 630048 542782 630057
rect 542726 629983 542782 629992
rect 542726 629504 542782 629513
rect 542726 629439 542782 629448
rect 542634 385792 542690 385801
rect 542634 385727 542690 385736
rect 542740 384946 542768 629439
rect 542818 626784 542874 626793
rect 542818 626719 542874 626728
rect 542728 384940 542780 384946
rect 542728 384882 542780 384888
rect 542832 384878 542860 626719
rect 542910 617264 542966 617273
rect 542910 617199 542966 617208
rect 542924 616894 542952 617199
rect 542912 616888 542964 616894
rect 542912 616830 542964 616836
rect 542910 615904 542966 615913
rect 542910 615839 542966 615848
rect 542924 389201 542952 615839
rect 543752 564398 543780 655522
rect 543740 564392 543792 564398
rect 543740 564334 543792 564340
rect 543752 563718 543780 564334
rect 543740 563712 543792 563718
rect 543740 563654 543792 563660
rect 543740 554872 543792 554878
rect 543740 554814 543792 554820
rect 542910 389192 542966 389201
rect 542910 389127 542966 389136
rect 542820 384872 542872 384878
rect 542820 384814 542872 384820
rect 542542 383072 542598 383081
rect 542542 383007 542598 383016
rect 542450 382256 542506 382265
rect 542450 382191 542506 382200
rect 542358 371376 542414 371385
rect 542358 371311 542414 371320
rect 541164 351416 541216 351422
rect 541164 351358 541216 351364
rect 543752 179314 543780 554814
rect 543832 536988 543884 536994
rect 543832 536930 543884 536936
rect 543740 179308 543792 179314
rect 543740 179250 543792 179256
rect 543844 179110 543872 536930
rect 543936 389026 543964 700334
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 547878 699816 547934 699825
rect 547878 699751 547934 699760
rect 546592 657484 546644 657490
rect 546592 657426 546644 657432
rect 544108 657348 544160 657354
rect 544108 657290 544160 657296
rect 544016 657212 544068 657218
rect 544016 657154 544068 657160
rect 543924 389020 543976 389026
rect 543924 388962 543976 388968
rect 544028 386374 544056 657154
rect 544120 387734 544148 657290
rect 544200 657280 544252 657286
rect 544200 657222 544252 657228
rect 544212 390182 544240 657222
rect 545396 657144 545448 657150
rect 545396 657086 545448 657092
rect 545118 647184 545174 647193
rect 545118 647119 545174 647128
rect 544382 630048 544438 630057
rect 544382 629983 544438 629992
rect 544290 597952 544346 597961
rect 544290 597887 544346 597896
rect 544200 390176 544252 390182
rect 544200 390118 544252 390124
rect 544304 388385 544332 597887
rect 544396 460193 544424 629983
rect 545132 601089 545160 647119
rect 545118 601080 545174 601089
rect 545118 601015 545174 601024
rect 544476 533520 544528 533526
rect 544476 533462 544528 533468
rect 544488 460902 544516 533462
rect 545120 527196 545172 527202
rect 545120 527138 545172 527144
rect 544566 526552 544622 526561
rect 544566 526487 544622 526496
rect 544580 476241 544608 526487
rect 544566 476232 544622 476241
rect 544566 476167 544622 476176
rect 544476 460896 544528 460902
rect 544476 460838 544528 460844
rect 544382 460184 544438 460193
rect 544382 460119 544438 460128
rect 544290 388376 544346 388385
rect 544290 388311 544346 388320
rect 544108 387728 544160 387734
rect 544108 387670 544160 387676
rect 544016 386368 544068 386374
rect 544016 386310 544068 386316
rect 545132 179178 545160 527138
rect 545212 523184 545264 523190
rect 545212 523126 545264 523132
rect 545120 179172 545172 179178
rect 545120 179114 545172 179120
rect 543832 179104 543884 179110
rect 543832 179046 543884 179052
rect 545224 179042 545252 523126
rect 545304 520396 545356 520402
rect 545304 520338 545356 520344
rect 545316 179246 545344 520338
rect 545408 386306 545436 657086
rect 545488 657008 545540 657014
rect 545488 656950 545540 656956
rect 546498 656976 546554 656985
rect 545500 390114 545528 656950
rect 546498 656911 546554 656920
rect 545580 616888 545632 616894
rect 545580 616830 545632 616836
rect 545488 390108 545540 390114
rect 545488 390050 545540 390056
rect 545592 388890 545620 616830
rect 545672 544672 545724 544678
rect 545672 544614 545724 544620
rect 545684 431934 545712 544614
rect 545764 535628 545816 535634
rect 545764 535570 545816 535576
rect 545776 442950 545804 535570
rect 545764 442944 545816 442950
rect 545764 442886 545816 442892
rect 545672 431928 545724 431934
rect 545672 431870 545724 431876
rect 545580 388884 545632 388890
rect 545580 388826 545632 388832
rect 545396 386300 545448 386306
rect 545396 386242 545448 386248
rect 546512 386209 546540 656911
rect 546604 387802 546632 657426
rect 546682 657112 546738 657121
rect 546682 657047 546738 657056
rect 546696 388793 546724 657047
rect 546682 388784 546738 388793
rect 546682 388719 546738 388728
rect 546592 387796 546644 387802
rect 546592 387738 546644 387744
rect 546498 386200 546554 386209
rect 546498 386135 546554 386144
rect 545304 179240 545356 179246
rect 545304 179182 545356 179188
rect 545212 179036 545264 179042
rect 545212 178978 545264 178984
rect 541072 178832 541124 178838
rect 541072 178774 541124 178780
rect 540980 177268 541032 177274
rect 540980 177210 541032 177216
rect 531320 176588 531372 176594
rect 531320 176530 531372 176536
rect 529202 169008 529258 169017
rect 529202 168943 529258 168952
rect 524328 167000 524380 167006
rect 524328 166942 524380 166948
rect 524340 166297 524368 166942
rect 524326 166288 524382 166297
rect 524326 166223 524382 166232
rect 500222 159760 500278 159769
rect 500222 159695 500278 159704
rect 547892 158681 547920 699751
rect 580262 697232 580318 697241
rect 580262 697167 580318 697176
rect 548062 657248 548118 657257
rect 548062 657183 548118 657192
rect 547972 657076 548024 657082
rect 547972 657018 548024 657024
rect 547984 387530 548012 657018
rect 548076 388249 548104 657183
rect 549260 650072 549312 650078
rect 549260 650014 549312 650020
rect 548062 388240 548118 388249
rect 548062 388175 548118 388184
rect 547972 387524 548024 387530
rect 547972 387466 548024 387472
rect 549272 376650 549300 650014
rect 580172 617568 580224 617574
rect 580170 617536 580172 617545
rect 580224 617536 580226 617545
rect 580170 617471 580226 617480
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 549260 376644 549312 376650
rect 549260 376586 549312 376592
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580276 351286 580304 697167
rect 580354 644056 580410 644065
rect 580354 643991 580410 644000
rect 580368 384334 580396 643991
rect 580446 431624 580502 431633
rect 580446 431559 580502 431568
rect 580356 384328 580408 384334
rect 580356 384270 580408 384276
rect 580460 354686 580488 431559
rect 580448 354680 580500 354686
rect 580448 354622 580500 354628
rect 580264 351280 580316 351286
rect 580264 351222 580316 351228
rect 580264 349308 580316 349314
rect 580264 349250 580316 349256
rect 580276 325281 580304 349250
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580262 272232 580318 272241
rect 580262 272167 580318 272176
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 244934 580212 245511
rect 580172 244928 580224 244934
rect 580172 244870 580224 244876
rect 580172 206304 580224 206310
rect 580172 206246 580224 206252
rect 580184 205737 580212 206246
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580276 169182 580304 272167
rect 580354 232384 580410 232393
rect 580354 232319 580410 232328
rect 580264 169176 580316 169182
rect 580264 169118 580316 169124
rect 580368 169114 580396 232319
rect 580446 219056 580502 219065
rect 580446 218991 580502 219000
rect 580356 169108 580408 169114
rect 580356 169050 580408 169056
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580460 160721 580488 218991
rect 580538 192536 580594 192545
rect 580538 192471 580594 192480
rect 580552 169046 580580 192471
rect 580540 169040 580592 169046
rect 580540 168982 580592 168988
rect 580446 160712 580502 160721
rect 580446 160647 580502 160656
rect 547878 158672 547934 158681
rect 547878 158607 547934 158616
rect 580170 152688 580226 152697
rect 580170 152623 580226 152632
rect 580184 151842 580212 152623
rect 580172 151836 580224 151842
rect 580172 151778 580224 151784
rect 407764 144356 407816 144362
rect 407764 144298 407816 144304
rect 407210 139224 407266 139233
rect 407210 139159 407266 139168
rect 407776 128081 407804 144298
rect 407762 128072 407818 128081
rect 407762 128007 407818 128016
rect 407210 116920 407266 116929
rect 407210 116855 407266 116864
rect 407118 105768 407174 105777
rect 407118 105703 407174 105712
rect 407224 100609 407252 116855
rect 407210 100600 407266 100609
rect 407210 100535 407266 100544
rect 382476 97889 382504 100028
rect 382462 97880 382518 97889
rect 382462 97815 382518 97824
rect 360660 89004 360712 89010
rect 360660 88946 360712 88952
rect 537484 89004 537536 89010
rect 537484 88946 537536 88952
rect 358084 86964 358136 86970
rect 358084 86906 358136 86912
rect 336278 85640 336334 85649
rect 336278 85575 336334 85584
rect 332690 9072 332746 9081
rect 332690 9007 332746 9016
rect 331864 6860 331916 6866
rect 331864 6802 331916 6808
rect 332704 480 332732 9007
rect 336292 480 336320 85575
rect 364614 85096 364670 85105
rect 364614 85031 364670 85040
rect 357530 84960 357586 84969
rect 357530 84895 357586 84904
rect 343362 84688 343418 84697
rect 343362 84623 343418 84632
rect 339866 3360 339922 3369
rect 339866 3295 339922 3304
rect 339880 480 339908 3295
rect 343376 480 343404 84623
rect 350448 69692 350500 69698
rect 350448 69634 350500 69640
rect 346952 54528 347004 54534
rect 346952 54470 347004 54476
rect 346964 480 346992 54470
rect 350460 480 350488 69634
rect 354036 50380 354088 50386
rect 354036 50322 354088 50328
rect 354048 480 354076 50322
rect 357544 480 357572 84895
rect 361118 84552 361174 84561
rect 361118 84487 361174 84496
rect 361132 480 361160 84487
rect 364628 480 364656 85031
rect 368202 83464 368258 83473
rect 368202 83399 368258 83408
rect 368216 480 368244 83399
rect 435362 83056 435418 83065
rect 435362 82991 435418 83000
rect 432602 81696 432658 81705
rect 432602 81631 432658 81640
rect 428554 80336 428610 80345
rect 428554 80271 428610 80280
rect 421562 77616 421618 77625
rect 421562 77551 421618 77560
rect 417422 76256 417478 76265
rect 417422 76191 417478 76200
rect 414662 74896 414718 74905
rect 414662 74831 414718 74840
rect 411902 57216 411958 57225
rect 411902 57151 411958 57160
rect 389454 40760 389510 40769
rect 389454 40695 389510 40704
rect 385958 16008 386014 16017
rect 385958 15943 386014 15952
rect 378874 14648 378930 14657
rect 378874 14583 378930 14592
rect 375286 11792 375342 11801
rect 375286 11727 375342 11736
rect 371700 10328 371752 10334
rect 371700 10270 371752 10276
rect 371712 480 371740 10270
rect 375300 480 375328 11727
rect 378888 480 378916 14583
rect 382370 13152 382426 13161
rect 382370 13087 382426 13096
rect 382384 480 382412 13087
rect 385972 480 386000 15943
rect 389468 480 389496 40695
rect 400126 39400 400182 39409
rect 400126 39335 400182 39344
rect 396538 21448 396594 21457
rect 396538 21383 396594 21392
rect 393042 18728 393098 18737
rect 393042 18663 393098 18672
rect 393056 480 393084 18663
rect 396552 480 396580 21383
rect 400140 480 400168 39335
rect 407210 38040 407266 38049
rect 407210 37975 407266 37984
rect 403622 17368 403678 17377
rect 403622 17303 403678 17312
rect 403636 480 403664 17303
rect 407224 480 407252 37975
rect 411916 4865 411944 57151
rect 410798 4856 410854 4865
rect 410798 4791 410854 4800
rect 411902 4856 411958 4865
rect 411902 4791 411958 4800
rect 414294 4856 414350 4865
rect 414294 4791 414350 4800
rect 410812 480 410840 4791
rect 414308 480 414336 4791
rect 414676 3097 414704 74831
rect 417436 3505 417464 76191
rect 418802 61296 418858 61305
rect 418802 61231 418858 61240
rect 417882 7712 417938 7721
rect 417882 7647 417938 7656
rect 417422 3496 417478 3505
rect 417422 3431 417478 3440
rect 414662 3088 414718 3097
rect 414662 3023 414718 3032
rect 417896 480 417924 7647
rect 418816 4865 418844 61231
rect 421378 53272 421434 53281
rect 421378 53207 421434 53216
rect 418802 4856 418858 4865
rect 418802 4791 418858 4800
rect 421392 480 421420 53207
rect 421576 3913 421604 77551
rect 422942 68096 422998 68105
rect 422942 68031 422998 68040
rect 422956 7585 422984 68031
rect 425702 62656 425758 62665
rect 425702 62591 425758 62600
rect 422942 7576 422998 7585
rect 422942 7511 422998 7520
rect 424966 4856 425022 4865
rect 424966 4791 425022 4800
rect 421562 3904 421618 3913
rect 421562 3839 421618 3848
rect 424980 480 425008 4791
rect 425716 4185 425744 62591
rect 425702 4176 425758 4185
rect 425702 4111 425758 4120
rect 428462 4176 428518 4185
rect 428462 4111 428518 4120
rect 428476 480 428504 4111
rect 428568 3777 428596 80271
rect 431222 65376 431278 65385
rect 431222 65311 431278 65320
rect 429842 64016 429898 64025
rect 429842 63951 429898 63960
rect 429856 4865 429884 63951
rect 431236 5001 431264 65311
rect 431222 4992 431278 5001
rect 431222 4927 431278 4936
rect 429842 4856 429898 4865
rect 429842 4791 429898 4800
rect 432050 4856 432106 4865
rect 432050 4791 432106 4800
rect 428554 3768 428610 3777
rect 428554 3703 428610 3712
rect 432064 480 432092 4791
rect 432616 3233 432644 81631
rect 435376 3641 435404 82991
rect 450542 73536 450598 73545
rect 450542 73471 450598 73480
rect 447782 72176 447838 72185
rect 447782 72111 447838 72120
rect 443642 70816 443698 70825
rect 443642 70751 443698 70760
rect 436742 66736 436798 66745
rect 436742 66671 436798 66680
rect 435546 4992 435602 5001
rect 435546 4927 435602 4936
rect 435362 3632 435418 3641
rect 435362 3567 435418 3576
rect 432602 3224 432658 3233
rect 432602 3159 432658 3168
rect 435560 480 435588 4927
rect 436756 4185 436784 66671
rect 439502 47832 439558 47841
rect 439502 47767 439558 47776
rect 436742 4176 436798 4185
rect 436742 4111 436798 4120
rect 439134 4176 439190 4185
rect 439134 4111 439190 4120
rect 439148 480 439176 4111
rect 439516 4049 439544 47767
rect 442262 47696 442318 47705
rect 442262 47631 442318 47640
rect 439502 4040 439558 4049
rect 439502 3975 439558 3984
rect 442276 3369 442304 47631
rect 442630 7576 442686 7585
rect 442630 7511 442686 7520
rect 442262 3360 442318 3369
rect 442262 3295 442318 3304
rect 442644 480 442672 7511
rect 443656 4185 443684 70751
rect 446402 47560 446458 47569
rect 446402 47495 446458 47504
rect 443642 4176 443698 4185
rect 443642 4111 443698 4120
rect 446218 4176 446274 4185
rect 446218 4111 446274 4120
rect 442906 4040 442962 4049
rect 442906 3975 442962 3984
rect 442920 2854 442948 3975
rect 442908 2848 442960 2854
rect 442908 2790 442960 2796
rect 446232 480 446260 4111
rect 446416 3466 446444 47495
rect 447796 4185 447824 72111
rect 450556 4865 450584 73471
rect 467470 55856 467526 55865
rect 467470 55791 467526 55800
rect 450542 4856 450598 4865
rect 450542 4791 450598 4800
rect 453302 4856 453358 4865
rect 453302 4791 453358 4800
rect 447782 4176 447838 4185
rect 447782 4111 447838 4120
rect 449806 4176 449862 4185
rect 449806 4111 449862 4120
rect 446404 3460 446456 3466
rect 446404 3402 446456 3408
rect 449820 480 449848 4111
rect 453316 480 453344 4791
rect 463974 3904 464030 3913
rect 463974 3839 464030 3848
rect 460386 3496 460442 3505
rect 460386 3431 460442 3440
rect 456890 3088 456946 3097
rect 456890 3023 456946 3032
rect 456904 480 456932 3023
rect 460400 480 460428 3431
rect 463988 480 464016 3839
rect 467484 480 467512 55791
rect 517150 49056 517206 49065
rect 517150 48991 517206 49000
rect 481730 46336 481786 46345
rect 481730 46271 481786 46280
rect 471058 3768 471114 3777
rect 471058 3703 471114 3712
rect 471072 480 471100 3703
rect 478142 3632 478198 3641
rect 478142 3567 478198 3576
rect 474554 3224 474610 3233
rect 474554 3159 474610 3168
rect 474568 480 474596 3159
rect 478156 480 478184 3567
rect 481744 480 481772 46271
rect 499394 43480 499450 43489
rect 499394 43415 499450 43424
rect 495898 13016 495954 13025
rect 495898 12951 495954 12960
rect 492310 11656 492366 11665
rect 492310 11591 492366 11600
rect 488814 10296 488870 10305
rect 488814 10231 488870 10240
rect 485226 8936 485282 8945
rect 485226 8871 485282 8880
rect 485240 480 485268 8871
rect 488828 480 488856 10231
rect 492324 480 492352 11591
rect 495912 480 495940 12951
rect 499408 480 499436 43415
rect 506478 42120 506534 42129
rect 506478 42055 506534 42064
rect 502982 14512 503038 14521
rect 502982 14447 503038 14456
rect 502996 480 503024 14447
rect 506492 480 506520 42055
rect 512642 40624 512698 40633
rect 512642 40559 512698 40568
rect 510066 15872 510122 15881
rect 510066 15807 510122 15816
rect 510080 480 510108 15807
rect 512656 3505 512684 40559
rect 512642 3496 512698 3505
rect 512642 3431 512698 3440
rect 513562 3496 513618 3505
rect 513562 3431 513618 3440
rect 513576 480 513604 3431
rect 517164 480 517192 48991
rect 537496 46918 537524 88946
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 576122 48920 576178 48929
rect 576122 48855 576178 48864
rect 537484 46912 537536 46918
rect 537484 46854 537536 46860
rect 549074 44840 549130 44849
rect 549074 44775 549130 44784
rect 520738 39264 520794 39273
rect 520738 39199 520794 39208
rect 520752 480 520780 39199
rect 524234 37904 524290 37913
rect 524234 37839 524290 37848
rect 524248 480 524276 37839
rect 527822 36544 527878 36553
rect 527822 36479 527878 36488
rect 527836 480 527864 36479
rect 534906 35184 534962 35193
rect 534906 35119 534962 35128
rect 531318 17232 531374 17241
rect 531318 17167 531374 17176
rect 531332 480 531360 17167
rect 534920 480 534948 35119
rect 538402 33824 538458 33833
rect 538402 33759 538458 33768
rect 538416 480 538444 33759
rect 541990 30968 542046 30977
rect 541990 30903 542046 30912
rect 542004 480 542032 30903
rect 545486 29608 545542 29617
rect 545486 29543 545542 29552
rect 545500 480 545528 29543
rect 549088 480 549116 44775
rect 552662 28248 552718 28257
rect 552662 28183 552718 28192
rect 552676 480 552704 28183
rect 559746 26888 559802 26897
rect 559746 26823 559802 26832
rect 555422 18592 555478 18601
rect 555422 18527 555478 18536
rect 555436 16574 555464 18527
rect 555436 16546 556108 16574
rect 556080 3482 556108 16546
rect 556080 3454 556200 3482
rect 556172 480 556200 3454
rect 559760 480 559788 26823
rect 562322 25528 562378 25537
rect 562322 25463 562378 25472
rect 562336 3505 562364 25463
rect 566830 24168 566886 24177
rect 566830 24103 566886 24112
rect 562322 3496 562378 3505
rect 562322 3431 562378 3440
rect 563242 3496 563298 3505
rect 563242 3431 563298 3440
rect 563256 480 563284 3431
rect 566844 480 566872 24103
rect 570326 22672 570382 22681
rect 570326 22607 570382 22616
rect 570340 480 570368 22607
rect 573914 21312 573970 21321
rect 573914 21247 573970 21256
rect 573928 480 573956 21247
rect 576136 4049 576164 48855
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 576122 4040 576178 4049
rect 576122 3975 576178 3984
rect 577410 4040 577466 4049
rect 577410 3975 577466 3984
rect 577424 480 577452 3975
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 581000 2848 581052 2854
rect 581000 2790 581052 2796
rect 581012 480 581040 2790
rect 582208 480 582236 3295
rect 583404 480 583432 3402
rect 50130 326 50476 354
rect 50130 -960 50242 326
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3422 579944 3478 580000
rect 3422 527856 3478 527912
rect 3422 475632 3478 475688
rect 3422 423544 3478 423600
rect 4066 398112 4122 398168
rect 3422 371320 3478 371376
rect 4066 358672 4122 358728
rect 3422 319232 3478 319288
rect 24306 700304 24362 700360
rect 31022 700304 31078 700360
rect 25686 645088 25742 645144
rect 25502 542816 25558 542872
rect 25502 432248 25558 432304
rect 25870 644136 25926 644192
rect 25686 481208 25742 481264
rect 26054 643184 26110 643240
rect 25870 475768 25926 475824
rect 26054 471416 26110 471472
rect 27434 655016 27490 655072
rect 26790 654200 26846 654256
rect 27250 549616 27306 549672
rect 26974 538464 27030 538520
rect 27066 534112 27122 534168
rect 26974 420824 27030 420880
rect 27066 400696 27122 400752
rect 26790 393624 26846 393680
rect 27250 410488 27306 410544
rect 30194 654472 30250 654528
rect 28262 652840 28318 652896
rect 27434 395800 27490 395856
rect 30010 641280 30066 641336
rect 28538 638560 28594 638616
rect 28446 553016 28502 553072
rect 28354 544040 28410 544096
rect 28722 633936 28778 633992
rect 28538 467608 28594 467664
rect 28446 409944 28502 410000
rect 28354 408856 28410 408912
rect 28262 394168 28318 394224
rect 28814 633800 28870 633856
rect 28722 461080 28778 461136
rect 28814 460536 28870 460592
rect 30102 542272 30158 542328
rect 30010 468152 30066 468208
rect 30286 654336 30342 654392
rect 30286 391448 30342 391504
rect 30194 390904 30250 390960
rect 43074 700304 43130 700360
rect 33046 654608 33102 654664
rect 31666 651616 31722 651672
rect 31298 642368 31354 642424
rect 31206 532888 31262 532944
rect 31114 525136 31170 525192
rect 31114 503648 31170 503704
rect 31390 514800 31446 514856
rect 31298 480664 31354 480720
rect 31206 420280 31262 420336
rect 31390 354456 31446 354512
rect 31022 354320 31078 354376
rect 30102 350376 30158 350432
rect 32862 641960 32918 642016
rect 32678 539824 32734 539880
rect 32586 535608 32642 535664
rect 32494 526904 32550 526960
rect 32402 523368 32458 523424
rect 32402 498616 32458 498672
rect 32494 427352 32550 427408
rect 32678 423000 32734 423056
rect 32586 421912 32642 421968
rect 31666 393080 31722 393136
rect 32954 638016 33010 638072
rect 32862 469240 32918 469296
rect 32954 464888 33010 464944
rect 41326 653656 41382 653712
rect 33782 652976 33838 653032
rect 39670 651072 39726 651128
rect 35714 640464 35770 640520
rect 34334 640056 34390 640112
rect 34242 553696 34298 553752
rect 33874 546760 33930 546816
rect 34150 542408 34206 542464
rect 34058 533704 34114 533760
rect 33966 530712 34022 530768
rect 33874 504600 33930 504656
rect 33966 401240 34022 401296
rect 35622 549480 35678 549536
rect 35530 545944 35586 546000
rect 35254 538600 35310 538656
rect 35162 526496 35218 526552
rect 34334 467064 34390 467120
rect 35346 536968 35402 537024
rect 35254 426808 35310 426864
rect 35162 421368 35218 421424
rect 35438 524592 35494 524648
rect 35346 412120 35402 412176
rect 34242 408312 34298 408368
rect 35438 400152 35494 400208
rect 35530 399608 35586 399664
rect 34150 399064 34206 399120
rect 34058 398520 34114 398576
rect 37186 639240 37242 639296
rect 35806 638152 35862 638208
rect 35714 480120 35770 480176
rect 35622 397976 35678 398032
rect 36634 557776 36690 557832
rect 36542 533024 36598 533080
rect 37002 550976 37058 551032
rect 36910 545264 36966 545320
rect 36818 543904 36874 543960
rect 36726 539688 36782 539744
rect 36634 429528 36690 429584
rect 36542 413208 36598 413264
rect 36726 403960 36782 404016
rect 36818 403416 36874 403472
rect 37002 405048 37058 405104
rect 36910 402872 36966 402928
rect 35806 395256 35862 395312
rect 33782 392536 33838 392592
rect 33046 391992 33102 392048
rect 38474 635024 38530 635080
rect 38106 552336 38162 552392
rect 37922 531936 37978 531992
rect 38014 523640 38070 523696
rect 37922 504056 37978 504112
rect 37922 503648 37978 503704
rect 37922 491816 37978 491872
rect 38382 547848 38438 547904
rect 38198 541184 38254 541240
rect 38106 506232 38162 506288
rect 38014 488824 38070 488880
rect 37186 462712 37242 462768
rect 38290 534928 38346 534984
rect 38198 404504 38254 404560
rect 38474 477400 38530 477456
rect 38382 406136 38438 406192
rect 38290 396888 38346 396944
rect 8114 312432 8170 312488
rect 3422 267144 3478 267200
rect 3422 214920 3478 214976
rect 35162 214104 35218 214160
rect 5262 213016 5318 213072
rect 3422 162832 3478 162888
rect 570 46144 626 46200
rect 4066 17176 4122 17232
rect 2870 8880 2926 8936
rect 1674 5208 1730 5264
rect 31022 211928 31078 211984
rect 6458 210840 6514 210896
rect 21822 118088 21878 118144
rect 7562 115912 7618 115968
rect 13542 112648 13598 112704
rect 9954 104080 10010 104136
rect 7562 71576 7618 71632
rect 8758 20168 8814 20224
rect 7654 3440 7710 3496
rect 11702 100000 11758 100056
rect 12346 6160 12402 6216
rect 11702 3440 11758 3496
rect 18234 109792 18290 109848
rect 14738 98776 14794 98832
rect 17038 3440 17094 3496
rect 18602 106936 18658 106992
rect 18602 3440 18658 3496
rect 19430 2760 19486 2816
rect 30102 117408 30158 117464
rect 26514 117272 26570 117328
rect 24214 94424 24270 94480
rect 23018 93336 23074 93392
rect 28906 88984 28962 89040
rect 27710 16088 27766 16144
rect 33598 117680 33654 117736
rect 32402 109656 32458 109712
rect 31022 17176 31078 17232
rect 31298 6296 31354 6352
rect 34794 97144 34850 97200
rect 39486 558184 39542 558240
rect 39210 552608 39266 552664
rect 39394 527312 39450 527368
rect 39302 521192 39358 521248
rect 39210 507864 39266 507920
rect 39578 535472 39634 535528
rect 39486 431704 39542 431760
rect 39394 402328 39450 402384
rect 39302 397432 39358 397488
rect 39762 650936 39818 650992
rect 39670 502288 39726 502344
rect 39854 650664 39910 650720
rect 39762 494672 39818 494728
rect 40774 650392 40830 650448
rect 40682 536832 40738 536888
rect 40498 532752 40554 532808
rect 39854 491136 39910 491192
rect 39578 396344 39634 396400
rect 40590 530032 40646 530088
rect 40498 419192 40554 419248
rect 40590 405592 40646 405648
rect 41234 648896 41290 648952
rect 40774 506504 40830 506560
rect 40682 401784 40738 401840
rect 41234 473048 41290 473104
rect 42154 650528 42210 650584
rect 42062 557912 42118 557968
rect 41878 530576 41934 530632
rect 41970 520648 42026 520704
rect 41878 508952 41934 509008
rect 41326 461624 41382 461680
rect 42706 650256 42762 650312
rect 42522 642096 42578 642152
rect 42154 498072 42210 498128
rect 42062 434968 42118 435024
rect 41970 419736 42026 419792
rect 42522 479032 42578 479088
rect 42706 469784 42762 469840
rect 43994 647536 44050 647592
rect 43902 582120 43958 582176
rect 43442 558048 43498 558104
rect 43166 547984 43222 548040
rect 43258 527584 43314 527640
rect 43258 498752 43314 498808
rect 43258 496712 43314 496768
rect 43166 496032 43222 496088
rect 43074 353232 43130 353288
rect 43902 552472 43958 552528
rect 43810 521872 43866 521928
rect 43442 493312 43498 493368
rect 45006 638968 45062 639024
rect 44914 578856 44970 578912
rect 44822 576680 44878 576736
rect 44822 555736 44878 555792
rect 44914 555464 44970 555520
rect 44638 549752 44694 549808
rect 44178 527448 44234 527504
rect 44178 525136 44234 525192
rect 44086 521736 44142 521792
rect 44730 538192 44786 538248
rect 44638 510040 44694 510096
rect 44914 533568 44970 533624
rect 44822 528672 44878 528728
rect 44730 500792 44786 500848
rect 44822 475496 44878 475552
rect 45098 591912 45154 591968
rect 45190 589736 45246 589792
rect 45098 560088 45154 560144
rect 45374 590824 45430 590880
rect 45374 558592 45430 558648
rect 45190 557368 45246 557424
rect 45006 493992 45062 494048
rect 44914 472640 44970 472696
rect 43994 471960 44050 472016
rect 53562 649576 53618 649632
rect 51446 649304 51502 649360
rect 46846 644000 46902 644056
rect 46754 594088 46810 594144
rect 46662 579944 46718 580000
rect 46570 577768 46626 577824
rect 46570 556960 46626 557016
rect 46754 559816 46810 559872
rect 46662 555192 46718 555248
rect 46570 551248 46626 551304
rect 46386 545400 46442 545456
rect 46294 534248 46350 534304
rect 46110 522552 46166 522608
rect 46018 519424 46074 519480
rect 46202 520784 46258 520840
rect 46110 508408 46166 508464
rect 46202 498888 46258 498944
rect 46478 520376 46534 520432
rect 46570 516568 46626 516624
rect 46478 496168 46534 496224
rect 46386 418648 46442 418704
rect 46294 418104 46350 418160
rect 46018 363568 46074 363624
rect 49606 643728 49662 643784
rect 48042 643456 48098 643512
rect 47950 581032 48006 581088
rect 47858 575592 47914 575648
rect 47950 556688 48006 556744
rect 47858 556008 47914 556064
rect 47766 548120 47822 548176
rect 47674 545536 47730 545592
rect 47582 522008 47638 522064
rect 47490 521056 47546 521112
rect 47398 519152 47454 519208
rect 47398 508544 47454 508600
rect 47398 506504 47454 506560
rect 46846 394712 46902 394768
rect 47490 499704 47546 499760
rect 47582 496304 47638 496360
rect 47674 425720 47730 425776
rect 47858 521872 47914 521928
rect 47858 505824 47914 505880
rect 47766 424632 47822 424688
rect 48226 642640 48282 642696
rect 48134 640872 48190 640928
rect 48042 458904 48098 458960
rect 49514 595176 49570 595232
rect 49422 587560 49478 587616
rect 49330 586336 49386 586392
rect 49238 585384 49294 585440
rect 49238 557232 49294 557288
rect 49330 557096 49386 557152
rect 49514 560496 49570 560552
rect 49422 555600 49478 555656
rect 49422 552064 49478 552120
rect 49330 544584 49386 544640
rect 49238 541456 49294 541512
rect 49146 538736 49202 538792
rect 49054 537104 49110 537160
rect 48962 535880 49018 535936
rect 48870 521736 48926 521792
rect 48226 457272 48282 457328
rect 48134 456728 48190 456784
rect 48870 506776 48926 506832
rect 49054 438232 49110 438288
rect 49146 437144 49202 437200
rect 48962 436600 49018 436656
rect 50618 641824 50674 641880
rect 50066 639920 50122 639976
rect 50526 550024 50582 550080
rect 50434 546896 50490 546952
rect 50342 545128 50398 545184
rect 50250 539960 50306 540016
rect 50158 523096 50214 523152
rect 50066 463256 50122 463312
rect 49606 459448 49662 459504
rect 49422 436056 49478 436112
rect 49330 433336 49386 433392
rect 49238 432792 49294 432848
rect 50250 435512 50306 435568
rect 50342 430616 50398 430672
rect 50158 426264 50214 426320
rect 50434 424088 50490 424144
rect 50710 637744 50766 637800
rect 50618 482976 50674 483032
rect 50618 482840 50674 482896
rect 50526 422456 50582 422512
rect 50894 637472 50950 637528
rect 50710 464344 50766 464400
rect 52274 649168 52330 649224
rect 51814 648080 51870 648136
rect 51630 533296 51686 533352
rect 50986 527176 51042 527232
rect 50986 520240 51042 520296
rect 51538 526632 51594 526688
rect 51538 520240 51594 520296
rect 51446 465432 51502 465488
rect 50894 462168 50950 462224
rect 51722 528944 51778 529000
rect 51630 434424 51686 434480
rect 51538 433880 51594 433936
rect 52182 647672 52238 647728
rect 52090 647400 52146 647456
rect 51906 642912 51962 642968
rect 51814 482296 51870 482352
rect 51722 417560 51778 417616
rect 51998 641416 52054 641472
rect 51906 476312 51962 476368
rect 51906 475496 51962 475552
rect 52090 476856 52146 476912
rect 52182 474680 52238 474736
rect 53010 646720 53066 646776
rect 52918 639512 52974 639568
rect 52366 520240 52422 520296
rect 52366 519288 52422 519344
rect 52366 476176 52422 476232
rect 52274 474136 52330 474192
rect 52182 472640 52238 472696
rect 51998 472504 52054 472560
rect 52182 407768 52238 407824
rect 51906 407224 51962 407280
rect 53378 640328 53434 640384
rect 53102 503648 53158 503704
rect 53010 470328 53066 470384
rect 52918 463800 52974 463856
rect 53194 425176 53250 425232
rect 53470 574504 53526 574560
rect 53470 556824 53526 556880
rect 54850 649032 54906 649088
rect 54114 647944 54170 648000
rect 53838 558048 53894 558104
rect 53930 557912 53986 557968
rect 53838 556144 53894 556200
rect 53838 554920 53894 554976
rect 53746 529760 53802 529816
rect 53838 523096 53894 523152
rect 53562 478488 53618 478544
rect 53378 475224 53434 475280
rect 54114 470872 54170 470928
rect 54758 641688 54814 641744
rect 54666 635432 54722 635488
rect 54574 634616 54630 634672
rect 54574 599528 54630 599584
rect 54666 597352 54722 597408
rect 54666 588648 54722 588704
rect 54574 584296 54630 584352
rect 54482 572328 54538 572384
rect 54482 558728 54538 558784
rect 54574 558456 54630 558512
rect 54666 556552 54722 556608
rect 54666 544176 54722 544232
rect 54390 538328 54446 538384
rect 54298 459992 54354 460048
rect 54390 412664 54446 412720
rect 54574 513304 54630 513360
rect 54758 481752 54814 481808
rect 56230 648760 56286 648816
rect 55586 640736 55642 640792
rect 54942 640600 54998 640656
rect 54850 477944 54906 478000
rect 55126 583208 55182 583264
rect 55034 573416 55090 573472
rect 55126 559272 55182 559328
rect 55034 555328 55090 555384
rect 55126 527176 55182 527232
rect 55034 520104 55090 520160
rect 56046 635568 56102 635624
rect 56138 612584 56194 612640
rect 56046 596264 56102 596320
rect 55954 570152 56010 570208
rect 55770 566752 55826 566808
rect 56046 558184 56102 558240
rect 56046 557912 56102 557968
rect 55770 552880 55826 552936
rect 56046 552744 56102 552800
rect 56046 546624 56102 546680
rect 55678 542680 55734 542736
rect 55586 466520 55642 466576
rect 54942 465976 54998 466032
rect 54666 411576 54722 411632
rect 55954 542544 56010 542600
rect 55770 541320 55826 541376
rect 55678 431160 55734 431216
rect 55862 499840 55918 499896
rect 55770 411032 55826 411088
rect 55954 409400 56010 409456
rect 56138 545808 56194 545864
rect 56046 406680 56102 406736
rect 56414 647808 56470 647864
rect 56322 641008 56378 641064
rect 56230 479576 56286 479632
rect 56230 478896 56286 478952
rect 56506 640484 56562 640520
rect 56506 640464 56508 640484
rect 56508 640464 56560 640484
rect 56560 640464 56562 640484
rect 57702 635704 57758 635760
rect 57610 624552 57666 624608
rect 56966 622376 57022 622432
rect 56506 567976 56562 568032
rect 57242 621288 57298 621344
rect 57058 604968 57114 605024
rect 56506 554784 56562 554840
rect 56506 552064 56562 552120
rect 56506 545128 56562 545184
rect 57150 562400 57206 562456
rect 57334 611496 57390 611552
rect 57426 609320 57482 609376
rect 57242 549888 57298 549944
rect 57150 542952 57206 543008
rect 57058 536152 57114 536208
rect 56966 532344 57022 532400
rect 56506 513984 56562 514040
rect 57150 532208 57206 532264
rect 57058 526360 57114 526416
rect 57058 512760 57114 512816
rect 56966 511672 57022 511728
rect 57518 593000 57574 593056
rect 57886 642776 57942 642832
rect 57886 641824 57942 641880
rect 58530 637336 58586 637392
rect 58346 634752 58402 634808
rect 57794 631080 57850 631136
rect 57886 625640 57942 625696
rect 57794 623464 57850 623520
rect 57702 600616 57758 600672
rect 57702 563488 57758 563544
rect 57610 560224 57666 560280
rect 57426 547032 57482 547088
rect 57518 532072 57574 532128
rect 57334 517112 57390 517168
rect 57426 515480 57482 515536
rect 57242 513304 57298 513360
rect 57794 550568 57850 550624
rect 57702 544448 57758 544504
rect 58254 615848 58310 615904
rect 58070 603880 58126 603936
rect 58438 614760 58494 614816
rect 58346 598440 58402 598496
rect 58346 564576 58402 564632
rect 58346 553288 58402 553344
rect 58254 547304 58310 547360
rect 58070 540368 58126 540424
rect 57886 539416 57942 539472
rect 57794 531528 57850 531584
rect 57702 523096 57758 523152
rect 57610 516024 57666 516080
rect 57518 512216 57574 512272
rect 57150 511128 57206 511184
rect 57518 510584 57574 510640
rect 57058 496032 57114 496088
rect 57426 503648 57482 503704
rect 57334 500656 57390 500712
rect 57150 493312 57206 493368
rect 57150 491136 57206 491192
rect 57058 489912 57114 489968
rect 56414 473592 56470 473648
rect 56322 468696 56378 468752
rect 57150 428440 57206 428496
rect 57610 505824 57666 505880
rect 57886 531392 57942 531448
rect 57794 514936 57850 514992
rect 66534 646856 66590 646912
rect 62670 645224 62726 645280
rect 59266 642368 59322 642424
rect 59082 642232 59138 642288
rect 59174 641824 59230 641880
rect 59266 641688 59322 641744
rect 59174 640464 59230 640520
rect 59082 633256 59138 633312
rect 59266 640328 59322 640384
rect 66074 639784 66130 639840
rect 66166 638968 66222 639024
rect 63958 636248 64014 636304
rect 66074 636248 66130 636304
rect 65246 635160 65302 635216
rect 71686 646176 71742 646232
rect 67822 646040 67878 646096
rect 70398 636928 70454 636984
rect 69110 636248 69166 636304
rect 89166 700304 89222 700360
rect 135902 700304 135958 700360
rect 87602 657464 87658 657520
rect 115846 646720 115902 646776
rect 115478 646584 115534 646640
rect 112902 646448 112958 646504
rect 73066 646312 73122 646368
rect 91098 645088 91154 645144
rect 92294 645088 92350 645144
rect 84566 644952 84622 645008
rect 80702 644816 80758 644872
rect 76838 644680 76894 644736
rect 75550 644544 75606 644600
rect 74262 637064 74318 637120
rect 73158 636248 73214 636304
rect 79414 638696 79470 638752
rect 78126 638288 78182 638344
rect 82818 638288 82874 638344
rect 83278 638288 83334 638344
rect 81438 638152 81494 638208
rect 81990 637608 82046 637664
rect 88982 640056 89038 640112
rect 88246 639784 88302 639840
rect 89718 639784 89774 639840
rect 87142 639104 87198 639160
rect 86866 638560 86922 638616
rect 85854 638424 85910 638480
rect 109038 639920 109094 639976
rect 110326 639920 110382 639976
rect 107566 639784 107622 639840
rect 106186 639104 106242 639160
rect 106462 639104 106518 639160
rect 105174 638968 105230 639024
rect 102598 638832 102654 638888
rect 102138 638288 102194 638344
rect 98734 635976 98790 636032
rect 95146 635196 95148 635216
rect 95148 635196 95200 635216
rect 95200 635196 95202 635216
rect 95146 635160 95202 635196
rect 92478 635024 92534 635080
rect 93766 635024 93822 635080
rect 94870 634888 94926 634944
rect 98090 634888 98146 634944
rect 99378 635024 99434 635080
rect 100022 634888 100078 634944
rect 104254 635024 104310 635080
rect 104806 634888 104862 634944
rect 108302 637064 108358 637120
rect 107750 636248 107806 636304
rect 109130 635976 109186 636032
rect 109038 635160 109094 635216
rect 111614 638560 111670 638616
rect 110418 637608 110474 637664
rect 114190 645904 114246 645960
rect 116122 646584 116178 646640
rect 116122 645904 116178 645960
rect 131118 645224 131174 645280
rect 132222 645224 132278 645280
rect 126886 644136 126942 644192
rect 124126 644000 124182 644056
rect 125782 644000 125838 644056
rect 123206 643864 123262 643920
rect 118698 638696 118754 638752
rect 119342 638152 119398 638208
rect 117226 636928 117282 636984
rect 116766 636792 116822 636848
rect 118054 636792 118110 636848
rect 117962 636248 118018 636304
rect 121458 637472 121514 637528
rect 121918 636384 121974 636440
rect 125506 636520 125562 636576
rect 125690 636520 125746 636576
rect 127622 641416 127678 641472
rect 127070 641144 127126 641200
rect 129738 638424 129794 638480
rect 130934 637608 130990 637664
rect 128358 637200 128414 637256
rect 128450 636656 128506 636712
rect 128818 636656 128874 636712
rect 129646 636248 129702 636304
rect 133878 636656 133934 636712
rect 133878 634480 133934 634536
rect 120630 634208 120686 634264
rect 59266 632168 59322 632224
rect 59174 629992 59230 630048
rect 58806 618024 58862 618080
rect 58714 607144 58770 607200
rect 58530 601704 58586 601760
rect 58622 571240 58678 571296
rect 58438 529760 58494 529816
rect 58990 616936 59046 616992
rect 58898 613672 58954 613728
rect 58806 559680 58862 559736
rect 58714 559136 58770 559192
rect 58806 558048 58862 558104
rect 58622 529216 58678 529272
rect 57886 513848 57942 513904
rect 57518 498752 57574 498808
rect 57518 498072 57574 498128
rect 57518 496304 57574 496360
rect 57518 492632 57574 492688
rect 57702 496168 57758 496224
rect 57702 491000 57758 491056
rect 57610 486648 57666 486704
rect 57518 437688 57574 437744
rect 59726 608232 59782 608288
rect 59634 569064 59690 569120
rect 59266 565800 59322 565856
rect 59542 561380 59598 561436
rect 59266 557776 59322 557832
rect 59174 552608 59230 552664
rect 59174 551384 59230 551440
rect 59082 548256 59138 548312
rect 58990 544312 59046 544368
rect 58990 534384 59046 534440
rect 58898 529080 58954 529136
rect 58806 491136 58862 491192
rect 58990 430072 59046 430128
rect 58898 428984 58954 429040
rect 59082 427896 59138 427952
rect 59634 553968 59690 554024
rect 59818 606056 59874 606112
rect 59818 602792 59874 602848
rect 59726 548528 59782 548584
rect 59266 538872 59322 538928
rect 59818 536696 59874 536752
rect 60646 560224 60702 560280
rect 60002 553696 60058 553752
rect 59910 532480 59966 532536
rect 59634 531528 59690 531584
rect 59634 527176 59690 527232
rect 59266 519424 59322 519480
rect 59726 519968 59782 520024
rect 59818 519832 59874 519888
rect 60002 522960 60058 523016
rect 59818 518200 59874 518256
rect 59174 423544 59230 423600
rect 60830 552336 60886 552392
rect 60830 538736 60886 538792
rect 60094 517928 60150 517984
rect 60186 505280 60242 505336
rect 60002 500520 60058 500576
rect 59910 390632 59966 390688
rect 60278 497120 60334 497176
rect 61566 552608 61622 552664
rect 61474 539144 61530 539200
rect 64510 558184 64566 558240
rect 63590 558048 63646 558104
rect 63498 548936 63554 548992
rect 62486 535064 62542 535120
rect 60646 519832 60702 519888
rect 60646 519560 60702 519616
rect 60646 519288 60702 519344
rect 62026 526632 62082 526688
rect 61750 526088 61806 526144
rect 61842 520260 61898 520296
rect 61842 520240 61844 520260
rect 61844 520240 61896 520260
rect 61896 520240 61898 520260
rect 68282 558184 68338 558240
rect 67546 551656 67602 551712
rect 66534 547576 66590 547632
rect 67546 546896 67602 546952
rect 65522 533160 65578 533216
rect 68558 537784 68614 537840
rect 69570 525544 69626 525600
rect 69018 525000 69074 525056
rect 71594 543360 71650 543416
rect 72606 542000 72662 542056
rect 74630 546216 74686 546272
rect 75826 545536 75882 545592
rect 75642 544992 75698 545048
rect 75826 544584 75882 544640
rect 73618 540640 73674 540696
rect 76654 536288 76710 536344
rect 70582 525272 70638 525328
rect 70398 524864 70454 524920
rect 68282 524184 68338 524240
rect 68926 523368 68982 523424
rect 62118 520104 62174 520160
rect 78678 549072 78734 549128
rect 79322 548392 79378 548448
rect 81438 551384 81494 551440
rect 81714 551112 81770 551168
rect 80702 550160 80758 550216
rect 80058 550024 80114 550080
rect 82726 543632 82782 543688
rect 83738 542272 83794 542328
rect 82818 541456 82874 541512
rect 79690 540912 79746 540968
rect 86774 545536 86830 545592
rect 86866 545400 86922 545456
rect 88798 547712 88854 547768
rect 88982 546760 89038 546816
rect 88246 544176 88302 544232
rect 88430 544176 88486 544232
rect 85762 539280 85818 539336
rect 86866 538600 86922 538656
rect 84750 537240 84806 537296
rect 85486 537104 85542 537160
rect 77666 523912 77722 523968
rect 78586 523232 78642 523288
rect 80794 527992 80850 528048
rect 89718 535880 89774 535936
rect 89810 534520 89866 534576
rect 91098 539960 91154 540016
rect 90822 536424 90878 536480
rect 92846 550024 92902 550080
rect 92478 549752 92534 549808
rect 91834 540096 91890 540152
rect 93858 529488 93914 529544
rect 94870 528808 94926 528864
rect 95882 529624 95938 529680
rect 95514 529488 95570 529544
rect 95146 528944 95202 529000
rect 96526 529352 96582 529408
rect 97814 553152 97870 553208
rect 97906 553016 97962 553072
rect 98918 553016 98974 553072
rect 98642 552200 98698 552256
rect 99930 550296 99986 550352
rect 99378 549616 99434 549672
rect 100758 538464 100814 538520
rect 101954 538464 102010 538520
rect 100942 535200 100998 535256
rect 100758 534384 100814 534440
rect 95514 528808 95570 528864
rect 95054 528672 95110 528728
rect 104806 539416 104862 539472
rect 103978 539008 104034 539064
rect 102966 527720 103022 527776
rect 107014 540776 107070 540832
rect 107566 539824 107622 539880
rect 109038 538056 109094 538112
rect 112074 551928 112130 551984
rect 111798 551248 111854 551304
rect 111062 549208 111118 549264
rect 110418 548256 110474 548312
rect 110050 537920 110106 537976
rect 109222 535880 109278 535936
rect 109038 535608 109094 535664
rect 108026 535336 108082 535392
rect 108302 534792 108358 534848
rect 106002 533840 106058 533896
rect 106186 533296 106242 533352
rect 104990 526224 105046 526280
rect 114466 553288 114522 553344
rect 114098 552336 114154 552392
rect 116122 537104 116178 537160
rect 117226 536968 117282 537024
rect 117226 535744 117282 535800
rect 117134 535608 117190 535664
rect 115110 533976 115166 534032
rect 115846 533024 115902 533080
rect 113086 527040 113142 527096
rect 106186 526904 106242 526960
rect 111798 526496 111854 526552
rect 119158 551792 119214 551848
rect 118698 550976 118754 551032
rect 120078 527992 120134 528048
rect 121182 527992 121238 528048
rect 120170 527856 120226 527912
rect 122194 528400 122250 528456
rect 123206 528264 123262 528320
rect 121458 527584 121514 527640
rect 120906 527176 120962 527232
rect 118146 524864 118202 524920
rect 117962 524728 118018 524784
rect 126242 545400 126298 545456
rect 126886 545264 126942 545320
rect 127254 543496 127310 543552
rect 127622 542816 127678 542872
rect 128358 541320 128414 541376
rect 129278 541456 129334 541512
rect 131118 550568 131174 550624
rect 131302 550432 131358 550488
rect 132314 544856 132370 544912
rect 131118 544040 131174 544096
rect 130290 541592 130346 541648
rect 129738 541184 129794 541240
rect 125230 527584 125286 527640
rect 135166 530304 135222 530360
rect 125506 528128 125562 528184
rect 125414 527448 125470 527504
rect 124126 527312 124182 527368
rect 124586 527312 124642 527368
rect 135994 636928 136050 636984
rect 136178 636384 136234 636440
rect 137282 638696 137338 638752
rect 137282 638016 137338 638072
rect 137374 636656 137430 636712
rect 137374 626184 137430 626240
rect 137282 620880 137338 620936
rect 137466 618568 137522 618624
rect 137282 611360 137338 611416
rect 137190 575456 137246 575512
rect 137098 572056 137154 572112
rect 137098 555872 137154 555928
rect 137190 554920 137246 554976
rect 136178 546896 136234 546952
rect 136546 546624 136602 546680
rect 135994 538600 136050 538656
rect 136546 538328 136602 538384
rect 137374 606328 137430 606384
rect 137650 607960 137706 608016
rect 137558 604424 137614 604480
rect 137742 592456 137798 592512
rect 137558 531256 137614 531312
rect 137374 530984 137430 531040
rect 137190 530440 137246 530496
rect 163502 700440 163558 700496
rect 154118 700304 154174 700360
rect 202786 700440 202842 700496
rect 176934 700304 176990 700360
rect 218978 700304 219034 700360
rect 235170 700304 235226 700360
rect 173162 698264 173218 698320
rect 176934 698264 176990 698320
rect 160098 687112 160154 687168
rect 163502 687112 163558 687168
rect 164422 688472 164478 688528
rect 173162 688472 173218 688528
rect 158718 685072 158774 685128
rect 160098 685072 160154 685128
rect 162122 677456 162178 677512
rect 163686 677456 163742 677512
rect 153842 674736 153898 674792
rect 158626 674736 158682 674792
rect 158810 667800 158866 667856
rect 162122 667800 162178 667856
rect 157338 665760 157394 665816
rect 158810 665760 158866 665816
rect 151082 662496 151138 662552
rect 153842 662496 153898 662552
rect 137926 588376 137982 588432
rect 149702 649440 149758 649496
rect 151174 657600 151230 657656
rect 157338 657600 157394 657656
rect 323582 700304 323638 700360
rect 178038 655016 178094 655072
rect 177854 654880 177910 654936
rect 177670 654744 177726 654800
rect 151174 649440 151230 649496
rect 153842 639784 153898 639840
rect 154486 639920 154542 639976
rect 176566 647300 176568 647320
rect 176568 647300 176620 647320
rect 176620 647300 176622 647320
rect 176566 647264 176622 647300
rect 176566 645924 176622 645960
rect 176566 645904 176568 645924
rect 176568 645904 176620 645924
rect 176620 645904 176622 645924
rect 177578 640328 177634 640384
rect 175094 637200 175150 637256
rect 173898 635568 173954 635624
rect 166354 626456 166410 626512
rect 166262 623192 166318 623248
rect 164882 607688 164938 607744
rect 163594 603608 163650 603664
rect 162398 595176 162454 595232
rect 162122 594632 162178 594688
rect 159362 581576 159418 581632
rect 153842 530576 153898 530632
rect 159546 581168 159602 581224
rect 159454 579672 159510 579728
rect 159454 555192 159510 555248
rect 159730 581032 159786 581088
rect 159638 578448 159694 578504
rect 159730 556688 159786 556744
rect 159638 555464 159694 555520
rect 159546 552472 159602 552528
rect 162214 571784 162270 571840
rect 162122 530576 162178 530632
rect 162490 592048 162546 592104
rect 162398 560496 162454 560552
rect 163502 591368 163558 591424
rect 162306 559816 162362 559872
rect 162766 576816 162822 576872
rect 162674 576544 162730 576600
rect 162582 558592 162638 558648
rect 162766 556960 162822 557016
rect 163502 556416 163558 556472
rect 162674 555736 162730 555792
rect 162490 554784 162546 554840
rect 164974 589600 165030 589656
rect 165158 587968 165214 588024
rect 165066 569880 165122 569936
rect 164974 557368 165030 557424
rect 166170 569336 166226 569392
rect 165250 556552 165306 556608
rect 166170 559544 166226 559600
rect 165526 556144 165582 556200
rect 165434 556008 165490 556064
rect 165066 555600 165122 555656
rect 164882 555192 164938 555248
rect 163594 531120 163650 531176
rect 164146 530984 164202 531040
rect 166170 546488 166226 546544
rect 166170 530168 166226 530224
rect 169022 624824 169078 624880
rect 167642 624008 167698 624064
rect 166446 605240 166502 605296
rect 166630 590552 166686 590608
rect 166446 530848 166502 530904
rect 166446 521464 166502 521520
rect 166262 520648 166318 520704
rect 166906 582120 166962 582176
rect 166906 581168 166962 581224
rect 166814 560224 166870 560280
rect 166630 556552 166686 556608
rect 166814 546760 166870 546816
rect 166906 537512 166962 537568
rect 166998 521056 167054 521112
rect 167090 520784 167146 520840
rect 167826 622376 167882 622432
rect 167734 589736 167790 589792
rect 167734 556960 167790 557016
rect 167642 521600 167698 521656
rect 168286 585248 168342 585304
rect 168102 585112 168158 585168
rect 168286 558456 168342 558512
rect 168102 557232 168158 557288
rect 168010 557096 168066 557152
rect 168378 549480 168434 549536
rect 168378 535472 168434 535528
rect 167826 521328 167882 521384
rect 168378 520512 168434 520568
rect 171782 619928 171838 619984
rect 170494 600344 170550 600400
rect 170402 598712 170458 598768
rect 169390 591912 169446 591968
rect 169114 573416 169170 573472
rect 169574 590824 169630 590880
rect 170310 588104 170366 588160
rect 169482 581032 169538 581088
rect 169390 559816 169446 559872
rect 169206 556824 169262 556880
rect 169942 578448 169998 578504
rect 169666 577768 169722 577824
rect 169666 576816 169722 576872
rect 169574 558184 169630 558240
rect 169482 550568 169538 550624
rect 169850 559680 169906 559736
rect 169758 559428 169814 559464
rect 169758 559408 169760 559428
rect 169760 559408 169812 559428
rect 169812 559408 169814 559428
rect 170310 556280 170366 556336
rect 170034 555328 170090 555384
rect 170034 552472 170090 552528
rect 169942 548256 169998 548312
rect 169758 548120 169814 548176
rect 169758 543904 169814 543960
rect 169758 539688 169814 539744
rect 169666 536560 169722 536616
rect 170586 599528 170642 599584
rect 170770 597896 170826 597952
rect 170678 592184 170734 592240
rect 171046 596808 171102 596864
rect 170862 594088 170918 594144
rect 171138 574504 171194 574560
rect 171046 559952 171102 560008
rect 170954 559680 171010 559736
rect 170678 544584 170734 544640
rect 170494 540504 170550 540560
rect 170402 534656 170458 534712
rect 169758 534248 169814 534304
rect 169022 520784 169078 520840
rect 171874 615032 171930 615088
rect 173254 615848 173310 615904
rect 173162 612584 173218 612640
rect 171966 601976 172022 602032
rect 172058 601160 172114 601216
rect 172426 586336 172482 586392
rect 172150 583208 172206 583264
rect 172978 579672 173034 579728
rect 172150 559272 172206 559328
rect 172886 561584 172942 561640
rect 172426 557096 172482 557152
rect 172334 555464 172390 555520
rect 172242 551248 172298 551304
rect 172426 550704 172482 550760
rect 172426 541728 172482 541784
rect 173070 575048 173126 575104
rect 172978 560496 173034 560552
rect 172978 559272 173034 559328
rect 172978 558592 173034 558648
rect 173070 554920 173126 554976
rect 173438 614216 173494 614272
rect 173346 602792 173402 602848
rect 174726 634752 174782 634808
rect 174634 613400 174690 613456
rect 174542 610952 174598 611008
rect 173898 596808 173954 596864
rect 173714 587560 173770 587616
rect 173530 587288 173586 587344
rect 173714 575592 173770 575648
rect 174450 574232 174506 574288
rect 173806 569880 173862 569936
rect 173530 557368 173586 557424
rect 174266 558864 174322 558920
rect 173714 554512 173770 554568
rect 173806 553832 173862 553888
rect 174450 555328 174506 555384
rect 173714 549616 173770 549672
rect 173806 549344 173862 549400
rect 176658 636792 176714 636848
rect 176658 635704 176714 635760
rect 175186 634616 175242 634672
rect 175186 633528 175242 633584
rect 177762 636928 177818 636984
rect 177762 629992 177818 630048
rect 189170 653520 189226 653576
rect 184018 652296 184074 652352
rect 178682 642504 178738 642560
rect 178038 642096 178094 642152
rect 177946 641688 178002 641744
rect 177946 640348 178002 640384
rect 177946 640328 177948 640348
rect 177948 640328 178000 640348
rect 178000 640328 178002 640348
rect 177854 627816 177910 627872
rect 177670 626728 177726 626784
rect 177578 623464 177634 623520
rect 177026 611360 177082 611416
rect 175922 610136 175978 610192
rect 174726 598440 174782 598496
rect 174818 597080 174874 597136
rect 174726 593816 174782 593872
rect 174910 585656 174966 585712
rect 175186 585248 175242 585304
rect 175094 585112 175150 585168
rect 175830 584840 175886 584896
rect 175186 584296 175242 584352
rect 174910 572328 174966 572384
rect 175002 570152 175058 570208
rect 174910 558456 174966 558512
rect 174818 548392 174874 548448
rect 173806 530848 173862 530904
rect 173346 530440 173402 530496
rect 175554 570968 175610 571024
rect 175462 560224 175518 560280
rect 175186 558320 175242 558376
rect 175094 556688 175150 556744
rect 175186 556180 175188 556200
rect 175188 556180 175240 556200
rect 175240 556180 175242 556200
rect 175186 556144 175242 556180
rect 175186 547848 175242 547904
rect 175186 547168 175242 547224
rect 175186 540504 175242 540560
rect 175370 540504 175426 540560
rect 175738 559000 175794 559056
rect 175830 556824 175886 556880
rect 175830 556416 175886 556472
rect 175830 554784 175886 554840
rect 175830 550840 175886 550896
rect 175554 533432 175610 533488
rect 176014 606056 176070 606112
rect 176290 595448 176346 595504
rect 176198 583072 176254 583128
rect 176106 579808 176162 579864
rect 176014 556008 176070 556064
rect 175922 536152 175978 536208
rect 175922 532888 175978 532944
rect 175922 531256 175978 531312
rect 176566 588648 176622 588704
rect 176566 587968 176622 588024
rect 176382 584296 176438 584352
rect 176474 582528 176530 582584
rect 176382 559272 176438 559328
rect 176290 555736 176346 555792
rect 176566 559408 176622 559464
rect 176474 550976 176530 551032
rect 176566 549752 176622 549808
rect 176198 536016 176254 536072
rect 176106 530848 176162 530904
rect 177302 609728 177358 609784
rect 177210 607144 177266 607200
rect 177118 569880 177174 569936
rect 177394 608504 177450 608560
rect 177486 601704 177542 601760
rect 179142 638424 179198 638480
rect 179050 637608 179106 637664
rect 178958 635568 179014 635624
rect 178774 633664 178830 633720
rect 178682 621560 178738 621616
rect 177854 610680 177910 610736
rect 177670 607008 177726 607064
rect 177762 604424 177818 604480
rect 178038 593000 178094 593056
rect 178038 592048 178094 592104
rect 178590 584024 178646 584080
rect 178498 573280 178554 573336
rect 178406 568520 178462 568576
rect 178130 556960 178186 557016
rect 178038 556552 178094 556608
rect 178590 556960 178646 557016
rect 178498 555600 178554 555656
rect 178038 555192 178094 555248
rect 177946 554648 178002 554704
rect 178038 554104 178094 554160
rect 178682 548800 178738 548856
rect 178038 547984 178094 548040
rect 178038 541048 178094 541104
rect 177946 532616 178002 532672
rect 178038 531120 178094 531176
rect 178222 530032 178278 530088
rect 178130 529896 178186 529952
rect 178038 526360 178094 526416
rect 177946 525680 178002 525736
rect 177946 523368 178002 523424
rect 178038 522552 178094 522608
rect 179326 636404 179382 636440
rect 179326 636384 179328 636404
rect 179328 636384 179380 636404
rect 179380 636384 179382 636404
rect 179234 635432 179290 635488
rect 179142 634752 179198 634808
rect 179142 633528 179198 633584
rect 179050 601704 179106 601760
rect 178958 600616 179014 600672
rect 179142 599528 179198 599584
rect 185306 652024 185362 652080
rect 187882 651344 187938 651400
rect 186318 650392 186374 650448
rect 186594 650120 186650 650176
rect 185674 635568 185730 635624
rect 185398 635432 185454 635488
rect 190458 653384 190514 653440
rect 194322 653248 194378 653304
rect 191746 637064 191802 637120
rect 191746 636792 191802 636848
rect 227718 652296 227774 652352
rect 211066 651888 211122 651944
rect 208490 651752 208546 651808
rect 207202 651480 207258 651536
rect 205914 649712 205970 649768
rect 196898 648624 196954 648680
rect 198738 648644 198794 648680
rect 198738 648624 198740 648644
rect 198740 648624 198792 648644
rect 198792 648624 198794 648644
rect 200762 648624 200818 648680
rect 205638 648624 205694 648680
rect 213826 651616 213882 651672
rect 214102 651616 214158 651672
rect 227810 652160 227866 652216
rect 212446 650664 212502 650720
rect 212354 650392 212410 650448
rect 226338 651072 226394 651128
rect 214562 650936 214618 650992
rect 214930 650664 214986 650720
rect 226522 650800 226578 650856
rect 224222 649712 224278 649768
rect 223946 649440 224002 649496
rect 227718 638832 227774 638888
rect 231766 650528 231822 650584
rect 232042 650528 232098 650584
rect 227902 638288 227958 638344
rect 227902 637472 227958 637528
rect 229466 636792 229522 636848
rect 233146 652024 233202 652080
rect 233422 652024 233478 652080
rect 234618 648080 234674 648136
rect 235538 648080 235594 648136
rect 323582 657600 323638 657656
rect 359370 654608 359426 654664
rect 356794 654472 356850 654528
rect 305274 653656 305330 653712
rect 235998 636928 236054 636984
rect 237286 637336 237342 637392
rect 240046 637064 240102 637120
rect 237378 636520 237434 636576
rect 239678 636520 239734 636576
rect 238390 636384 238446 636440
rect 261666 644000 261722 644056
rect 259642 643864 259698 643920
rect 251086 641280 251142 641336
rect 249706 641008 249762 641064
rect 259366 641008 259422 641064
rect 249706 640328 249762 640384
rect 242806 637336 242862 637392
rect 242438 636928 242494 636984
rect 245014 637064 245070 637120
rect 247130 637064 247186 637120
rect 246946 636540 247002 636576
rect 246946 636520 246948 636540
rect 246948 636520 247000 636540
rect 247000 636520 247002 636540
rect 247130 636520 247186 636576
rect 245566 636384 245622 636440
rect 246118 636384 246174 636440
rect 258722 638424 258778 638480
rect 250902 638288 250958 638344
rect 249706 636248 249762 636304
rect 258078 638288 258134 638344
rect 256606 638152 256662 638208
rect 255594 635704 255650 635760
rect 248372 634752 248428 634808
rect 237378 634616 237434 634672
rect 243220 634208 243276 634264
rect 179970 633392 180026 633448
rect 179234 597352 179290 597408
rect 179970 594904 180026 594960
rect 179050 593000 179106 593056
rect 178866 580760 178922 580816
rect 178958 578312 179014 578368
rect 179234 579128 179290 579184
rect 179142 577496 179198 577552
rect 179050 560088 179106 560144
rect 179326 576680 179382 576736
rect 179878 576680 179934 576736
rect 179234 541728 179290 541784
rect 179694 563556 179750 563612
rect 179602 563080 179658 563136
rect 179418 556280 179474 556336
rect 179418 556008 179474 556064
rect 254582 588648 254638 588704
rect 253018 560360 253074 560416
rect 233422 560224 233478 560280
rect 180614 558864 180670 558920
rect 180706 558728 180762 558784
rect 179970 557232 180026 557288
rect 179878 555192 179934 555248
rect 180062 551384 180118 551440
rect 185490 551384 185546 551440
rect 185490 550976 185546 551032
rect 179326 531256 179382 531312
rect 179142 531120 179198 531176
rect 178958 530984 179014 531040
rect 178866 526496 178922 526552
rect 179050 522824 179106 522880
rect 184202 541592 184258 541648
rect 184202 522416 184258 522472
rect 184846 521736 184902 521792
rect 204810 541592 204866 541648
rect 216908 560088 216964 560144
rect 208858 542816 208914 542872
rect 208398 542680 208454 542736
rect 214930 526904 214986 526960
rect 214562 526088 214618 526144
rect 216678 559136 216734 559192
rect 217966 544040 218022 544096
rect 216678 543768 216734 543824
rect 215942 532616 215998 532672
rect 215298 531392 215354 531448
rect 218058 539552 218114 539608
rect 218978 540232 219034 540288
rect 219990 520648 220046 520704
rect 221002 521056 221058 521112
rect 220726 520376 220782 520432
rect 222014 539552 222070 539608
rect 222106 538192 222162 538248
rect 224130 545944 224186 546000
rect 224038 545264 224094 545320
rect 223026 533296 223082 533352
rect 223486 532752 223542 532808
rect 222106 521228 222108 521248
rect 222108 521228 222160 521248
rect 222160 521228 222162 521248
rect 222106 521192 222162 521228
rect 224130 522960 224186 523016
rect 226246 558456 226302 558512
rect 225510 539552 225566 539608
rect 225050 538736 225106 538792
rect 224314 533160 224370 533216
rect 225326 524864 225382 524920
rect 224958 524592 225014 524648
rect 224314 522144 224370 522200
rect 226338 555736 226394 555792
rect 227258 555056 227314 555112
rect 227718 557368 227774 557424
rect 227350 553288 227406 553344
rect 227258 552472 227314 552528
rect 226982 539008 227038 539064
rect 226982 522960 227038 523016
rect 226338 522008 226394 522064
rect 228270 556416 228326 556472
rect 228270 551248 228326 551304
rect 228086 548664 228142 548720
rect 227718 548392 227774 548448
rect 227718 521872 227774 521928
rect 228362 549888 228418 549944
rect 230202 557368 230258 557424
rect 229282 549752 229338 549808
rect 228362 522552 228418 522608
rect 230202 555192 230258 555248
rect 230202 553696 230258 553752
rect 230386 556588 230388 556608
rect 230388 556588 230440 556608
rect 230440 556588 230442 556608
rect 230386 556552 230442 556588
rect 230386 554412 230388 554432
rect 230388 554412 230440 554432
rect 230440 554412 230442 554432
rect 230386 554376 230442 554412
rect 230386 551248 230442 551304
rect 230202 549752 230258 549808
rect 231214 558048 231270 558104
rect 231766 557640 231822 557696
rect 231122 547168 231178 547224
rect 231766 547304 231822 547360
rect 231306 536560 231362 536616
rect 232318 549752 232374 549808
rect 232318 548256 232374 548312
rect 233698 560088 233754 560144
rect 233146 536560 233202 536616
rect 234342 555736 234398 555792
rect 234618 553288 234674 553344
rect 234342 550568 234398 550624
rect 234158 526632 234214 526688
rect 233882 525952 233938 526008
rect 236366 558592 236422 558648
rect 235354 552472 235410 552528
rect 235170 547304 235226 547360
rect 235998 551520 236054 551576
rect 235354 546760 235410 546816
rect 235998 541592 236054 541648
rect 236458 550976 236514 551032
rect 237378 559272 237434 559328
rect 237194 541592 237250 541648
rect 238390 558320 238446 558376
rect 237470 526904 237526 526960
rect 238206 526904 238262 526960
rect 240138 559408 240194 559464
rect 240046 555464 240102 555520
rect 240138 554784 240194 554840
rect 239402 554648 239458 554704
rect 240046 554648 240102 554704
rect 239218 543224 239274 543280
rect 240046 553560 240102 553616
rect 240046 542544 240102 542600
rect 240414 559136 240470 559192
rect 240414 554512 240470 554568
rect 240230 523232 240286 523288
rect 241426 556008 241482 556064
rect 241426 554784 241482 554840
rect 241334 536560 241390 536616
rect 241242 536152 241298 536208
rect 241334 523776 241390 523832
rect 242438 557096 242494 557152
rect 242254 543088 242310 543144
rect 243450 558728 243506 558784
rect 243450 558184 243506 558240
rect 243266 549888 243322 549944
rect 242806 542816 242862 542872
rect 244462 559816 244518 559872
rect 245474 559952 245530 560008
rect 244370 542816 244426 542872
rect 244278 542408 244334 542464
rect 244278 540232 244334 540288
rect 245290 539960 245346 540016
rect 248602 560088 248658 560144
rect 246394 559680 246450 559736
rect 246394 558864 246450 558920
rect 245658 557504 245714 557560
rect 247130 557232 247186 557288
rect 247130 555192 247186 555248
rect 247038 554920 247094 554976
rect 247038 540368 247094 540424
rect 247498 555192 247554 555248
rect 247314 540232 247370 540288
rect 247038 524456 247094 524512
rect 248510 553288 248566 553344
rect 248326 525000 248382 525056
rect 249522 553832 249578 553888
rect 249338 526360 249394 526416
rect 249706 552744 249762 552800
rect 250534 557232 250590 557288
rect 250350 534792 250406 534848
rect 249706 525816 249762 525872
rect 251546 557504 251602 557560
rect 251362 544720 251418 544776
rect 251086 534112 251142 534168
rect 252558 559000 252614 559056
rect 252466 557912 252522 557968
rect 252466 544040 252522 544096
rect 252374 537512 252430 537568
rect 252466 536832 252522 536888
rect 253202 552880 253258 552936
rect 253570 552880 253626 552936
rect 253386 539008 253442 539064
rect 253202 522688 253258 522744
rect 255042 577768 255098 577824
rect 254950 576408 255006 576464
rect 254766 575592 254822 575648
rect 254582 556008 254638 556064
rect 253938 546352 253994 546408
rect 253662 539144 253718 539200
rect 254582 538600 254638 538656
rect 253662 522008 253718 522064
rect 254766 553696 254822 553752
rect 255226 574504 255282 574560
rect 255134 573144 255190 573200
rect 255042 558048 255098 558104
rect 254950 557368 255006 557424
rect 255226 556416 255282 556472
rect 255134 555056 255190 555112
rect 255962 633392 256018 633448
rect 255962 600208 256018 600264
rect 255962 594088 256018 594144
rect 255870 584296 255926 584352
rect 255870 559272 255926 559328
rect 256054 589736 256110 589792
rect 255962 558864 256018 558920
rect 256422 587560 256478 587616
rect 256330 585384 256386 585440
rect 256238 582120 256294 582176
rect 256146 578856 256202 578912
rect 256054 557096 256110 557152
rect 256514 569200 256570 569256
rect 256422 559136 256478 559192
rect 256330 558320 256386 558376
rect 256514 553288 256570 553344
rect 256238 552472 256294 552528
rect 256146 549752 256202 549808
rect 257986 598848 258042 598904
rect 257710 575456 257766 575512
rect 257526 572872 257582 572928
rect 257618 571784 257674 571840
rect 257526 558320 257582 558376
rect 257802 572736 257858 572792
rect 257710 559680 257766 559736
rect 257618 555464 257674 555520
rect 257894 572600 257950 572656
rect 257802 554376 257858 554432
rect 256698 553424 256754 553480
rect 256698 553288 256754 553344
rect 256698 552880 256754 552936
rect 257986 554512 258042 554568
rect 256698 530440 256754 530496
rect 257894 530440 257950 530496
rect 256698 526632 256754 526688
rect 258170 599528 258226 599584
rect 259366 638288 259422 638344
rect 258906 635568 258962 635624
rect 258722 598440 258778 598496
rect 258906 597352 258962 597408
rect 258170 557504 258226 557560
rect 259090 595176 259146 595232
rect 259366 591912 259422 591968
rect 258814 557232 258870 557288
rect 259090 561720 259146 561776
rect 258998 559816 259054 559872
rect 258906 555192 258962 555248
rect 258722 553832 258778 553888
rect 258630 546896 258686 546952
rect 258078 524864 258134 524920
rect 257526 522824 257582 522880
rect 256698 522688 256754 522744
rect 259090 533704 259146 533760
rect 260194 637200 260250 637256
rect 260286 635432 260342 635488
rect 260194 601704 260250 601760
rect 260654 634616 260710 634672
rect 260286 600616 260342 600672
rect 260286 559000 260342 559056
rect 260194 553288 260250 553344
rect 297270 643728 297326 643784
rect 294050 642912 294106 642968
rect 293958 642388 294014 642424
rect 293958 642368 293960 642388
rect 293960 642368 294012 642388
rect 294012 642368 294014 642388
rect 294786 642232 294842 642288
rect 294602 642096 294658 642152
rect 262678 641144 262734 641200
rect 287702 636792 287758 636848
rect 285034 634752 285090 634808
rect 263690 634480 263746 634536
rect 284206 611496 284262 611552
rect 270774 551656 270830 551712
rect 266726 548936 266782 548992
rect 264242 547576 264298 547632
rect 265714 535064 265770 535120
rect 264242 522824 264298 522880
rect 264610 522008 264666 522064
rect 270222 537784 270278 537840
rect 267738 524184 267794 524240
rect 269670 522824 269726 522880
rect 268750 522144 268806 522200
rect 269026 522144 269082 522200
rect 270222 522824 270278 522880
rect 277858 546216 277914 546272
rect 274822 543360 274878 543416
rect 272706 525544 272762 525600
rect 271602 522824 271658 522880
rect 271970 522824 272026 522880
rect 271970 522144 272026 522200
rect 273810 525272 273866 525328
rect 275834 542000 275890 542056
rect 276846 540640 276902 540696
rect 278870 544992 278926 545048
rect 279882 536288 279938 536344
rect 283930 550160 283986 550216
rect 281906 549072 281962 549128
rect 280710 523912 280766 523968
rect 282918 540912 282974 540968
rect 284942 551112 284998 551168
rect 284206 546488 284262 546544
rect 285954 543632 286010 543688
rect 285034 534928 285090 534984
rect 285678 528536 285734 528592
rect 286966 542272 287022 542328
rect 288346 578176 288402 578232
rect 288346 550160 288402 550216
rect 288990 539280 289046 539336
rect 287978 537240 288034 537296
rect 288346 526904 288402 526960
rect 288346 520648 288402 520704
rect 291106 585112 291162 585168
rect 289174 581168 289230 581224
rect 290922 581032 290978 581088
rect 289266 579944 289322 580000
rect 289726 570152 289782 570208
rect 289450 567976 289506 568032
rect 289266 560224 289322 560280
rect 289634 564440 289690 564496
rect 289542 563080 289598 563136
rect 289450 556144 289506 556200
rect 289174 555736 289230 555792
rect 289542 552744 289598 552800
rect 289726 549072 289782 549128
rect 290002 545536 290058 545592
rect 290830 544176 290886 544232
rect 291014 580896 291070 580952
rect 291014 542136 291070 542192
rect 290922 539280 290978 539336
rect 291750 572328 291806 572384
rect 291750 558456 291806 558512
rect 291934 622376 291990 622432
rect 295982 638696 296038 638752
rect 294786 625640 294842 625696
rect 294602 624824 294658 624880
rect 292210 596536 292266 596592
rect 292026 590824 292082 590880
rect 292118 586608 292174 586664
rect 292026 558728 292082 558784
rect 292394 583208 292450 583264
rect 292210 569200 292266 569256
rect 292302 566888 292358 566944
rect 292210 558728 292266 558784
rect 292118 554648 292174 554704
rect 291934 554240 291990 554296
rect 292026 547712 292082 547768
rect 291106 524048 291162 524104
rect 291842 521056 291898 521112
rect 292486 562264 292542 562320
rect 292394 558592 292450 558648
rect 292302 551656 292358 551712
rect 295246 601024 295302 601080
rect 294602 593000 294658 593056
rect 293774 568520 293830 568576
rect 292486 543632 292542 543688
rect 293038 534520 293094 534576
rect 292210 533568 292266 533624
rect 293866 565800 293922 565856
rect 293774 555736 293830 555792
rect 295154 590552 295210 590608
rect 295062 589192 295118 589248
rect 294970 586472 295026 586528
rect 294878 569880 294934 569936
rect 294602 560088 294658 560144
rect 294970 559816 295026 559872
rect 294878 552880 294934 552936
rect 295062 547712 295118 547768
rect 293866 546488 293922 546544
rect 295062 540096 295118 540152
rect 294050 536424 294106 536480
rect 295154 538600 295210 538656
rect 295246 535064 295302 535120
rect 296166 636656 296222 636712
rect 296074 550024 296130 550080
rect 295982 522280 296038 522336
rect 297914 643456 297970 643512
rect 297730 643320 297786 643376
rect 297546 642640 297602 642696
rect 297270 633256 297326 633312
rect 297362 623464 297418 623520
rect 297362 621288 297418 621344
rect 296626 597488 296682 597544
rect 296534 596128 296590 596184
rect 296534 587152 296590 587208
rect 296534 586336 296590 586392
rect 296534 577360 296590 577416
rect 296534 576680 296590 576736
rect 296534 567432 296590 567488
rect 296534 567024 296590 567080
rect 296534 557776 296590 557832
rect 296534 557232 296590 557288
rect 296534 550160 296590 550216
rect 296718 587152 296774 587208
rect 296718 586472 296774 586528
rect 297638 640872 297694 640928
rect 297546 628904 297602 628960
rect 297822 635432 297878 635488
rect 297730 631080 297786 631136
rect 297638 627816 297694 627872
rect 298098 642504 298154 642560
rect 298006 640192 298062 640248
rect 297914 632168 297970 632224
rect 298006 629992 298062 630048
rect 297822 626728 297878 626784
rect 298006 620200 298062 620256
rect 298006 619112 298062 619168
rect 298006 618024 298062 618080
rect 297454 616936 297510 616992
rect 297546 609320 297602 609376
rect 297454 608232 297510 608288
rect 297638 606056 297694 606112
rect 298006 613672 298062 613728
rect 298006 612584 298062 612640
rect 297914 603880 297970 603936
rect 297730 569064 297786 569120
rect 297914 561312 297970 561368
rect 298006 542408 298062 542464
rect 298006 526224 298062 526280
rect 296626 525408 296682 525464
rect 296902 522280 296958 522336
rect 296166 522144 296222 522200
rect 298006 522008 298062 522064
rect 324594 650256 324650 650312
rect 314290 649304 314346 649360
rect 307850 639240 307906 639296
rect 310426 639512 310482 639568
rect 311714 637744 311770 637800
rect 323306 641960 323362 642016
rect 316866 640736 316922 640792
rect 315578 640600 315634 640656
rect 345202 649576 345258 649632
rect 334898 649168 334954 649224
rect 332322 648896 332378 648952
rect 327170 647944 327226 648000
rect 329746 647536 329802 647592
rect 328458 643184 328514 643240
rect 333610 647808 333666 647864
rect 343914 649032 343970 649088
rect 336186 647672 336242 647728
rect 341338 647400 341394 647456
rect 347778 648760 347834 648816
rect 358082 654336 358138 654392
rect 363234 654200 363290 654256
rect 360658 652976 360714 653032
rect 364522 652840 364578 652896
rect 370962 641008 371018 641064
rect 369674 640328 369730 640384
rect 369674 636248 369730 636304
rect 304262 634480 304318 634536
rect 299662 634344 299718 634400
rect 302698 634344 302754 634400
rect 303986 634208 304042 634264
rect 299662 633936 299718 633992
rect 374458 636248 374514 636304
rect 374458 632576 374514 632632
rect 374734 626184 374790 626240
rect 374550 624960 374606 625016
rect 375470 639784 375526 639840
rect 374826 624552 374882 624608
rect 374458 623600 374514 623656
rect 374642 618432 374698 618488
rect 374550 613944 374606 614000
rect 374458 612040 374514 612096
rect 299846 604424 299902 604480
rect 299754 602928 299810 602984
rect 299386 601840 299442 601896
rect 299202 594768 299258 594824
rect 299110 571104 299166 571160
rect 299018 561720 299074 561776
rect 298742 560496 298798 560552
rect 299018 560224 299074 560280
rect 299110 551112 299166 551168
rect 299294 592048 299350 592104
rect 299202 543768 299258 543824
rect 299202 543632 299258 543688
rect 298742 540640 298798 540696
rect 299754 552472 299810 552528
rect 299386 536696 299442 536752
rect 299938 597488 299994 597544
rect 299846 534520 299902 534576
rect 299386 529760 299442 529816
rect 299294 529352 299350 529408
rect 302238 560496 302294 560552
rect 305550 560224 305606 560280
rect 307206 553152 307262 553208
rect 306194 529624 306250 529680
rect 305182 528944 305238 529000
rect 302238 528808 302294 528864
rect 299938 523368 299994 523424
rect 302238 522280 302294 522336
rect 304078 522280 304134 522336
rect 303066 522144 303122 522200
rect 301134 521600 301190 521656
rect 300030 521464 300086 521520
rect 299018 521328 299074 521384
rect 302054 520784 302110 520840
rect 303618 522144 303674 522200
rect 308218 553016 308274 553072
rect 309230 550296 309286 550352
rect 310242 535200 310298 535256
rect 311254 538464 311310 538520
rect 310610 530712 310666 530768
rect 312174 527720 312230 527776
rect 313922 555872 313978 555928
rect 320362 549208 320418 549264
rect 316314 540776 316370 540832
rect 313370 523096 313426 523152
rect 313278 522960 313334 523016
rect 315302 533840 315358 533896
rect 314014 522280 314070 522336
rect 314290 522008 314346 522064
rect 319350 537920 319406 537976
rect 318338 535880 318394 535936
rect 317326 535336 317382 535392
rect 321374 551928 321430 551984
rect 322754 558728 322810 558784
rect 323398 552336 323454 552392
rect 322386 527040 322442 527096
rect 328458 551792 328514 551848
rect 325422 537104 325478 537160
rect 324410 533976 324466 534032
rect 326434 535744 326490 535800
rect 327354 524728 327410 524784
rect 331494 528400 331550 528456
rect 330390 527992 330446 528048
rect 329378 527856 329434 527912
rect 336922 552608 336978 552664
rect 335542 545400 335598 545456
rect 332322 528264 332378 528320
rect 334530 527584 334586 527640
rect 333426 527312 333482 527368
rect 336554 543496 336610 543552
rect 338578 541456 338634 541512
rect 340602 550432 340658 550488
rect 339498 522416 339554 522472
rect 341614 544856 341670 544912
rect 345662 553968 345718 554024
rect 347686 529216 347742 529272
rect 350722 544448 350778 544504
rect 349710 542952 349766 543008
rect 350538 542816 350594 542872
rect 350538 539416 350594 539472
rect 352746 538872 352802 538928
rect 356794 532480 356850 532536
rect 358818 548528 358874 548584
rect 359830 547032 359886 547088
rect 362866 545808 362922 545864
rect 361854 522552 361910 522608
rect 363878 529080 363934 529136
rect 366914 544312 366970 544368
rect 374826 607280 374882 607336
rect 374734 569880 374790 569936
rect 387154 646856 387210 646912
rect 383106 645224 383162 645280
rect 380070 642776 380126 642832
rect 379058 640464 379114 640520
rect 375654 621560 375710 621616
rect 376206 619112 376262 619168
rect 375746 617480 375802 617536
rect 375654 610952 375710 611008
rect 375562 608504 375618 608560
rect 375470 606872 375526 606928
rect 375562 603608 375618 603664
rect 375378 602792 375434 602848
rect 375838 613400 375894 613456
rect 375930 601976 375986 602032
rect 376022 597080 376078 597136
rect 376114 595448 376170 595504
rect 375654 532344 375710 532400
rect 376298 615848 376354 615904
rect 377218 622412 377220 622432
rect 377220 622412 377272 622432
rect 377272 622412 377274 622432
rect 377218 622376 377274 622412
rect 376850 620744 376906 620800
rect 378598 619928 378654 619984
rect 378322 616664 378378 616720
rect 378046 606056 378102 606112
rect 377034 605240 377090 605296
rect 378046 604460 378048 604480
rect 378048 604460 378100 604480
rect 378100 604460 378102 604480
rect 378046 604424 378102 604460
rect 376758 600344 376814 600400
rect 376850 598712 376906 598768
rect 376758 597896 376814 597952
rect 377954 594632 378010 594688
rect 378046 593816 378102 593872
rect 378046 593000 378102 593056
rect 378046 592184 378102 592240
rect 378046 591368 378102 591424
rect 378046 590552 378102 590608
rect 378046 589736 378102 589792
rect 376942 588920 376998 588976
rect 378046 588104 378102 588160
rect 377770 587288 377826 587344
rect 378046 586472 378102 586528
rect 378046 585656 378102 585712
rect 378046 584840 378102 584896
rect 378046 584024 378102 584080
rect 378046 583208 378102 583264
rect 378046 582412 378102 582448
rect 378046 582392 378048 582412
rect 378048 582392 378100 582412
rect 378100 582392 378102 582412
rect 377862 581576 377918 581632
rect 377126 580760 377182 580816
rect 377586 579944 377642 580000
rect 377034 579128 377090 579184
rect 377862 578332 377918 578368
rect 377862 578312 377864 578332
rect 377864 578312 377916 578332
rect 377916 578312 377918 578332
rect 377126 575864 377182 575920
rect 376942 575048 376998 575104
rect 378046 573416 378102 573472
rect 378046 572600 378102 572656
rect 378046 571784 378102 571840
rect 378046 570288 378102 570344
rect 377034 569336 377090 569392
rect 377770 568520 377826 568576
rect 376666 522688 376722 522744
rect 378414 611768 378470 611824
rect 378506 610136 378562 610192
rect 378874 609320 378930 609376
rect 378690 601160 378746 601216
rect 378782 596264 378838 596320
rect 378506 532208 378562 532264
rect 378414 532072 378470 532128
rect 377954 522824 378010 522880
rect 378782 522144 378838 522200
rect 381082 641824 381138 641880
rect 380990 576680 381046 576736
rect 380990 523640 381046 523696
rect 380898 522960 380954 523016
rect 386510 599528 386566 599584
rect 386510 531936 386566 531992
rect 392214 646312 392270 646368
rect 391202 646176 391258 646232
rect 388166 646040 388222 646096
rect 392582 634480 392638 634536
rect 392582 613264 392638 613320
rect 395250 644680 395306 644736
rect 394238 644544 394294 644600
rect 393962 635160 394018 635216
rect 393962 522416 394018 522472
rect 407394 645088 407450 645144
rect 401322 644952 401378 645008
rect 398286 644816 398342 644872
rect 397550 613264 397606 613320
rect 397550 607144 397606 607200
rect 397458 599664 397514 599720
rect 400954 607144 401010 607200
rect 400954 596808 401010 596864
rect 429842 657736 429898 657792
rect 461582 652160 461638 652216
rect 425610 646720 425666 646776
rect 424598 646584 424654 646640
rect 423586 646448 423642 646504
rect 418526 639104 418582 639160
rect 417514 638968 417570 639024
rect 416502 635024 416558 635080
rect 416042 596808 416098 596864
rect 416042 536696 416098 536752
rect 420458 522416 420514 522472
rect 422574 638560 422630 638616
rect 427634 559544 427690 559600
rect 426622 548800 426678 548856
rect 432694 555600 432750 555656
rect 428646 540504 428702 540560
rect 429658 533432 429714 533488
rect 431682 522280 431738 522336
rect 433706 555328 433762 555384
rect 445850 556960 445906 557016
rect 443826 551384 443882 551440
rect 439778 541728 439834 541784
rect 436374 536696 436430 536752
rect 436374 532480 436430 532536
rect 436742 531256 436798 531312
rect 437754 531120 437810 531176
rect 438766 530984 438822 531040
rect 440882 532480 440938 532536
rect 440790 530848 440846 530904
rect 440882 528400 440938 528456
rect 441710 526496 441766 526552
rect 444838 536016 444894 536072
rect 444286 528400 444342 528456
rect 444286 526496 444342 526552
rect 446862 556824 446918 556880
rect 447874 556688 447930 556744
rect 455970 544584 456026 544640
rect 459006 530576 459062 530632
rect 461030 554104 461086 554160
rect 461766 650800 461822 650856
rect 461674 648080 461730 648136
rect 461582 523640 461638 523696
rect 475382 654880 475438 654936
rect 463146 653520 463202 653576
rect 461766 530712 461822 530768
rect 461674 521464 461730 521520
rect 465722 653384 465778 653440
rect 463146 533432 463202 533488
rect 464066 534656 464122 534712
rect 471334 653248 471390 653304
rect 469862 651888 469918 651944
rect 468482 651752 468538 651808
rect 467378 650664 467434 650720
rect 467194 650392 467250 650448
rect 465722 533568 465778 533624
rect 465906 636928 465962 636984
rect 465906 536016 465962 536072
rect 467286 649440 467342 649496
rect 467286 530576 467342 530632
rect 467194 527856 467250 527912
rect 467378 527720 467434 527776
rect 468574 636520 468630 636576
rect 468482 528128 468538 528184
rect 468574 521600 468630 521656
rect 470046 636384 470102 636440
rect 469862 523504 469918 523560
rect 471334 533840 471390 533896
rect 478234 651344 478290 651400
rect 475566 642232 475622 642288
rect 475382 533024 475438 533080
rect 475750 642096 475806 642152
rect 475566 522416 475622 522472
rect 475750 522280 475806 522336
rect 478234 533976 478290 534032
rect 507766 670656 507822 670712
rect 482466 654744 482522 654800
rect 479614 652024 479670 652080
rect 480994 650120 481050 650176
rect 480902 632576 480958 632632
rect 480902 613264 480958 613320
rect 479614 527040 479670 527096
rect 481546 524320 481602 524376
rect 482466 530848 482522 530904
rect 485042 650528 485098 650584
rect 485042 533160 485098 533216
rect 485042 533060 485044 533080
rect 485044 533060 485096 533080
rect 485096 533060 485098 533080
rect 485042 533024 485098 533060
rect 488170 654472 488226 654528
rect 487986 651616 488042 651672
rect 487802 651480 487858 651536
rect 487066 613264 487122 613320
rect 487066 599528 487122 599584
rect 488078 641144 488134 641200
rect 488078 600072 488134 600128
rect 488170 599800 488226 599856
rect 487986 528264 488042 528320
rect 487802 525680 487858 525736
rect 489274 633664 489330 633720
rect 489826 657872 489882 657928
rect 494702 657872 494758 657928
rect 489826 599936 489882 599992
rect 489550 520512 489606 520568
rect 491114 657736 491170 657792
rect 543462 699760 543518 699816
rect 507766 657328 507822 657384
rect 515586 657600 515642 657656
rect 515586 657056 515642 657112
rect 521106 657464 521162 657520
rect 537666 657192 537722 657248
rect 535458 657056 535514 657112
rect 536286 657056 536342 657112
rect 535458 655560 535514 655616
rect 539046 656920 539102 656976
rect 540242 655424 540298 655480
rect 500406 654472 500462 654528
rect 539598 640464 539654 640520
rect 539414 608640 539470 608696
rect 539414 601704 539470 601760
rect 539506 601024 539562 601080
rect 537298 600480 537354 600536
rect 490746 598168 490802 598224
rect 494886 598440 494942 598496
rect 497646 598304 497702 598360
rect 490562 522144 490618 522200
rect 498106 521600 498162 521656
rect 498106 520512 498162 520568
rect 497370 520104 497426 520160
rect 499026 598712 499082 598768
rect 499026 550160 499082 550216
rect 500406 598576 500462 598632
rect 501418 559680 501474 559736
rect 500038 555736 500094 555792
rect 499762 549888 499818 549944
rect 499670 547304 499726 547360
rect 499578 534148 499580 534168
rect 499580 534148 499632 534168
rect 499632 534148 499634 534168
rect 499578 534112 499634 534148
rect 499578 531428 499580 531448
rect 499580 531428 499632 531448
rect 499632 531428 499634 531448
rect 499578 531392 499634 531428
rect 499578 520104 499634 520160
rect 499578 519560 499634 519616
rect 499854 543224 499910 543280
rect 500038 521872 500094 521928
rect 501142 541592 501198 541648
rect 500130 521056 500186 521112
rect 500958 539416 501014 539472
rect 500958 533704 501014 533760
rect 500958 529216 501014 529272
rect 500958 528572 500960 528592
rect 500960 528572 501012 528592
rect 501012 528572 501014 528592
rect 500958 528536 501014 528572
rect 500314 520512 500370 520568
rect 500314 520104 500370 520160
rect 500406 519968 500462 520024
rect 500222 487192 500278 487248
rect 500222 482840 500278 482896
rect 500222 474544 500278 474600
rect 500130 451288 500186 451344
rect 500130 444508 500186 444544
rect 500130 444488 500132 444508
rect 500132 444488 500184 444508
rect 500184 444488 500186 444508
rect 500130 443400 500186 443456
rect 500130 442312 500186 442368
rect 500222 442040 500278 442096
rect 499578 391856 499634 391912
rect 60922 390632 60978 390688
rect 498290 390632 498346 390688
rect 323582 390360 323638 390416
rect 316590 390224 316646 390280
rect 60922 389000 60978 389056
rect 66902 389000 66958 389056
rect 66902 384920 66958 384976
rect 68926 384920 68982 384976
rect 69202 381928 69258 381984
rect 71778 381928 71834 381984
rect 70122 380432 70178 380488
rect 71778 380160 71834 380216
rect 73618 380296 73674 380352
rect 71870 355544 71926 355600
rect 77574 380160 77630 380216
rect 77574 377032 77630 377088
rect 80610 384920 80666 384976
rect 80702 377032 80758 377088
rect 78862 373496 78918 373552
rect 81438 367648 81494 367704
rect 77114 359624 77170 359680
rect 82358 359080 82414 359136
rect 75366 351736 75422 351792
rect 68374 348200 68430 348256
rect 71686 347792 71742 347848
rect 62026 345072 62082 345128
rect 50342 340040 50398 340096
rect 49330 303184 49386 303240
rect 48042 302912 48098 302968
rect 41878 184728 41934 184784
rect 37186 117816 37242 117872
rect 35990 101360 36046 101416
rect 35162 8880 35218 8936
rect 40682 117544 40738 117600
rect 38382 91840 38438 91896
rect 39578 90344 39634 90400
rect 44270 117952 44326 118008
rect 43074 106800 43130 106856
rect 45466 185816 45522 185872
rect 47950 301008 48006 301064
rect 47858 119992 47914 120048
rect 48134 302368 48190 302424
rect 48226 255040 48282 255096
rect 49606 303048 49662 303104
rect 49514 301144 49570 301200
rect 49422 300872 49478 300928
rect 49330 237360 49386 237416
rect 48226 185000 48282 185056
rect 48226 173168 48282 173224
rect 49422 120400 49478 120456
rect 50526 302776 50582 302832
rect 50434 302232 50490 302288
rect 50434 120536 50490 120592
rect 62026 303184 62082 303240
rect 61290 301144 61346 301200
rect 63498 302368 63554 302424
rect 66166 303048 66222 303104
rect 68926 302912 68982 302968
rect 66074 301008 66130 301064
rect 71594 302812 71596 302832
rect 71596 302812 71648 302832
rect 71648 302812 71650 302832
rect 71594 302776 71650 302812
rect 85854 347656 85910 347712
rect 84106 346296 84162 346352
rect 86222 321544 86278 321600
rect 75826 302912 75882 302968
rect 71226 300872 71282 300928
rect 74262 302232 74318 302288
rect 81070 302232 81126 302288
rect 86222 302912 86278 302968
rect 88154 367648 88210 367704
rect 88154 365744 88210 365800
rect 87602 346160 87658 346216
rect 89350 344936 89406 344992
rect 91098 341536 91154 341592
rect 94502 365744 94558 365800
rect 94502 350512 94558 350568
rect 94594 348880 94650 348936
rect 92846 343576 92902 343632
rect 96342 385736 96398 385792
rect 95882 350512 95938 350568
rect 95882 339360 95938 339416
rect 97262 339360 97318 339416
rect 96526 302232 96582 302288
rect 99838 349696 99894 349752
rect 98090 347520 98146 347576
rect 101586 346024 101642 346080
rect 105082 352688 105138 352744
rect 103334 343440 103390 343496
rect 98642 339496 98698 339552
rect 104806 339768 104862 339824
rect 97722 300872 97778 300928
rect 97262 300056 97318 300112
rect 106830 365200 106886 365256
rect 108578 344800 108634 344856
rect 112074 351600 112130 351656
rect 113822 348744 113878 348800
rect 110326 341400 110382 341456
rect 119066 367648 119122 367704
rect 122562 379208 122618 379264
rect 120814 366288 120870 366344
rect 129554 377576 129610 377632
rect 127806 370776 127862 370832
rect 126058 349832 126114 349888
rect 124310 347384 124366 347440
rect 134798 386008 134854 386064
rect 136546 383016 136602 383072
rect 133050 381792 133106 381848
rect 143538 384512 143594 384568
rect 141790 376488 141846 376544
rect 140042 373768 140098 373824
rect 138294 345752 138350 345808
rect 145286 344528 145342 344584
rect 131302 344256 131358 344312
rect 117318 343304 117374 343360
rect 115570 340720 115626 340776
rect 113822 321408 113878 321464
rect 105910 301008 105966 301064
rect 110326 300056 110382 300112
rect 107244 299648 107300 299704
rect 108900 299512 108956 299568
rect 110418 291760 110474 291816
rect 52918 238040 52974 238096
rect 53102 237360 53158 237416
rect 56230 238312 56286 238368
rect 59266 238176 59322 238232
rect 57794 237904 57850 237960
rect 61198 237360 61254 237416
rect 62854 236952 62910 237008
rect 66166 238448 66222 238504
rect 64510 235728 64566 235784
rect 56506 235320 56562 235376
rect 54574 234504 54630 234560
rect 55126 187312 55182 187368
rect 59266 232600 59322 232656
rect 58622 230424 58678 230480
rect 57518 202136 57574 202192
rect 57426 199280 57482 199336
rect 57334 185272 57390 185328
rect 57150 184864 57206 184920
rect 57242 173168 57298 173224
rect 57150 144744 57206 144800
rect 56506 124616 56562 124672
rect 57702 198056 57758 198112
rect 57610 185408 57666 185464
rect 57518 176432 57574 176488
rect 57426 175208 57482 175264
rect 57886 191120 57942 191176
rect 57794 187176 57850 187232
rect 57886 179424 57942 179480
rect 57794 177928 57850 177984
rect 58990 196560 59046 196616
rect 58898 193976 58954 194032
rect 58806 185680 58862 185736
rect 57886 174936 57942 174992
rect 58622 174936 58678 174992
rect 57886 172352 57942 172408
rect 57702 158752 57758 158808
rect 58898 162696 58954 162752
rect 59082 192616 59138 192672
rect 58990 160112 59046 160168
rect 58806 156576 58862 156632
rect 59174 187720 59230 187776
rect 59082 155896 59138 155952
rect 57610 154400 57666 154456
rect 57794 143384 57850 143440
rect 57794 134136 57850 134192
rect 57334 128424 57390 128480
rect 61382 223896 61438 223952
rect 60278 221720 60334 221776
rect 59910 220632 59966 220688
rect 60002 220088 60058 220144
rect 59910 182008 59966 182064
rect 59266 167048 59322 167104
rect 60094 217232 60150 217288
rect 60002 143384 60058 143440
rect 60186 197920 60242 197976
rect 60094 132504 60150 132560
rect 61474 222808 61530 222864
rect 69478 237224 69534 237280
rect 71134 237088 71190 237144
rect 77436 240080 77492 240136
rect 79414 239944 79470 240000
rect 74446 237768 74502 237824
rect 72790 236816 72846 236872
rect 81438 238040 81494 238096
rect 82726 238040 82782 238096
rect 81070 236680 81126 236736
rect 88706 240080 88762 240136
rect 88706 239536 88762 239592
rect 88246 238312 88302 238368
rect 88982 238176 89038 238232
rect 86866 237904 86922 237960
rect 87694 237904 87750 237960
rect 86038 237632 86094 237688
rect 90684 240080 90740 240136
rect 93306 240080 93362 240136
rect 93490 240080 93546 240136
rect 92340 239808 92396 239864
rect 93306 239808 93362 239864
rect 93490 239536 93546 239592
rect 95974 239536 96030 239592
rect 94318 239400 94374 239456
rect 97630 238584 97686 238640
rect 89350 237496 89406 237552
rect 98642 238448 98698 238504
rect 100666 238448 100722 238504
rect 99194 238312 99250 238368
rect 102598 238176 102654 238232
rect 102138 238040 102194 238096
rect 104254 238040 104310 238096
rect 107566 239264 107622 239320
rect 108394 238448 108450 238504
rect 108118 238312 108174 238368
rect 104806 237904 104862 237960
rect 105910 237904 105966 237960
rect 99378 237768 99434 237824
rect 106186 237632 106242 237688
rect 108854 237768 108910 237824
rect 108302 237496 108358 237552
rect 97906 237360 97962 237416
rect 84106 236544 84162 236600
rect 75826 235592 75882 235648
rect 67546 219272 67602 219328
rect 64142 215328 64198 215384
rect 61474 185408 61530 185464
rect 112442 291760 112498 291816
rect 112442 275304 112498 275360
rect 92386 187040 92442 187096
rect 64142 185272 64198 185328
rect 61382 184864 61438 184920
rect 148782 352960 148838 353016
rect 152278 384648 152334 384704
rect 154026 365336 154082 365392
rect 150530 348608 150586 348664
rect 147034 341808 147090 341864
rect 159270 364112 159326 364168
rect 161018 362480 161074 362536
rect 157522 361392 157578 361448
rect 162766 343168 162822 343224
rect 166262 367920 166318 367976
rect 169758 379344 169814 379400
rect 171506 375128 171562 375184
rect 168010 366560 168066 366616
rect 180246 381928 180302 381984
rect 183742 383288 183798 383344
rect 181994 377984 182050 378040
rect 178498 374992 178554 375048
rect 185490 372000 185546 372056
rect 176750 370912 176806 370968
rect 175002 349968 175058 350024
rect 187238 348472 187294 348528
rect 173254 346976 173310 347032
rect 188986 345480 189042 345536
rect 164514 341672 164570 341728
rect 155774 340584 155830 340640
rect 192482 380840 192538 380896
rect 195978 375808 196034 375864
rect 194230 369280 194286 369336
rect 199474 353096 199530 353152
rect 204718 368192 204774 368248
rect 202970 365608 203026 365664
rect 201222 351192 201278 351248
rect 197726 344392 197782 344448
rect 211710 372272 211766 372328
rect 213458 366696 213514 366752
rect 209962 362888 210018 362944
rect 208214 361528 208270 361584
rect 216954 386144 217010 386200
rect 211802 350648 211858 350704
rect 209042 350512 209098 350568
rect 206466 342080 206522 342136
rect 190734 340448 190790 340504
rect 113914 275304 113970 275360
rect 113914 264968 113970 265024
rect 115202 264968 115258 265024
rect 115202 242800 115258 242856
rect 116582 242800 116638 242856
rect 116582 224984 116638 225040
rect 118054 224984 118110 225040
rect 118054 222264 118110 222320
rect 122102 222128 122158 222184
rect 122102 207984 122158 208040
rect 124126 207984 124182 208040
rect 124126 204040 124182 204096
rect 113822 187312 113878 187368
rect 60278 168680 60334 168736
rect 60186 130872 60242 130928
rect 59174 126520 59230 126576
rect 57242 122712 57298 122768
rect 57242 121488 57298 121544
rect 86314 120536 86370 120592
rect 82818 120400 82874 120456
rect 55126 120264 55182 120320
rect 88062 120264 88118 120320
rect 53102 119856 53158 119912
rect 46846 117000 46902 117056
rect 70398 119992 70454 120048
rect 74078 119856 74134 119912
rect 93306 119856 93362 119912
rect 95054 119720 95110 119776
rect 96802 119584 96858 119640
rect 100298 117136 100354 117192
rect 106186 117156 106242 117192
rect 106186 117136 106188 117156
rect 106188 117136 106240 117156
rect 106240 117136 106242 117156
rect 98550 117000 98606 117056
rect 107566 117000 107622 117056
rect 68834 116864 68890 116920
rect 106922 116456 106978 116512
rect 63590 115232 63646 115288
rect 85670 112512 85726 112568
rect 46662 102720 46718 102776
rect 52918 86944 52974 87000
rect 50986 85856 51042 85912
rect 54666 87760 54722 87816
rect 63866 87624 63922 87680
rect 62026 87488 62082 87544
rect 59266 87352 59322 87408
rect 57610 87216 57666 87272
rect 56230 87080 56286 87136
rect 60738 86944 60794 87000
rect 60738 86128 60794 86184
rect 60646 85720 60702 85776
rect 65614 87896 65670 87952
rect 84842 87624 84898 87680
rect 68650 85992 68706 86048
rect 66994 85584 67050 85640
rect 69800 84768 69856 84824
rect 80748 85040 80804 85096
rect 77620 84904 77676 84960
rect 71364 84632 71420 84688
rect 79184 84496 79240 84552
rect 82312 84224 82368 84280
rect 48134 81640 48190 81696
rect 47674 65320 47730 65376
rect 47582 62600 47638 62656
rect 47490 55800 47546 55856
rect 47950 63960 48006 64016
rect 47858 59880 47914 59936
rect 47766 58520 47822 58576
rect 47674 43560 47730 43616
rect 47766 25472 47822 25528
rect 48042 61240 48098 61296
rect 47950 48864 48006 48920
rect 47858 24112 47914 24168
rect 48226 80280 48282 80336
rect 85026 87352 85082 87408
rect 85210 87080 85266 87136
rect 85210 82048 85266 82104
rect 85026 80688 85082 80744
rect 84842 79328 84898 79384
rect 49330 78920 49386 78976
rect 49238 68040 49294 68096
rect 49054 66680 49110 66736
rect 48226 49272 48282 49328
rect 49146 54440 49202 54496
rect 49054 49000 49110 49056
rect 48134 42200 48190 42256
rect 50250 77288 50306 77344
rect 49606 76200 49662 76256
rect 49514 73480 49570 73536
rect 49422 70760 49478 70816
rect 49330 44784 49386 44840
rect 49238 39208 49294 39264
rect 49422 36488 49478 36544
rect 49514 35128 49570 35184
rect 50158 71848 50214 71904
rect 49606 30912 49662 30968
rect 49146 28192 49202 28248
rect 48042 22616 48098 22672
rect 47582 21256 47638 21312
rect 47490 18536 47546 18592
rect 50342 74568 50398 74624
rect 50434 68992 50490 69048
rect 50526 56616 50582 56672
rect 50434 37848 50490 37904
rect 50342 33768 50398 33824
rect 50434 29688 50490 29744
rect 50250 29552 50306 29608
rect 50158 17176 50214 17232
rect 48962 5072 49018 5128
rect 47858 3440 47914 3496
rect 85578 53216 85634 53272
rect 50618 52536 50674 52592
rect 84474 51448 84530 51504
rect 82082 50224 82138 50280
rect 50986 47776 51042 47832
rect 52366 47640 52422 47696
rect 53746 47504 53802 47560
rect 53746 44920 53802 44976
rect 51354 36624 51410 36680
rect 50618 32544 50674 32600
rect 50526 26832 50582 26888
rect 51722 22888 51778 22944
rect 52550 10376 52606 10432
rect 51722 3440 51778 3496
rect 56506 46280 56562 46336
rect 55862 35264 55918 35320
rect 55034 19896 55090 19952
rect 56046 32680 56102 32736
rect 54942 3984 54998 4040
rect 55862 3984 55918 4040
rect 58438 24248 58494 24304
rect 57794 8880 57850 8936
rect 57242 3168 57298 3224
rect 60646 47912 60702 47968
rect 62762 47912 62818 47968
rect 61934 12960 61990 13016
rect 64786 46960 64842 47016
rect 65614 46960 65670 47016
rect 63314 43424 63370 43480
rect 62854 33904 62910 33960
rect 62762 11600 62818 11656
rect 59174 10240 59230 10296
rect 59634 7792 59690 7848
rect 65522 25608 65578 25664
rect 63222 20032 63278 20088
rect 62026 3440 62082 3496
rect 62854 3440 62910 3496
rect 60830 3304 60886 3360
rect 64326 3576 64382 3632
rect 66074 42064 66130 42120
rect 67914 49136 67970 49192
rect 67454 15816 67510 15872
rect 65614 14456 65670 14512
rect 66718 9152 66774 9208
rect 68834 40568 68890 40624
rect 69110 26968 69166 27024
rect 70306 17448 70362 17504
rect 71502 22752 71558 22808
rect 71042 4800 71098 4856
rect 72606 31048 72662 31104
rect 72422 11736 72478 11792
rect 74446 46960 74502 47016
rect 75182 46960 75238 47016
rect 74998 46144 75054 46200
rect 72974 14592 73030 14648
rect 73802 11872 73858 11928
rect 76194 28328 76250 28384
rect 75182 13096 75238 13152
rect 77114 40704 77170 40760
rect 81254 39344 81310 39400
rect 80702 21392 80758 21448
rect 79322 18672 79378 18728
rect 76562 15952 76618 16008
rect 80886 14728 80942 14784
rect 77390 13232 77446 13288
rect 79690 6432 79746 6488
rect 78586 4936 78642 4992
rect 83278 29824 83334 29880
rect 84014 37984 84070 38040
rect 83462 17312 83518 17368
rect 85578 5208 85634 5264
rect 87970 111152 88026 111208
rect 86866 98912 86922 98968
rect 86406 87760 86462 87816
rect 86222 87216 86278 87272
rect 86406 53080 86462 53136
rect 86222 51720 86278 51776
rect 87786 87896 87842 87952
rect 87602 87488 87658 87544
rect 87786 9016 87842 9072
rect 87602 7520 87658 7576
rect 98642 108432 98698 108488
rect 93950 102856 94006 102912
rect 91558 101496 91614 101552
rect 90362 95784 90418 95840
rect 89166 72392 89222 72448
rect 90454 62736 90510 62792
rect 90454 3576 90510 3632
rect 92754 3576 92810 3632
rect 97446 97280 97502 97336
rect 95146 94560 95202 94616
rect 97262 87488 97318 87544
rect 96250 64096 96306 64152
rect 97262 3576 97318 3632
rect 104530 105576 104586 105632
rect 99838 105440 99894 105496
rect 101034 104216 101090 104272
rect 102782 100136 102838 100192
rect 102230 3576 102286 3632
rect 102782 3440 102838 3496
rect 103334 3440 103390 3496
rect 105542 78920 105598 78976
rect 105542 55800 105598 55856
rect 105726 3712 105782 3768
rect 121458 118088 121514 118144
rect 122286 118088 122342 118144
rect 121274 115640 121330 115696
rect 119526 115504 119582 115560
rect 112810 114144 112866 114200
rect 110510 113736 110566 113792
rect 108118 89120 108174 89176
rect 109314 3848 109370 3904
rect 111614 90480 111670 90536
rect 114006 111016 114062 111072
rect 119526 110608 119582 110664
rect 119894 109928 119950 109984
rect 116398 102992 116454 103048
rect 115202 91704 115258 91760
rect 118790 93064 118846 93120
rect 117594 58656 117650 58712
rect 121090 60016 121146 60072
rect 178682 312432 178738 312488
rect 125690 302232 125746 302288
rect 126886 301552 126942 301608
rect 126334 300736 126390 300792
rect 126886 300736 126942 300792
rect 126242 204312 126298 204368
rect 125506 116320 125562 116376
rect 125230 115776 125286 115832
rect 123574 115368 123630 115424
rect 123482 57296 123538 57352
rect 124678 61376 124734 61432
rect 123574 32408 123630 32464
rect 126426 205400 126482 205456
rect 126334 119856 126390 119912
rect 126610 203224 126666 203280
rect 126426 3848 126482 3904
rect 126242 3712 126298 3768
rect 127714 141752 127770 141808
rect 127622 140120 127678 140176
rect 127438 131960 127494 132016
rect 127346 130328 127402 130384
rect 127254 127064 127310 127120
rect 126978 119720 127034 119776
rect 127346 120808 127402 120864
rect 127898 138488 127954 138544
rect 127806 128696 127862 128752
rect 127714 121080 127770 121136
rect 127622 120012 127678 120048
rect 127622 119992 127624 120012
rect 127624 119992 127676 120012
rect 127676 119992 127678 120012
rect 127438 119448 127494 119504
rect 127530 119312 127586 119368
rect 127622 119040 127678 119096
rect 128082 135224 128138 135280
rect 128266 133592 128322 133648
rect 127898 120944 127954 121000
rect 128082 125432 128138 125488
rect 127806 119584 127862 119640
rect 127990 119584 128046 119640
rect 128266 119176 128322 119232
rect 127254 118904 127310 118960
rect 129094 204040 129150 204096
rect 129094 196016 129150 196072
rect 129094 120672 129150 120728
rect 130290 196016 130346 196072
rect 130290 193160 130346 193216
rect 130382 178200 130438 178256
rect 129830 117136 129886 117192
rect 126978 116592 127034 116648
rect 126610 3576 126666 3632
rect 131210 299648 131266 299704
rect 131486 193160 131542 193216
rect 131486 184864 131542 184920
rect 131210 117000 131266 117056
rect 131210 115640 131266 115696
rect 133878 301008 133934 301064
rect 132590 300872 132646 300928
rect 133142 184864 133198 184920
rect 133142 176704 133198 176760
rect 135258 299512 135314 299568
rect 134522 176704 134578 176760
rect 134522 167048 134578 167104
rect 133878 115504 133934 115560
rect 175922 244568 175978 244624
rect 159362 208664 159418 208720
rect 155222 206488 155278 206544
rect 146942 190168 146998 190224
rect 140042 187992 140098 188048
rect 137282 183640 137338 183696
rect 136546 167048 136602 167104
rect 136638 160112 136694 160168
rect 135258 115368 135314 115424
rect 130382 109792 130438 109848
rect 138662 174936 138718 174992
rect 137650 113872 137706 113928
rect 137282 91840 137338 91896
rect 130566 77832 130622 77888
rect 134154 76472 134210 76528
rect 138662 53216 138718 53272
rect 141422 179288 141478 179344
rect 142802 176024 142858 176080
rect 141422 93336 141478 93392
rect 141238 93200 141294 93256
rect 140042 10376 140098 10432
rect 143446 160112 143502 160168
rect 143446 155896 143502 155952
rect 144734 109792 144790 109848
rect 142802 20168 142858 20224
rect 151082 180376 151138 180432
rect 147678 155896 147734 155952
rect 147678 153312 147734 153368
rect 148322 114008 148378 114064
rect 146942 7792 146998 7848
rect 155222 114144 155278 114200
rect 175922 187176 175978 187232
rect 209042 239400 209098 239456
rect 209318 338544 209374 338600
rect 212262 349016 212318 349072
rect 212078 348336 212134 348392
rect 211894 347928 211950 347984
rect 211802 236544 211858 236600
rect 212262 347792 212318 347848
rect 212170 345208 212226 345264
rect 212078 240080 212134 240136
rect 212446 348200 212502 348256
rect 214562 344936 214618 344992
rect 213182 344664 213238 344720
rect 212354 343984 212410 344040
rect 212262 239944 212318 240000
rect 212446 343032 212502 343088
rect 212446 239264 212502 239320
rect 212354 237904 212410 237960
rect 212170 237768 212226 237824
rect 214746 344120 214802 344176
rect 214378 343576 214434 343632
rect 214286 342624 214342 342680
rect 214470 343440 214526 343496
rect 214654 343304 214710 343360
rect 214562 343168 214618 343224
rect 216678 345072 216734 345128
rect 216678 344800 216734 344856
rect 215114 343576 215170 343632
rect 214930 342352 214986 342408
rect 214286 238448 214342 238504
rect 214838 342216 214894 342272
rect 214654 341264 214710 341320
rect 214654 239536 214710 239592
rect 216678 341556 216734 341592
rect 216678 341536 216680 341556
rect 216680 341536 216732 341556
rect 216732 341536 216734 341556
rect 216770 340720 216826 340776
rect 216678 339768 216734 339824
rect 216862 339496 216918 339552
rect 215114 339088 215170 339144
rect 215114 238584 215170 238640
rect 214930 238312 214986 238368
rect 214746 238176 214802 238232
rect 214562 238040 214618 238096
rect 218794 350920 218850 350976
rect 218702 347112 218758 347168
rect 218058 344256 218114 344312
rect 217966 340992 218022 341048
rect 217782 339904 217838 339960
rect 217598 339768 217654 339824
rect 217966 298016 218022 298072
rect 217782 239808 217838 239864
rect 217598 239672 217654 239728
rect 213182 236952 213238 237008
rect 218978 350784 219034 350840
rect 220082 348064 220138 348120
rect 218978 247968 219034 248024
rect 220726 348880 220782 348936
rect 220726 347656 220782 347712
rect 220450 347248 220506 347304
rect 220726 346296 220782 346352
rect 221002 346296 221058 346352
rect 220266 345888 220322 345944
rect 221002 345888 221058 345944
rect 220726 341400 220782 341456
rect 220726 340584 220782 340640
rect 220358 243480 220414 243536
rect 220266 236816 220322 236872
rect 220082 236680 220138 236736
rect 218794 235728 218850 235784
rect 211894 235592 211950 235648
rect 216126 224984 216182 225040
rect 199382 209752 199438 209808
rect 188342 195608 188398 195664
rect 186962 177112 187018 177168
rect 178682 157528 178738 157584
rect 180246 115096 180302 115152
rect 176658 114416 176714 114472
rect 166078 114280 166134 114336
rect 162490 114144 162546 114200
rect 159362 109928 159418 109984
rect 155406 108296 155462 108352
rect 151818 73752 151874 73808
rect 151082 16088 151138 16144
rect 158902 91840 158958 91896
rect 170402 112784 170458 112840
rect 173162 79464 173218 79520
rect 169574 3576 169630 3632
rect 170402 3576 170458 3632
rect 186962 112648 187018 112704
rect 183742 111288 183798 111344
rect 187330 101632 187386 101688
rect 198002 186904 198058 186960
rect 191746 117136 191802 117192
rect 190826 116728 190882 116784
rect 188342 13232 188398 13288
rect 195242 109928 195298 109984
rect 197910 107072 197966 107128
rect 194414 3576 194470 3632
rect 195242 3576 195298 3632
rect 211802 207440 211858 207496
rect 209042 201048 209098 201104
rect 206282 191256 206338 191312
rect 205086 112648 205142 112704
rect 201498 94696 201554 94752
rect 199382 57296 199438 57352
rect 198002 5072 198058 5128
rect 208582 108568 208638 108624
rect 206282 20032 206338 20088
rect 210422 189080 210478 189136
rect 209042 94560 209098 94616
rect 216126 198056 216182 198112
rect 215942 197784 215998 197840
rect 214562 196696 214618 196752
rect 213182 182552 213238 182608
rect 212446 116320 212502 116376
rect 212170 116184 212226 116240
rect 211802 102992 211858 103048
rect 210422 32680 210478 32736
rect 213182 97144 213238 97200
rect 215666 114960 215722 115016
rect 214562 14728 214618 14784
rect 220082 194520 220138 194576
rect 219254 105712 219310 105768
rect 215942 51448 215998 51504
rect 221554 347792 221610 347848
rect 221462 235320 221518 235376
rect 222106 351736 222162 351792
rect 222014 351328 222070 351384
rect 223486 381656 223542 381712
rect 223394 376216 223450 376272
rect 222198 350104 222254 350160
rect 222106 348744 222162 348800
rect 223302 347520 223358 347576
rect 223210 346160 223266 346216
rect 223118 346024 223174 346080
rect 223026 345888 223082 345944
rect 222842 345072 222898 345128
rect 222014 339668 222016 339688
rect 222016 339668 222068 339688
rect 222068 339668 222070 339688
rect 222014 339632 222070 339668
rect 221922 339496 221978 339552
rect 222106 255312 222162 255368
rect 223302 345752 223358 345808
rect 223302 341808 223358 341864
rect 223394 292440 223450 292496
rect 224774 389816 224830 389872
rect 223946 369416 224002 369472
rect 224222 351600 224278 351656
rect 224222 348608 224278 348664
rect 224222 346568 224278 346624
rect 224222 344528 224278 344584
rect 224222 342488 224278 342544
rect 224222 340176 224278 340232
rect 224222 339632 224278 339688
rect 224406 348200 224462 348256
rect 224682 351464 224738 351520
rect 223486 290264 223542 290320
rect 224314 326304 224370 326360
rect 224222 259392 224278 259448
rect 223026 237224 223082 237280
rect 222842 237088 222898 237144
rect 221554 234504 221610 234560
rect 222842 202000 222898 202056
rect 220358 191120 220414 191176
rect 222750 111424 222806 111480
rect 220082 11872 220138 11928
rect 224222 192344 224278 192400
rect 222842 108432 222898 108488
rect 224406 261024 224462 261080
rect 225694 386960 225750 387016
rect 226246 375944 226302 376000
rect 226154 373224 226210 373280
rect 224866 351872 224922 351928
rect 224774 293528 224830 293584
rect 224682 256672 224738 256728
rect 225050 347384 225106 347440
rect 224958 346976 225014 347032
rect 225786 346976 225842 347032
rect 225878 345344 225934 345400
rect 224958 341672 225014 341728
rect 225970 289720 226026 289776
rect 226154 298968 226210 299024
rect 227626 387912 227682 387968
rect 227534 376352 227590 376408
rect 227442 364248 227498 364304
rect 226338 350396 226394 350432
rect 226338 350376 226340 350396
rect 226340 350376 226392 350396
rect 226392 350376 226394 350396
rect 227350 349560 227406 349616
rect 227166 349424 227222 349480
rect 226982 349288 227038 349344
rect 226430 348472 226486 348528
rect 226338 347928 226394 347984
rect 226522 347792 226578 347848
rect 226338 345480 226394 345536
rect 226246 295704 226302 295760
rect 226062 282240 226118 282296
rect 227074 348608 227130 348664
rect 227074 283872 227130 283928
rect 227534 318688 227590 318744
rect 227350 292032 227406 292088
rect 227166 278976 227222 279032
rect 226982 277344 227038 277400
rect 224866 253952 224922 254008
rect 227166 240216 227222 240272
rect 227166 199280 227222 199336
rect 226982 198872 227038 198928
rect 224314 164056 224370 164112
rect 229006 382880 229062 382936
rect 228914 378800 228970 378856
rect 228822 377304 228878 377360
rect 228730 376080 228786 376136
rect 227718 345072 227774 345128
rect 228730 326440 228786 326496
rect 228822 323584 228878 323640
rect 228914 311072 228970 311128
rect 228546 300736 228602 300792
rect 230386 383696 230442 383752
rect 230202 381112 230258 381168
rect 230110 378936 230166 378992
rect 230018 375400 230074 375456
rect 229190 371048 229246 371104
rect 229926 351092 229928 351112
rect 229928 351092 229980 351112
rect 229980 351092 229982 351112
rect 229926 351056 229982 351092
rect 229006 291352 229062 291408
rect 228362 219272 228418 219328
rect 228362 199960 228418 200016
rect 227626 148960 227682 149016
rect 226982 111152 227038 111208
rect 226338 108432 226394 108488
rect 224222 9152 224278 9208
rect 229926 340448 229982 340504
rect 230018 320864 230074 320920
rect 230110 313112 230166 313168
rect 230202 307672 230258 307728
rect 229834 301416 229890 301472
rect 229742 187040 229798 187096
rect 230294 252456 230350 252512
rect 231766 387776 231822 387832
rect 231674 384376 231730 384432
rect 231582 384240 231638 384296
rect 231490 381520 231546 381576
rect 231398 380976 231454 381032
rect 231306 378664 231362 378720
rect 230938 352416 230994 352472
rect 231122 342760 231178 342816
rect 231122 340992 231178 341048
rect 231122 338816 231178 338872
rect 231214 326304 231270 326360
rect 231306 312160 231362 312216
rect 231398 306584 231454 306640
rect 231122 302776 231178 302832
rect 231490 301144 231546 301200
rect 230386 219544 230442 219600
rect 231582 218456 231638 218512
rect 231582 217640 231638 217696
rect 231674 217368 231730 217424
rect 233146 388048 233202 388104
rect 233054 384104 233110 384160
rect 232778 383152 232834 383208
rect 232686 373088 232742 373144
rect 232594 367784 232650 367840
rect 232502 317328 232558 317384
rect 232594 285912 232650 285968
rect 232962 362752 233018 362808
rect 232870 359352 232926 359408
rect 232778 288088 232834 288144
rect 233054 258712 233110 258768
rect 232962 257624 233018 257680
rect 232870 256536 232926 256592
rect 232686 255448 232742 255504
rect 231766 151000 231822 151056
rect 234342 381384 234398 381440
rect 233606 378528 233662 378584
rect 234158 374856 234214 374912
rect 233882 370640 233938 370696
rect 233790 361256 233846 361312
rect 233698 355816 233754 355872
rect 233698 282648 233754 282704
rect 234066 369144 234122 369200
rect 233882 281560 233938 281616
rect 233790 279384 233846 279440
rect 233606 275032 233662 275088
rect 234250 372136 234306 372192
rect 234158 278296 234214 278352
rect 234066 273944 234122 274000
rect 234618 384920 234674 384976
rect 235814 384784 235870 384840
rect 235814 377848 235870 377904
rect 235630 377712 235686 377768
rect 234618 375400 234674 375456
rect 234434 375264 234490 375320
rect 235538 373904 235594 373960
rect 234526 368056 234582 368112
rect 234342 277208 234398 277264
rect 234250 272856 234306 272912
rect 235078 363976 235134 364032
rect 235446 362616 235502 362672
rect 235078 355136 235134 355192
rect 235078 352824 235134 352880
rect 234986 349152 235042 349208
rect 235262 353640 235318 353696
rect 235170 276120 235226 276176
rect 235078 270680 235134 270736
rect 235354 353232 235410 353288
rect 235262 261976 235318 262032
rect 235722 376624 235778 376680
rect 235630 269592 235686 269648
rect 235722 267416 235778 267472
rect 235538 266328 235594 266384
rect 235446 264152 235502 264208
rect 237286 380704 237342 380760
rect 236734 374584 236790 374640
rect 236182 372408 236238 372464
rect 236642 354184 236698 354240
rect 236550 354048 236606 354104
rect 235998 344392 236054 344448
rect 236366 343712 236422 343768
rect 235998 342080 236054 342136
rect 235906 265240 235962 265296
rect 235814 263064 235870 263120
rect 235354 260888 235410 260944
rect 234526 259800 234582 259856
rect 233974 254360 234030 254416
rect 236550 303320 236606 303376
rect 236826 372680 236882 372736
rect 236734 319776 236790 319832
rect 237194 365472 237250 365528
rect 237102 355000 237158 355056
rect 237010 354456 237066 354512
rect 237102 354320 237158 354376
rect 237010 341672 237066 341728
rect 236826 305496 236882 305552
rect 236642 302232 236698 302288
rect 236366 253272 236422 253328
rect 237102 323040 237158 323096
rect 238666 388456 238722 388512
rect 238482 388320 238538 388376
rect 237930 369008 237986 369064
rect 238298 363704 238354 363760
rect 237838 340176 237894 340232
rect 237746 327392 237802 327448
rect 237746 326440 237802 326496
rect 237838 323584 237894 323640
rect 237746 296792 237802 296848
rect 238206 355408 238262 355464
rect 238114 354864 238170 354920
rect 238022 325216 238078 325272
rect 238114 324128 238170 324184
rect 237930 321408 237986 321464
rect 238206 317600 238262 317656
rect 238022 317328 238078 317384
rect 238390 355972 238446 356008
rect 238390 355952 238392 355972
rect 238392 355952 238444 355972
rect 238444 355952 238446 355972
rect 238298 314336 238354 314392
rect 238022 297880 238078 297936
rect 237838 294616 237894 294672
rect 238574 379072 238630 379128
rect 238574 315424 238630 315480
rect 238574 313928 238630 313984
rect 238482 308760 238538 308816
rect 238390 280472 238446 280528
rect 237286 271768 237342 271824
rect 237194 268504 237250 268560
rect 237010 251096 237066 251152
rect 236918 250008 236974 250064
rect 233882 241304 233938 241360
rect 237378 236000 237434 236056
rect 238206 229336 238262 229392
rect 233882 202136 233938 202192
rect 233882 193432 233938 193488
rect 233146 150048 233202 150104
rect 233422 104352 233478 104408
rect 228362 101496 228418 101552
rect 229834 3848 229890 3904
rect 235906 172760 235962 172816
rect 235722 156576 235778 156632
rect 235354 153176 235410 153232
rect 235262 136856 235318 136912
rect 235814 155896 235870 155952
rect 235722 140256 235778 140312
rect 235354 120400 235410 120456
rect 238114 228248 238170 228304
rect 238022 227160 238078 227216
rect 237470 217368 237526 217424
rect 237378 216280 237434 216336
rect 237378 215328 237434 215384
rect 237470 197920 237526 197976
rect 239678 382200 239734 382256
rect 239494 361120 239550 361176
rect 239402 355272 239458 355328
rect 239402 354592 239458 354648
rect 239218 341400 239274 341456
rect 239218 339088 239274 339144
rect 239402 321952 239458 322008
rect 239678 354320 239734 354376
rect 239494 316512 239550 316568
rect 239310 313928 239366 313984
rect 239586 304408 239642 304464
rect 239770 339360 239826 339416
rect 239770 338680 239826 338736
rect 239678 300056 239734 300112
rect 238666 289176 238722 289232
rect 239770 252184 239826 252240
rect 238574 226344 238630 226400
rect 238298 226072 238354 226128
rect 238206 196560 238262 196616
rect 238114 193976 238170 194032
rect 238022 192616 238078 192672
rect 238206 187856 238262 187912
rect 238022 185000 238078 185056
rect 238114 181464 238170 181520
rect 238022 173848 238078 173904
rect 237378 155352 237434 155408
rect 237378 154264 237434 154320
rect 237286 152088 237342 152144
rect 238022 123528 238078 123584
rect 235814 120808 235870 120864
rect 235906 120672 235962 120728
rect 235722 120536 235778 120592
rect 235814 120264 235870 120320
rect 237286 120264 237342 120320
rect 237562 120264 237618 120320
rect 235906 119176 235962 119232
rect 235814 118904 235870 118960
rect 235262 118768 235318 118824
rect 237378 117816 237434 117872
rect 237470 117680 237526 117736
rect 237562 117408 237618 117464
rect 234618 117272 234674 117328
rect 234618 115232 234674 115288
rect 233882 17448 233938 17504
rect 237010 7656 237066 7712
rect 238574 216280 238630 216336
rect 238482 187720 238538 187776
rect 238298 185680 238354 185736
rect 238482 158616 238538 158672
rect 238390 156440 238446 156496
rect 238482 139032 238538 139088
rect 238390 137944 238446 138000
rect 238298 119992 238354 120048
rect 238666 215192 238722 215248
rect 238666 187856 238722 187912
rect 238666 173848 238722 173904
rect 238574 119468 238630 119504
rect 238574 119448 238576 119468
rect 238576 119448 238628 119468
rect 238628 119448 238630 119468
rect 239862 147804 239918 147860
rect 239862 146716 239918 146772
rect 240046 381112 240102 381168
rect 240046 353368 240102 353424
rect 240046 341672 240102 341728
rect 242990 359488 243046 359544
rect 241426 340040 241482 340096
rect 241610 340040 241666 340096
rect 243542 346976 243598 347032
rect 244094 346976 244150 347032
rect 243174 344392 243230 344448
rect 243542 343712 243598 343768
rect 244278 345752 244334 345808
rect 244830 345072 244886 345128
rect 244278 343576 244334 343632
rect 245750 357856 245806 357912
rect 244922 342896 244978 342952
rect 247590 359216 247646 359272
rect 246762 358536 246818 358592
rect 246670 357584 246726 357640
rect 248510 360032 248566 360088
rect 248326 348472 248382 348528
rect 249430 359896 249486 359952
rect 249706 349016 249762 349072
rect 251914 360712 251970 360768
rect 252190 359760 252246 359816
rect 251270 358944 251326 359000
rect 251086 344664 251142 344720
rect 250166 344256 250222 344312
rect 252374 359624 252430 359680
rect 252650 359624 252706 359680
rect 252466 359080 252522 359136
rect 252650 358944 252706 359000
rect 253110 345888 253166 345944
rect 254950 357312 255006 357368
rect 254030 356496 254086 356552
rect 253662 345752 253718 345808
rect 255318 344936 255374 344992
rect 255870 357176 255926 357232
rect 255410 343168 255466 343224
rect 256790 357040 256846 357096
rect 256698 341944 256754 342000
rect 257710 356904 257766 356960
rect 257158 341808 257214 341864
rect 258630 356768 258686 356824
rect 259550 356632 259606 356688
rect 258906 348744 258962 348800
rect 259366 348336 259422 348392
rect 259642 348744 259698 348800
rect 259642 348336 259698 348392
rect 262402 387096 262458 387152
rect 263230 380568 263286 380624
rect 262954 359760 263010 359816
rect 262678 359624 262734 359680
rect 260654 345888 260710 345944
rect 260746 345072 260802 345128
rect 265898 386280 265954 386336
rect 265070 385872 265126 385928
rect 264150 373360 264206 373416
rect 264150 365064 264206 365120
rect 266910 382064 266966 382120
rect 266358 380976 266414 381032
rect 265990 363840 266046 363896
rect 266358 346432 266414 346488
rect 268750 357720 268806 357776
rect 267830 355680 267886 355736
rect 267646 347384 267702 347440
rect 268382 340312 268438 340368
rect 268382 339904 268438 339960
rect 269026 354864 269082 354920
rect 269670 358264 269726 358320
rect 269394 341672 269450 341728
rect 270590 358128 270646 358184
rect 270406 341264 270462 341320
rect 272890 387640 272946 387696
rect 271786 358692 271842 358728
rect 271786 358672 271788 358692
rect 271788 358672 271840 358692
rect 271840 358672 271842 358692
rect 271786 358400 271842 358456
rect 271510 357992 271566 358048
rect 271142 344528 271198 344584
rect 271786 344120 271842 344176
rect 276018 372680 276074 372736
rect 274638 346024 274694 346080
rect 274638 345636 274694 345672
rect 274638 345616 274640 345636
rect 274640 345616 274692 345636
rect 274692 345616 274694 345636
rect 277030 373632 277086 373688
rect 276662 371184 276718 371240
rect 276386 355952 276442 356008
rect 276018 355000 276074 355056
rect 279606 387640 279662 387696
rect 279422 386960 279478 387016
rect 280066 387096 280122 387152
rect 250994 339496 251050 339552
rect 275742 339496 275798 339552
rect 279514 343712 279570 343768
rect 283378 386824 283434 386880
rect 282182 385600 282238 385656
rect 281630 384784 281686 384840
rect 282090 383696 282146 383752
rect 280894 373360 280950 373416
rect 280802 369008 280858 369064
rect 280434 351328 280490 351384
rect 280158 345616 280214 345672
rect 280066 339768 280122 339824
rect 250902 339360 250958 339416
rect 274638 339360 274694 339416
rect 278410 339360 278466 339416
rect 279974 339396 279976 339416
rect 279976 339396 280028 339416
rect 280028 339396 280030 339416
rect 279974 339360 280030 339396
rect 280158 339360 280214 339416
rect 280066 339088 280122 339144
rect 280066 338408 280122 338464
rect 280066 338272 280122 338328
rect 280066 338000 280122 338056
rect 280158 337864 280214 337920
rect 280066 336640 280122 336696
rect 280158 336232 280214 336288
rect 280434 305496 280490 305552
rect 280342 304408 280398 304464
rect 280250 303864 280306 303920
rect 280710 308760 280766 308816
rect 280618 307128 280674 307184
rect 280526 302776 280582 302832
rect 280986 357584 281042 357640
rect 280894 317736 280950 317792
rect 281078 343984 281134 344040
rect 281262 338680 281318 338736
rect 281906 338816 281962 338872
rect 281906 338408 281962 338464
rect 281354 336096 281410 336152
rect 281170 335960 281226 336016
rect 281814 307708 281816 307728
rect 281816 307708 281868 307728
rect 281868 307708 281870 307728
rect 281814 307672 281870 307708
rect 280986 306856 281042 306912
rect 280802 301416 280858 301472
rect 281906 298424 281962 298480
rect 281814 292984 281870 293040
rect 281906 292440 281962 292496
rect 281906 290808 281962 290864
rect 281906 289720 281962 289776
rect 281998 287000 282054 287056
rect 282090 284824 282146 284880
rect 282366 371864 282422 371920
rect 282274 285368 282330 285424
rect 282182 281560 282238 281616
rect 284942 372272 284998 372328
rect 282642 362344 282698 362400
rect 282550 286456 282606 286512
rect 282458 283736 282514 283792
rect 282366 279928 282422 279984
rect 282918 357448 282974 357504
rect 284298 355000 284354 355056
rect 283102 351872 283158 351928
rect 282826 351056 282882 351112
rect 282918 349016 282974 349072
rect 282918 308216 282974 308272
rect 284758 349424 284814 349480
rect 283286 348608 283342 348664
rect 283194 306584 283250 306640
rect 283102 304952 283158 305008
rect 283010 302232 283066 302288
rect 283010 293528 283066 293584
rect 282826 282648 282882 282704
rect 282734 278840 282790 278896
rect 282642 277752 282698 277808
rect 282090 269068 282146 269104
rect 282090 269048 282092 269068
rect 282092 269048 282144 269068
rect 282144 269048 282146 269068
rect 280158 268504 280214 268560
rect 282826 267960 282882 268016
rect 282826 265240 282882 265296
rect 282826 264152 282882 264208
rect 282826 263064 282882 263120
rect 282734 262520 282790 262576
rect 282826 261976 282882 262032
rect 282826 259800 282882 259856
rect 282826 259256 282882 259312
rect 282642 258712 282698 258768
rect 282734 258168 282790 258224
rect 282826 257624 282882 257680
rect 282734 257080 282790 257136
rect 282826 256572 282828 256592
rect 282828 256572 282880 256592
rect 282880 256572 282882 256592
rect 282826 256536 282882 256572
rect 282642 255992 282698 256048
rect 282734 255448 282790 255504
rect 282826 254360 282882 254416
rect 282826 253816 282882 253872
rect 282642 253272 282698 253328
rect 282734 252728 282790 252784
rect 282826 252184 282882 252240
rect 282734 251640 282790 251696
rect 282826 251132 282828 251152
rect 282828 251132 282880 251152
rect 282880 251132 282882 251152
rect 282826 251096 282882 251132
rect 282734 250552 282790 250608
rect 282550 250008 282606 250064
rect 282826 248920 282882 248976
rect 282734 248376 282790 248432
rect 282642 247832 282698 247888
rect 282826 246744 282882 246800
rect 282826 237496 282882 237552
rect 281538 235900 281540 235920
rect 281540 235900 281592 235920
rect 281592 235900 281594 235920
rect 281538 235864 281594 235900
rect 280250 229336 280306 229392
rect 280158 223352 280214 223408
rect 280066 192888 280122 192944
rect 280066 135088 280122 135144
rect 280066 134680 280122 134736
rect 238850 119312 238906 119368
rect 238850 118768 238906 118824
rect 238666 118632 238722 118688
rect 279974 120264 280030 120320
rect 279698 120128 279754 120184
rect 240506 116184 240562 116240
rect 238114 6296 238170 6352
rect 241426 116900 241428 116920
rect 241428 116900 241480 116920
rect 241480 116900 241482 116920
rect 241426 116864 241482 116900
rect 247774 118224 247830 118280
rect 247038 117544 247094 117600
rect 243358 106936 243414 106992
rect 251362 117952 251418 118008
rect 251178 113600 251234 113656
rect 240874 100000 240930 100056
rect 242070 6160 242126 6216
rect 247682 3848 247738 3904
rect 247590 3712 247646 3768
rect 244094 3576 244150 3632
rect 252466 113192 252522 113248
rect 254030 36624 254086 36680
rect 261758 117680 261814 117736
rect 255226 35264 255282 35320
rect 257618 33904 257674 33960
rect 261206 31048 261262 31104
rect 260010 26968 260066 27024
rect 258814 25608 258870 25664
rect 256422 24248 256478 24304
rect 252834 22888 252890 22944
rect 258262 3984 258318 4040
rect 254674 3848 254730 3904
rect 265346 117952 265402 118008
rect 264978 117408 265034 117464
rect 262402 28328 262458 28384
rect 264794 29824 264850 29880
rect 263598 6432 263654 6488
rect 271786 118360 271842 118416
rect 271142 117272 271198 117328
rect 270866 104216 270922 104272
rect 265990 98912 266046 98968
rect 268382 102856 268438 102912
rect 269578 97280 269634 97336
rect 267186 95784 267242 95840
rect 272890 117272 272946 117328
rect 273902 117272 273958 117328
rect 272062 105576 272118 105632
rect 277674 118088 277730 118144
rect 279422 118088 279478 118144
rect 276386 117272 276442 117328
rect 273902 93064 273958 93120
rect 275558 91704 275614 91760
rect 274362 90480 274418 90536
rect 271142 89120 271198 89176
rect 275282 85992 275338 86048
rect 271142 85856 271198 85912
rect 267002 54440 267058 54496
rect 268842 49272 268898 49328
rect 267002 6160 267058 6216
rect 278042 69400 278098 69456
rect 271142 3576 271198 3632
rect 270590 3440 270646 3496
rect 271050 3440 271106 3496
rect 272430 3576 272486 3632
rect 271786 2760 271842 2816
rect 278042 5616 278098 5672
rect 279514 4800 279570 4856
rect 279422 3304 279478 3360
rect 282550 228792 282606 228848
rect 281538 228248 281594 228304
rect 280342 226072 280398 226128
rect 280250 117680 280306 117736
rect 280526 222264 280582 222320
rect 280434 220632 280490 220688
rect 280342 116184 280398 116240
rect 280618 221720 280674 221776
rect 280894 218456 280950 218512
rect 280710 216280 280766 216336
rect 280618 116320 280674 116376
rect 280526 114960 280582 115016
rect 280802 214512 280858 214568
rect 280710 114416 280766 114472
rect 280434 112648 280490 112704
rect 280158 111424 280214 111480
rect 281630 227160 281686 227216
rect 281538 214512 281594 214568
rect 281998 226616 282054 226672
rect 281814 219000 281870 219056
rect 281722 217912 281778 217968
rect 280894 116728 280950 116784
rect 280802 3848 280858 3904
rect 281630 203224 281686 203280
rect 281906 217368 281962 217424
rect 282090 224440 282146 224496
rect 281998 120128 282054 120184
rect 282274 216824 282330 216880
rect 282182 215192 282238 215248
rect 282090 118224 282146 118280
rect 282366 198328 282422 198384
rect 282274 115096 282330 115152
rect 282182 112784 282238 112840
rect 281906 111288 281962 111344
rect 281814 109928 281870 109984
rect 281722 101632 281778 101688
rect 282734 215736 282790 215792
rect 282550 197376 282606 197432
rect 282642 167864 282698 167920
rect 282458 167320 282514 167376
rect 282642 162968 282698 163024
rect 282642 161880 282698 161936
rect 282366 100136 282422 100192
rect 281630 87488 281686 87544
rect 282182 84768 282238 84824
rect 280986 3712 281042 3768
rect 282918 197376 282974 197432
rect 282826 192344 282882 192400
rect 282826 170584 282882 170640
rect 282826 168428 282882 168464
rect 282826 168408 282828 168428
rect 282828 168408 282880 168428
rect 282880 168408 282882 168428
rect 282826 166776 282882 166832
rect 282826 165144 282882 165200
rect 282826 163512 282882 163568
rect 282826 162424 282882 162480
rect 282826 161372 282828 161392
rect 282828 161372 282880 161392
rect 282880 161372 282882 161392
rect 282826 161336 282882 161372
rect 282734 79464 282790 79520
rect 283194 291896 283250 291952
rect 283102 290264 283158 290320
rect 284298 348880 284354 348936
rect 284666 348200 284722 348256
rect 283654 347248 283710 347304
rect 283470 342624 283526 342680
rect 283562 306040 283618 306096
rect 283562 295296 283618 295352
rect 283470 266328 283526 266384
rect 283378 260888 283434 260944
rect 283286 244568 283342 244624
rect 284298 345616 284354 345672
rect 283654 290536 283710 290592
rect 283562 236952 283618 237008
rect 283838 339360 283894 339416
rect 283838 338816 283894 338872
rect 284390 294616 284446 294672
rect 283562 219544 283618 219600
rect 283378 209752 283434 209808
rect 283286 179016 283342 179072
rect 283286 178608 283342 178664
rect 283286 169768 283342 169824
rect 283010 119584 283066 119640
rect 283102 6160 283158 6216
rect 282918 3984 282974 4040
rect 282182 3304 282238 3360
rect 280066 3168 280122 3224
rect 283470 209208 283526 209264
rect 283746 213016 283802 213072
rect 283654 193432 283710 193488
rect 283562 107072 283618 107128
rect 284390 120944 284446 121000
rect 284298 119992 284354 120048
rect 284942 285096 284998 285152
rect 286690 386824 286746 386880
rect 286506 384648 286562 384704
rect 286322 379208 286378 379264
rect 285218 347112 285274 347168
rect 285126 337320 285182 337376
rect 285310 344528 285366 344584
rect 285402 341672 285458 341728
rect 285310 322088 285366 322144
rect 285678 341128 285734 341184
rect 285954 342352 286010 342408
rect 285402 321000 285458 321056
rect 285218 289448 285274 289504
rect 285770 295704 285826 295760
rect 284758 242936 284814 242992
rect 284666 236408 284722 236464
rect 285034 227704 285090 227760
rect 284758 220088 284814 220144
rect 284666 203768 284722 203824
rect 283746 108296 283802 108352
rect 283654 88984 283710 89040
rect 283470 77832 283526 77888
rect 283378 76472 283434 76528
rect 284850 213560 284906 213616
rect 284758 94696 284814 94752
rect 284942 210840 284998 210896
rect 285678 225528 285734 225584
rect 285126 221176 285182 221232
rect 285034 113600 285090 113656
rect 285126 108568 285182 108624
rect 284942 93200 284998 93256
rect 284850 91840 284906 91896
rect 284666 64096 284722 64152
rect 284942 43560 284998 43616
rect 285954 266872 286010 266928
rect 286230 229880 286286 229936
rect 285954 224984 286010 225040
rect 285862 212472 285918 212528
rect 285770 121080 285826 121136
rect 286138 223896 286194 223952
rect 286046 222808 286102 222864
rect 286414 365200 286470 365256
rect 286322 229608 286378 229664
rect 286782 345752 286838 345808
rect 286690 329704 286746 329760
rect 288162 386280 288218 386336
rect 288070 370912 288126 370968
rect 287702 355544 287758 355600
rect 287150 351464 287206 351520
rect 287058 349288 287114 349344
rect 286874 337456 286930 337512
rect 286782 311208 286838 311264
rect 286506 248104 286562 248160
rect 287150 295296 287206 295352
rect 287150 295160 287206 295216
rect 287058 242392 287114 242448
rect 286414 219816 286470 219872
rect 286414 211928 286470 211984
rect 286322 211384 286378 211440
rect 286230 117952 286286 118008
rect 286506 205400 286562 205456
rect 287058 201048 287114 201104
rect 286506 116456 286562 116512
rect 286414 114008 286470 114064
rect 286322 109792 286378 109848
rect 286138 108432 286194 108488
rect 286046 105712 286102 105768
rect 285954 104352 286010 104408
rect 285862 73752 285918 73808
rect 285678 7656 285734 7712
rect 286598 5616 286654 5672
rect 284942 3576 284998 3632
rect 283286 3440 283342 3496
rect 287610 206488 287666 206544
rect 287518 204312 287574 204368
rect 287426 202680 287482 202736
rect 287334 201592 287390 201648
rect 287242 200504 287298 200560
rect 287150 119040 287206 119096
rect 287886 349696 287942 349752
rect 287702 198056 287758 198112
rect 288254 341808 288310 341864
rect 288162 318824 288218 318880
rect 288254 313384 288310 313440
rect 288070 263336 288126 263392
rect 287886 215464 287942 215520
rect 287886 202136 287942 202192
rect 288530 349560 288586 349616
rect 289174 381792 289230 381848
rect 288622 337864 288678 337920
rect 288530 247288 288586 247344
rect 288714 208120 288770 208176
rect 288622 207576 288678 207632
rect 288530 207032 288586 207088
rect 287886 112512 287942 112568
rect 287610 111016 287666 111072
rect 287518 105440 287574 105496
rect 287426 72392 287482 72448
rect 289450 352688 289506 352744
rect 289174 236136 289230 236192
rect 290094 348064 290150 348120
rect 290002 338000 290058 338056
rect 292118 384784 292174 384840
rect 292026 383288 292082 383344
rect 291842 380432 291898 380488
rect 290738 375264 290794 375320
rect 290462 373768 290518 373824
rect 290370 334056 290426 334112
rect 290186 299376 290242 299432
rect 290094 260344 290150 260400
rect 290002 246200 290058 246256
rect 289450 218728 289506 218784
rect 289910 214104 289966 214160
rect 288898 196152 288954 196208
rect 288806 195064 288862 195120
rect 289082 195608 289138 195664
rect 288990 194520 289046 194576
rect 288898 102720 288954 102776
rect 290462 240488 290518 240544
rect 290738 299240 290794 299296
rect 291382 301144 291438 301200
rect 291290 294072 291346 294128
rect 291474 199416 291530 199472
rect 291382 131144 291438 131200
rect 291290 119312 291346 119368
rect 289910 114144 289966 114200
rect 289082 106800 289138 106856
rect 288990 101360 289046 101416
rect 288806 90344 288862 90400
rect 288714 61376 288770 61432
rect 288622 60016 288678 60072
rect 288530 58656 288586 58712
rect 287702 55664 287758 55720
rect 287334 50224 287390 50280
rect 287242 46144 287298 46200
rect 287058 4936 287114 4992
rect 291934 370776 291990 370832
rect 294694 383016 294750 383072
rect 293222 377576 293278 377632
rect 292302 345888 292358 345944
rect 292210 344392 292266 344448
rect 292118 328616 292174 328672
rect 292302 315560 292358 315616
rect 292210 304680 292266 304736
rect 292026 267688 292082 267744
rect 291934 232872 291990 232928
rect 291842 196968 291898 197024
rect 291566 170040 291622 170096
rect 291842 160656 291898 160712
rect 291842 153176 291898 153232
rect 291566 118768 291622 118824
rect 291842 118088 291898 118144
rect 291842 100544 291898 100600
rect 291474 49136 291530 49192
rect 289082 42200 289138 42256
rect 287702 4800 287758 4856
rect 290186 19896 290242 19952
rect 289082 3440 289138 3496
rect 293498 362888 293554 362944
rect 293406 349968 293462 350024
rect 294142 342216 294198 342272
rect 293958 298968 294014 299024
rect 293498 284008 293554 284064
rect 293406 262248 293462 262304
rect 293222 233960 293278 234016
rect 292762 210296 292818 210352
rect 293958 125432 294014 125488
rect 294234 341400 294290 341456
rect 294142 267416 294198 267472
rect 294234 265784 294290 265840
rect 294142 205944 294198 206000
rect 292762 113872 292818 113928
rect 294878 377984 294934 378040
rect 294694 238312 294750 238368
rect 294970 372408 295026 372464
rect 295062 346024 295118 346080
rect 295062 324264 295118 324320
rect 294970 300328 295026 300384
rect 294878 266600 294934 266656
rect 295430 337864 295486 337920
rect 295430 332968 295486 333024
rect 295430 299512 295486 299568
rect 296166 381928 296222 381984
rect 295982 376488 296038 376544
rect 295798 336232 295854 336288
rect 295798 263608 295854 263664
rect 295982 241576 296038 241632
rect 296258 352416 296314 352472
rect 296258 297064 296314 297120
rect 296166 265512 296222 265568
rect 296994 345208 297050 345264
rect 296994 269592 297050 269648
rect 297454 369280 297510 369336
rect 298742 367648 298798 367704
rect 298098 349152 298154 349208
rect 297546 339088 297602 339144
rect 297546 326440 297602 326496
rect 297454 274216 297510 274272
rect 299018 366696 299074 366752
rect 298926 365336 298982 365392
rect 298742 227432 298798 227488
rect 299018 286184 299074 286240
rect 298926 249192 298982 249248
rect 300122 385736 300178 385792
rect 299202 343168 299258 343224
rect 299202 312296 299258 312352
rect 299662 336096 299718 336152
rect 300490 364248 300546 364304
rect 300306 361392 300362 361448
rect 300214 349832 300270 349888
rect 300582 347384 300638 347440
rect 300582 319912 300638 319968
rect 304354 389000 304410 389056
rect 301594 372000 301650 372056
rect 301502 352960 301558 353016
rect 301134 350512 301190 350568
rect 300858 299376 300914 299432
rect 300490 294888 300546 294944
rect 301134 264696 301190 264752
rect 300306 251368 300362 251424
rect 301594 268776 301650 268832
rect 301502 245928 301558 245984
rect 300214 231784 300270 231840
rect 300122 213288 300178 213344
rect 298742 187720 298798 187776
rect 302606 350648 302662 350704
rect 304262 380296 304318 380352
rect 303250 369416 303306 369472
rect 302974 366288 303030 366344
rect 302606 261432 302662 261488
rect 303158 364112 303214 364168
rect 302974 228520 303030 228576
rect 303250 292712 303306 292768
rect 303158 252456 303214 252512
rect 303526 191664 303582 191720
rect 303526 187720 303582 187776
rect 304170 337456 304226 337512
rect 304170 331880 304226 331936
rect 305734 379344 305790 379400
rect 304446 362480 304502 362536
rect 304262 199144 304318 199200
rect 304998 350920 305054 350976
rect 304998 254904 305054 254960
rect 304446 253544 304502 253600
rect 305918 371048 305974 371104
rect 305734 258984 305790 259040
rect 307022 386008 307078 386064
rect 306378 350784 306434 350840
rect 305918 295976 305974 296032
rect 307206 374992 307262 375048
rect 307022 237224 307078 237280
rect 306378 232600 306434 232656
rect 307206 264424 307262 264480
rect 308586 351192 308642 351248
rect 309874 375808 309930 375864
rect 308586 278568 308642 278624
rect 309046 195880 309102 195936
rect 309046 191800 309102 191856
rect 308402 169768 308458 169824
rect 304354 167592 304410 167648
rect 308402 162832 308458 162888
rect 303986 162696 304042 162752
rect 303986 160792 304042 160848
rect 312542 386280 312598 386336
rect 311438 365608 311494 365664
rect 309874 275304 309930 275360
rect 310426 337320 310482 337376
rect 310426 330792 310482 330848
rect 310518 175208 310574 175264
rect 310426 169768 310482 169824
rect 298742 160248 298798 160304
rect 312542 302776 312598 302832
rect 311438 279656 311494 279712
rect 314198 367920 314254 367976
rect 315394 373496 315450 373552
rect 314198 256808 314254 256864
rect 318062 388864 318118 388920
rect 321834 390088 321890 390144
rect 315486 350104 315542 350160
rect 318154 384512 318210 384568
rect 315486 291624 315542 291680
rect 315394 202408 315450 202464
rect 315394 188400 315450 188456
rect 315394 175344 315450 175400
rect 316774 198736 316830 198792
rect 316774 188400 316830 188456
rect 321098 382200 321154 382256
rect 320914 380840 320970 380896
rect 318246 361528 318302 361584
rect 319626 368192 319682 368248
rect 318246 282784 318302 282840
rect 318154 242664 318210 242720
rect 318154 208528 318210 208584
rect 318338 208392 318394 208448
rect 318338 198736 318394 198792
rect 318154 196016 318210 196072
rect 318062 148416 318118 148472
rect 316682 148280 316738 148336
rect 297362 147328 297418 147384
rect 295614 146920 295670 146976
rect 295982 146920 296038 146976
rect 295430 120536 295486 120592
rect 319626 280744 319682 280800
rect 319626 255312 319682 255368
rect 320546 212472 320602 212528
rect 320914 273128 320970 273184
rect 320914 263608 320970 263664
rect 320914 255312 320970 255368
rect 322386 386144 322442 386200
rect 321098 302504 321154 302560
rect 320546 208528 320602 208584
rect 319626 208392 319682 208448
rect 320822 190712 320878 190768
rect 294142 113736 294198 113792
rect 323674 366560 323730 366616
rect 322386 288360 322442 288416
rect 322294 230424 322350 230480
rect 322294 212472 322350 212528
rect 323766 340040 323822 340096
rect 323766 303456 323822 303512
rect 323674 257896 323730 257952
rect 323674 252184 323730 252240
rect 323674 230424 323730 230480
rect 329102 353096 329158 353152
rect 327814 348472 327870 348528
rect 325882 272992 325938 273048
rect 325146 263608 325202 263664
rect 326986 253816 327042 253872
rect 326986 252184 327042 252240
rect 327814 307944 327870 308000
rect 327814 288224 327870 288280
rect 331862 339496 331918 339552
rect 329930 291080 329986 291136
rect 329930 288224 329986 288280
rect 330482 282240 330538 282296
rect 329102 277480 329158 277536
rect 329102 274624 329158 274680
rect 330482 274624 330538 274680
rect 327814 272992 327870 273048
rect 329102 253816 329158 253872
rect 323582 148552 323638 148608
rect 320822 97824 320878 97880
rect 304354 86128 304410 86184
rect 297270 32544 297326 32600
rect 293682 3576 293738 3632
rect 300766 3440 300822 3496
rect 322110 85720 322166 85776
rect 311438 82048 311494 82104
rect 307114 59880 307170 59936
rect 307114 53216 307170 53272
rect 307942 53080 307998 53136
rect 318522 80688 318578 80744
rect 315026 51720 315082 51776
rect 329194 79328 329250 79384
rect 324962 58520 325018 58576
rect 324962 7656 325018 7712
rect 325606 7520 325662 7576
rect 332046 300736 332102 300792
rect 331954 292576 332010 292632
rect 332046 291080 332102 291136
rect 331954 282240 332010 282296
rect 333518 343032 333574 343088
rect 333518 300736 333574 300792
rect 334714 342896 334770 342952
rect 334806 306448 334862 306504
rect 334714 305768 334770 305824
rect 334806 292576 334862 292632
rect 336094 177792 336150 177848
rect 336370 180376 336426 180432
rect 337382 347112 337438 347168
rect 336646 338816 336702 338872
rect 336646 327528 336702 327584
rect 337382 306448 337438 306504
rect 339406 345072 339462 345128
rect 339406 343032 339462 343088
rect 339130 302776 339186 302832
rect 338946 179016 339002 179072
rect 341614 363568 341670 363624
rect 346306 387912 346362 387968
rect 349802 388048 349858 388104
rect 341890 179288 341946 179344
rect 346214 349832 346270 349888
rect 346214 345072 346270 345128
rect 345662 344256 345718 344312
rect 345662 309032 345718 309088
rect 341614 176568 341670 176624
rect 347594 352552 347650 352608
rect 353298 387368 353354 387424
rect 351550 387232 351606 387288
rect 350078 386960 350134 387016
rect 353942 386960 353998 387016
rect 350446 360712 350502 360768
rect 347594 180240 347650 180296
rect 349894 178880 349950 178936
rect 351182 348336 351238 348392
rect 351182 314472 351238 314528
rect 350446 310120 350502 310176
rect 349802 177520 349858 177576
rect 353298 349696 353354 349752
rect 353298 347112 353354 347168
rect 339130 151136 339186 151192
rect 355966 383968 356022 384024
rect 355690 181736 355746 181792
rect 355506 177656 355562 177712
rect 355874 173168 355930 173224
rect 357346 387232 357402 387288
rect 357346 383832 357402 383888
rect 357254 347792 357310 347848
rect 358266 373088 358322 373144
rect 357254 299376 357310 299432
rect 352562 147600 352618 147656
rect 353942 147600 353998 147656
rect 350078 147056 350134 147112
rect 355322 146648 355378 146704
rect 352746 146512 352802 146568
rect 352930 146376 352986 146432
rect 352746 115640 352802 115696
rect 352562 115504 352618 115560
rect 355506 144336 355562 144392
rect 355966 147328 356022 147384
rect 357530 287816 357586 287872
rect 357530 282240 357586 282296
rect 357530 276800 357586 276856
rect 357530 272584 357586 272640
rect 357530 271360 357586 271416
rect 357530 270136 357586 270192
rect 357530 261568 357586 261624
rect 357530 256128 357586 256184
rect 357530 254904 357586 254960
rect 357530 250688 357586 250744
rect 357530 246880 357586 246936
rect 357530 245112 357586 245168
rect 357530 243888 357586 243944
rect 357530 239672 357586 239728
rect 357530 235456 357586 235512
rect 357530 231240 357586 231296
rect 357530 226228 357586 226264
rect 357530 226208 357532 226228
rect 357532 226208 357584 226228
rect 357584 226208 357586 226228
rect 357714 225664 357770 225720
rect 357530 224440 357586 224496
rect 357530 223216 357586 223272
rect 357530 222028 357532 222048
rect 357532 222028 357584 222048
rect 357584 222028 357586 222048
rect 357530 221992 357586 222028
rect 357714 221448 357770 221504
rect 357530 217776 357586 217832
rect 357530 216588 357532 216608
rect 357532 216588 357584 216608
rect 357584 216588 357586 216608
rect 357530 216552 357586 216588
rect 357530 214784 357586 214840
rect 357530 212336 357586 212392
rect 357530 211132 357586 211168
rect 357530 211112 357532 211132
rect 357532 211112 357584 211132
rect 357584 211112 357586 211132
rect 357530 209344 357586 209400
rect 357530 207984 357586 208040
rect 357530 206760 357586 206816
rect 357530 206216 357586 206272
rect 357530 204992 357586 205048
rect 357530 203768 357586 203824
rect 357530 201320 357586 201376
rect 357530 200776 357586 200832
rect 357530 195916 357532 195936
rect 357532 195916 357584 195936
rect 357584 195916 357586 195936
rect 357530 195880 357586 195916
rect 358450 355952 358506 356008
rect 358266 298696 358322 298752
rect 360014 387368 360070 387424
rect 359646 386688 359702 386744
rect 358726 351872 358782 351928
rect 358634 338680 358690 338736
rect 358542 335960 358598 336016
rect 358450 325488 358506 325544
rect 358634 323720 358690 323776
rect 358542 317192 358598 317248
rect 358358 293800 358414 293856
rect 358174 177928 358230 177984
rect 359554 180512 359610 180568
rect 359830 387096 359886 387152
rect 360014 386552 360070 386608
rect 359830 346976 359886 347032
rect 359922 180104 359978 180160
rect 358726 172488 358782 172544
rect 360014 171672 360070 171728
rect 360198 386452 360200 386472
rect 360200 386452 360252 386472
rect 360252 386452 360254 386472
rect 360198 386416 360254 386452
rect 362038 386824 362094 386880
rect 363786 386824 363842 386880
rect 369030 384104 369086 384160
rect 370778 368056 370834 368112
rect 367282 362752 367338 362808
rect 365534 359352 365590 359408
rect 372526 355136 372582 355192
rect 376022 377848 376078 377904
rect 379518 384920 379574 384976
rect 383014 376624 383070 376680
rect 381266 373904 381322 373960
rect 386510 377712 386566 377768
rect 384762 365472 384818 365528
rect 377770 362616 377826 362672
rect 374274 353640 374330 353696
rect 390006 380704 390062 380760
rect 391754 372136 391810 372192
rect 395250 378528 395306 378584
rect 393502 369144 393558 369200
rect 398930 388728 398986 388784
rect 398838 387776 398894 387832
rect 400218 388184 400274 388240
rect 400310 387912 400366 387968
rect 400218 387232 400274 387288
rect 398930 386960 398986 387016
rect 398746 381384 398802 381440
rect 400494 374856 400550 374912
rect 396998 363976 397054 364032
rect 403622 386960 403678 387016
rect 402242 361256 402298 361312
rect 404266 386552 404322 386608
rect 404266 386144 404322 386200
rect 405738 370640 405794 370696
rect 403622 357720 403678 357776
rect 407486 355816 407542 355872
rect 417974 387096 418030 387152
rect 416226 383152 416282 383208
rect 414478 377440 414534 377496
rect 412730 367784 412786 367840
rect 410982 366424 411038 366480
rect 421562 359352 421618 359408
rect 421470 357856 421526 357912
rect 409234 353776 409290 353832
rect 388258 352824 388314 352880
rect 401966 352688 402022 352744
rect 373998 351872 374054 351928
rect 426714 360032 426770 360088
rect 428462 359896 428518 359952
rect 431222 386008 431278 386064
rect 424966 359216 425022 359272
rect 423218 358536 423274 358592
rect 421562 352552 421618 352608
rect 431958 359760 432014 359816
rect 433706 359624 433762 359680
rect 438950 357312 439006 357368
rect 440698 357176 440754 357232
rect 442446 357040 442502 357096
rect 444194 356904 444250 356960
rect 445942 356768 445998 356824
rect 454682 380568 454738 380624
rect 458178 385872 458234 385928
rect 456430 365064 456486 365120
rect 461674 382064 461730 382120
rect 459926 363840 459982 363896
rect 447690 356632 447746 356688
rect 437202 356496 437258 356552
rect 460938 355952 460994 356008
rect 457902 352552 457958 352608
rect 429934 352008 429990 352064
rect 431222 352008 431278 352064
rect 465170 386960 465226 387016
rect 467838 360168 467894 360224
rect 466918 358264 466974 358320
rect 468666 358128 468722 358184
rect 471242 383152 471298 383208
rect 470414 357992 470470 358048
rect 467838 355952 467894 356008
rect 463422 355680 463478 355736
rect 473266 362072 473322 362128
rect 473266 360168 473322 360224
rect 476394 366968 476450 367024
rect 476394 362072 476450 362128
rect 478878 369824 478934 369880
rect 480902 387640 480958 387696
rect 478878 366968 478934 367024
rect 479522 362888 479578 362944
rect 471242 352552 471298 352608
rect 482282 372680 482338 372736
rect 482282 363160 482338 363216
rect 484398 387096 484454 387152
rect 486146 387232 486202 387288
rect 485870 386960 485926 387016
rect 485410 376624 485466 376680
rect 485778 375808 485834 375864
rect 485778 372680 485834 372736
rect 482834 371728 482890 371784
rect 485410 371728 485466 371784
rect 482834 369824 482890 369880
rect 482650 359488 482706 359544
rect 480902 359352 480958 359408
rect 476118 350648 476174 350704
rect 479522 350648 479578 350704
rect 460846 349832 460902 349888
rect 487894 384376 487950 384432
rect 491298 385872 491354 385928
rect 489642 384240 489698 384296
rect 491942 387368 491998 387424
rect 490930 380976 490986 381032
rect 487342 378528 487398 378584
rect 487250 377984 487306 378040
rect 499486 387368 499542 387424
rect 498106 385872 498162 385928
rect 497462 384240 497518 384296
rect 491942 380976 491998 381032
rect 491206 378528 491262 378584
rect 490930 377984 490986 378040
rect 487342 376624 487398 376680
rect 487250 375808 487306 375864
rect 485962 375400 486018 375456
rect 499946 388048 500002 388104
rect 499762 387096 499818 387152
rect 497462 352688 497518 352744
rect 476118 349696 476174 349752
rect 360474 345752 360530 345808
rect 387982 180512 388038 180568
rect 478050 180512 478106 180568
rect 392030 180376 392086 180432
rect 461858 180376 461914 180432
rect 405186 180240 405242 180296
rect 454774 180240 454830 180296
rect 372802 177928 372858 177984
rect 371790 177792 371846 177848
rect 374826 177656 374882 177712
rect 391018 176568 391074 176624
rect 407762 179832 407818 179888
rect 365718 173168 365774 173224
rect 357530 147056 357586 147112
rect 357346 146512 357402 146568
rect 355506 117000 355562 117056
rect 355322 115776 355378 115832
rect 358726 146956 358728 146976
rect 358728 146956 358780 146976
rect 358780 146956 358782 146976
rect 358726 146920 358782 146956
rect 358082 118632 358138 118688
rect 358542 144472 358598 144528
rect 364982 168952 365038 169008
rect 363602 166232 363658 166288
rect 369858 167592 369914 167648
rect 367466 147056 367522 147112
rect 407118 172488 407174 172544
rect 402978 171672 403034 171728
rect 375838 151136 375894 151192
rect 383014 148552 383070 148608
rect 379426 148416 379482 148472
rect 378230 148280 378286 148336
rect 394974 169088 395030 169144
rect 400954 147192 401010 147248
rect 399758 146648 399814 146704
rect 402150 146512 402206 146568
rect 402978 146376 403034 146432
rect 396170 144336 396226 144392
rect 352930 115368 352986 115424
rect 407210 144744 407266 144800
rect 410246 179288 410302 179344
rect 411258 179016 411314 179072
rect 415306 179288 415362 179344
rect 414294 178880 414350 178936
rect 413282 177520 413338 177576
rect 421378 180104 421434 180160
rect 420366 176568 420422 176624
rect 418342 175208 418398 175264
rect 424414 176024 424470 176080
rect 422390 175072 422446 175128
rect 425426 174936 425482 174992
rect 428462 174800 428518 174856
rect 433522 176296 433578 176352
rect 435546 176160 435602 176216
rect 438582 177248 438638 177304
rect 437570 176432 437626 176488
rect 432510 174664 432566 174720
rect 431498 174528 431554 174584
rect 441618 180104 441674 180160
rect 462870 179016 462926 179072
rect 457810 178880 457866 178936
rect 456798 178744 456854 178800
rect 474002 179696 474058 179752
rect 471978 177792 472034 177848
rect 481086 177520 481142 177576
rect 490194 177928 490250 177984
rect 487158 177656 487214 177712
rect 493230 177384 493286 177440
rect 499670 202680 499726 202736
rect 499762 179832 499818 179888
rect 439594 174392 439650 174448
rect 500866 521736 500922 521792
rect 500866 519832 500922 519888
rect 500866 519288 500922 519344
rect 500590 511808 500646 511864
rect 500590 488280 500646 488336
rect 500498 482296 500554 482352
rect 500498 474544 500554 474600
rect 500866 451152 500922 451208
rect 501142 442856 501198 442912
rect 501602 554512 501658 554568
rect 501510 523232 501566 523288
rect 501418 479848 501474 479904
rect 503166 598848 503222 598904
rect 504822 600072 504878 600128
rect 504546 598032 504602 598088
rect 505098 599528 505154 599584
rect 502338 552472 502394 552528
rect 502062 550976 502118 551032
rect 501970 522144 502026 522200
rect 501878 519152 501934 519208
rect 501602 483928 501658 483984
rect 501510 443672 501566 443728
rect 501326 443128 501382 443184
rect 501234 441496 501290 441552
rect 501050 438776 501106 438832
rect 500682 404912 500738 404968
rect 500590 391856 500646 391912
rect 500682 389000 500738 389056
rect 500498 388864 500554 388920
rect 500958 387232 501014 387288
rect 501050 360848 501106 360904
rect 501142 208256 501198 208312
rect 501234 196696 501290 196752
rect 501050 190304 501106 190360
rect 500958 181328 501014 181384
rect 501694 474544 501750 474600
rect 502246 520240 502302 520296
rect 502154 519016 502210 519072
rect 502246 511944 502302 512000
rect 503534 551112 503590 551168
rect 502522 547712 502578 547768
rect 502338 482024 502394 482080
rect 502338 481344 502394 481400
rect 502062 442584 502118 442640
rect 502614 543632 502670 543688
rect 502706 538600 502762 538656
rect 502798 534520 502854 534576
rect 502706 484472 502762 484528
rect 502706 483928 502762 483984
rect 502614 483656 502670 483712
rect 502522 483384 502578 483440
rect 502798 482840 502854 482896
rect 503074 525408 503130 525464
rect 503258 523368 503314 523424
rect 503166 520240 503222 520296
rect 503074 486376 503130 486432
rect 503166 485832 503222 485888
rect 502890 482568 502946 482624
rect 502890 469240 502946 469296
rect 502890 468424 502946 468480
rect 502798 468152 502854 468208
rect 502706 466792 502762 466848
rect 502890 467336 502946 467392
rect 502798 466520 502854 466576
rect 502890 466248 502946 466304
rect 502706 465976 502762 466032
rect 502798 465704 502854 465760
rect 502614 465432 502670 465488
rect 502890 464072 502946 464128
rect 502706 463256 502762 463312
rect 502890 462984 502946 463040
rect 502798 462712 502854 462768
rect 502614 462440 502670 462496
rect 502890 462204 502892 462224
rect 502892 462204 502944 462224
rect 502944 462204 502946 462224
rect 502890 462168 502946 462204
rect 502522 461896 502578 461952
rect 502614 461352 502670 461408
rect 502890 461624 502946 461680
rect 502798 461080 502854 461136
rect 502798 460536 502854 460592
rect 502890 460264 502946 460320
rect 502614 458904 502670 458960
rect 502890 459176 502946 459232
rect 502798 458632 502854 458688
rect 502706 458360 502762 458416
rect 502890 458088 502946 458144
rect 502798 457816 502854 457872
rect 502706 457272 502762 457328
rect 502614 457000 502670 457056
rect 502890 456728 502946 456784
rect 502890 456492 502892 456512
rect 502892 456492 502944 456512
rect 502944 456492 502946 456512
rect 502890 456456 502946 456492
rect 502798 455912 502854 455968
rect 502614 455640 502670 455696
rect 502798 455368 502854 455424
rect 502890 455116 502946 455152
rect 502890 455096 502892 455116
rect 502892 455096 502944 455116
rect 502944 455096 502946 455116
rect 502706 454824 502762 454880
rect 502614 454280 502670 454336
rect 502522 454008 502578 454064
rect 502890 453736 502946 453792
rect 502798 453192 502854 453248
rect 502706 452648 502762 452704
rect 502890 452412 502892 452432
rect 502892 452412 502944 452432
rect 502944 452412 502946 452432
rect 502890 452376 502946 452412
rect 502706 452104 502762 452160
rect 502798 451832 502854 451888
rect 502614 451560 502670 451616
rect 502706 450472 502762 450528
rect 502890 450200 502946 450256
rect 502614 449928 502670 449984
rect 502706 448840 502762 448896
rect 502890 449112 502946 449168
rect 502798 448568 502854 448624
rect 502890 448024 502946 448080
rect 502706 447752 502762 447808
rect 502614 447480 502670 447536
rect 502798 434152 502854 434208
rect 502614 432792 502670 432848
rect 502522 430888 502578 430944
rect 502706 430616 502762 430672
rect 502614 430072 502670 430128
rect 502522 428168 502578 428224
rect 502706 427624 502762 427680
rect 502798 427352 502854 427408
rect 502890 425448 502946 425504
rect 502614 423272 502670 423328
rect 502430 423000 502486 423056
rect 501970 390632 502026 390688
rect 502522 422728 502578 422784
rect 502706 422456 502762 422512
rect 502614 386960 502670 387016
rect 502522 386008 502578 386064
rect 502430 384240 502486 384296
rect 502706 383152 502762 383208
rect 502522 232872 502578 232928
rect 502798 250552 502854 250608
rect 502706 238312 502762 238368
rect 502614 226208 502670 226264
rect 502430 220768 502486 220824
rect 502338 214648 502394 214704
rect 503718 546488 503774 546544
rect 503718 523096 503774 523152
rect 503718 519596 503720 519616
rect 503720 519596 503772 519616
rect 503772 519596 503774 519616
rect 503718 519560 503774 519596
rect 503626 487464 503682 487520
rect 503626 484336 503682 484392
rect 503350 481752 503406 481808
rect 503258 480936 503314 480992
rect 503534 481344 503590 481400
rect 503626 451152 503682 451208
rect 503626 451052 503628 451072
rect 503628 451052 503680 451072
rect 503680 451052 503682 451072
rect 503626 451016 503682 451052
rect 503626 450744 503682 450800
rect 503626 449656 503682 449712
rect 503626 449384 503682 449440
rect 503626 448332 503628 448352
rect 503628 448332 503680 448352
rect 503680 448332 503682 448352
rect 503626 448296 503682 448332
rect 503626 445304 503682 445360
rect 503626 441768 503682 441824
rect 503626 440680 503682 440736
rect 503626 440172 503628 440192
rect 503628 440172 503680 440192
rect 503680 440172 503682 440192
rect 503626 440136 503682 440172
rect 503626 439864 503682 439920
rect 503626 437960 503682 438016
rect 503534 437688 503590 437744
rect 503626 437144 503682 437200
rect 503626 436872 503682 436928
rect 503626 435512 503682 435568
rect 503442 434696 503498 434752
rect 503626 434424 503682 434480
rect 503534 433880 503590 433936
rect 503442 433336 503498 433392
rect 503442 433064 503498 433120
rect 503534 432520 503590 432576
rect 503626 432248 503682 432304
rect 503442 431976 503498 432032
rect 504454 554376 504510 554432
rect 504178 536152 504234 536208
rect 504086 533296 504142 533352
rect 503994 452920 504050 452976
rect 504178 443944 504234 444000
rect 504086 439048 504142 439104
rect 504270 438504 504326 438560
rect 504638 552744 504694 552800
rect 504546 542272 504602 542328
rect 504638 520512 504694 520568
rect 504546 483112 504602 483168
rect 504454 479576 504510 479632
rect 504362 438232 504418 438288
rect 503902 433608 503958 433664
rect 503626 431740 503628 431760
rect 503628 431740 503680 431760
rect 503680 431740 503682 431760
rect 503626 431704 503682 431740
rect 503534 431432 503590 431488
rect 503442 431160 503498 431216
rect 503626 430344 503682 430400
rect 503626 429936 503682 429992
rect 503534 429528 503590 429584
rect 503442 429256 503498 429312
rect 503626 429020 503628 429040
rect 503628 429020 503680 429040
rect 503680 429020 503682 429040
rect 503626 428984 503682 429020
rect 503626 428712 503682 428768
rect 503626 428440 503682 428496
rect 503626 427896 503682 427952
rect 503442 426808 503498 426864
rect 503626 427080 503682 427136
rect 503534 426536 503590 426592
rect 503626 426300 503628 426320
rect 503628 426300 503680 426320
rect 503680 426300 503682 426320
rect 503626 426264 503682 426300
rect 503442 425720 503498 425776
rect 503534 425176 503590 425232
rect 503626 424904 503682 424960
rect 503626 424360 503682 424416
rect 503534 424088 503590 424144
rect 503442 423816 503498 423872
rect 503626 423580 503628 423600
rect 503628 423580 503680 423600
rect 503680 423580 503682 423600
rect 503626 423544 503682 423580
rect 505926 598032 505982 598088
rect 507306 598032 507362 598088
rect 507858 554784 507914 554840
rect 505098 387640 505154 387696
rect 504730 373632 504786 373688
rect 503626 346024 503682 346080
rect 503626 340312 503682 340368
rect 503626 333784 503682 333840
rect 503626 328072 503682 328128
rect 503626 322360 503682 322416
rect 503626 304408 503682 304464
rect 503626 297880 503682 297936
rect 503626 292168 503682 292224
rect 503626 286456 503682 286512
rect 503626 274216 503682 274272
rect 503626 184864 503682 184920
rect 503902 256672 503958 256728
rect 503810 244296 503866 244352
rect 506478 547848 506534 547904
rect 506478 541068 506534 541104
rect 506478 541048 506480 541068
rect 506480 541048 506532 541068
rect 506532 541048 506534 541068
rect 506018 519696 506074 519752
rect 505926 484336 505982 484392
rect 505834 480256 505890 480312
rect 505374 394576 505430 394632
rect 505374 390360 505430 390416
rect 507030 539960 507086 540016
rect 507306 530440 507362 530496
rect 507122 525000 507178 525056
rect 507306 472232 507362 472288
rect 507122 445848 507178 445904
rect 507030 445032 507086 445088
rect 507950 519696 508006 519752
rect 507950 519016 508006 519072
rect 508410 539008 508466 539064
rect 508410 447208 508466 447264
rect 508502 407768 508558 407824
rect 508502 394576 508558 394632
rect 507950 381656 508006 381712
rect 509698 552880 509754 552936
rect 509606 551248 509662 551304
rect 509238 550704 509294 550760
rect 508686 354048 508742 354104
rect 509422 519152 509478 519208
rect 509790 532752 509846 532808
rect 509698 477128 509754 477184
rect 509974 513440 510030 513496
rect 509606 440952 509662 441008
rect 509422 382880 509478 382936
rect 510710 519696 510766 519752
rect 510618 519288 510674 519344
rect 510894 548664 510950 548720
rect 510986 547168 511042 547224
rect 510986 441224 511042 441280
rect 510894 440408 510950 440464
rect 511998 559020 512054 559056
rect 511998 559000 512000 559020
rect 512000 559000 512052 559020
rect 512052 559000 512054 559020
rect 512090 545264 512146 545320
rect 511998 527176 512054 527232
rect 511998 524456 512054 524512
rect 511630 520512 511686 520568
rect 511538 519696 511594 519752
rect 511354 485288 511410 485344
rect 511354 481344 511410 481400
rect 510710 389816 510766 389872
rect 512274 544720 512330 544776
rect 512458 540232 512514 540288
rect 512366 532616 512422 532672
rect 512274 446664 512330 446720
rect 512090 439320 512146 439376
rect 512550 537512 512606 537568
rect 512734 534792 512790 534848
rect 512642 519016 512698 519072
rect 512642 486104 512698 486160
rect 512642 480800 512698 480856
rect 512550 446936 512606 446992
rect 512458 445576 512514 445632
rect 512366 437416 512422 437472
rect 512734 446392 512790 446448
rect 514758 532788 514760 532808
rect 514760 532788 514812 532808
rect 514812 532788 514814 532808
rect 514758 532752 514814 532788
rect 514022 529080 514078 529136
rect 514758 527176 514814 527232
rect 514206 525816 514262 525872
rect 514114 519832 514170 519888
rect 514758 520240 514814 520296
rect 514666 514664 514722 514720
rect 514666 505280 514722 505336
rect 514206 485560 514262 485616
rect 514114 476040 514170 476096
rect 514022 457544 514078 457600
rect 515402 558320 515458 558376
rect 515494 555464 515550 555520
rect 515402 471416 515458 471472
rect 515678 534928 515734 534984
rect 515494 471144 515550 471200
rect 515678 425992 515734 426048
rect 516690 530848 516746 530904
rect 516690 456184 516746 456240
rect 517518 527176 517574 527232
rect 517518 521736 517574 521792
rect 517058 521192 517114 521248
rect 516966 364928 517022 364984
rect 517886 536016 517942 536072
rect 518070 523096 518126 523152
rect 517886 424632 517942 424688
rect 518254 533704 518310 533760
rect 518254 526496 518310 526552
rect 518346 521464 518402 521520
rect 518346 469512 518402 469568
rect 518162 378936 518218 378992
rect 518990 532772 519046 532808
rect 518990 532752 518992 532772
rect 518992 532752 519044 532772
rect 519044 532752 519046 532772
rect 519450 543088 519506 543144
rect 519542 526360 519598 526416
rect 519726 523504 519782 523560
rect 519726 464344 519782 464400
rect 519542 446120 519598 446176
rect 519450 444216 519506 444272
rect 521658 539724 521660 539744
rect 521660 539724 521712 539744
rect 521712 539724 521714 539744
rect 521658 539688 521714 539724
rect 521658 539588 521660 539608
rect 521660 539588 521712 539608
rect 521712 539588 521714 539608
rect 521658 539552 521714 539588
rect 521106 535064 521162 535120
rect 520830 522688 520886 522744
rect 521658 531392 521714 531448
rect 521106 485016 521162 485072
rect 520830 435784 520886 435840
rect 522302 539280 522358 539336
rect 522026 538736 522082 538792
rect 522302 475496 522358 475552
rect 522026 439592 522082 439648
rect 523038 554784 523094 554840
rect 522486 363704 522542 363760
rect 523038 527212 523040 527232
rect 523040 527212 523092 527232
rect 523092 527212 523094 527232
rect 523038 527176 523094 527212
rect 523682 525680 523738 525736
rect 523590 522416 523646 522472
rect 523774 523640 523830 523696
rect 523774 468016 523830 468072
rect 523682 463528 523738 463584
rect 523590 436600 523646 436656
rect 523958 467880 524014 467936
rect 523866 379072 523922 379128
rect 525154 529352 525210 529408
rect 524786 522280 524842 522336
rect 525154 486920 525210 486976
rect 524786 436328 524842 436384
rect 525798 531392 525854 531448
rect 525798 523096 525854 523152
rect 525246 361120 525302 361176
rect 526442 530712 526498 530768
rect 526442 467608 526498 467664
rect 526626 355408 526682 355464
rect 527730 528128 527786 528184
rect 527730 463800 527786 463856
rect 528742 599936 528798 599992
rect 528650 598440 528706 598496
rect 528006 376352 528062 376408
rect 528742 390088 528798 390144
rect 528650 376216 528706 376272
rect 529846 597896 529902 597952
rect 529938 560360 529994 560416
rect 529846 531412 529902 531448
rect 529846 531392 529848 531412
rect 529848 531392 529900 531412
rect 529900 531392 529902 531412
rect 529386 374584 529442 374640
rect 529938 355952 529994 356008
rect 531318 597760 531374 597816
rect 531226 521600 531282 521656
rect 530582 181736 530638 181792
rect 531502 598304 531558 598360
rect 531870 528264 531926 528320
rect 531778 527856 531834 527912
rect 531962 527040 532018 527096
rect 532054 524048 532110 524104
rect 532054 486648 532110 486704
rect 531962 468968 532018 469024
rect 531870 464888 531926 464944
rect 531778 464616 531834 464672
rect 531502 377304 531558 377360
rect 532882 599800 532938 599856
rect 532698 598712 532754 598768
rect 532974 598304 533030 598360
rect 534078 598576 534134 598632
rect 533526 598032 533582 598088
rect 533066 533840 533122 533896
rect 533434 533160 533490 533216
rect 533066 460808 533122 460864
rect 533526 530576 533582 530632
rect 533434 468696 533490 468752
rect 533526 467064 533582 467120
rect 533342 427080 533398 427136
rect 533342 407768 533398 407824
rect 532882 404912 532938 404968
rect 535458 598848 535514 598904
rect 534906 598032 534962 598088
rect 534170 597760 534226 597816
rect 534262 559816 534318 559872
rect 535366 535508 535368 535528
rect 535368 535508 535420 535528
rect 535420 535508 535422 535528
rect 535366 535472 535422 535508
rect 534354 533432 534410 533488
rect 534262 480664 534318 480720
rect 534354 459720 534410 459776
rect 534814 527720 534870 527776
rect 534998 468424 535054 468480
rect 534814 465160 534870 465216
rect 534998 444760 535054 444816
rect 534170 378800 534226 378856
rect 534078 376080 534134 376136
rect 532698 375944 532754 376000
rect 535642 597624 535698 597680
rect 536930 598304 536986 598360
rect 535918 533976 535974 534032
rect 535918 459448 535974 459504
rect 535642 381520 535698 381576
rect 535458 373224 535514 373280
rect 532698 355952 532754 356008
rect 534078 355952 534134 356008
rect 536194 533568 536250 533624
rect 536378 460128 536434 460184
rect 536194 459992 536250 460048
rect 536378 427080 536434 427136
rect 532146 355272 532202 355328
rect 531410 347792 531466 347848
rect 537482 386280 537538 386336
rect 536930 378664 536986 378720
rect 538310 598168 538366 598224
rect 538310 388456 538366 388512
rect 539506 473184 539562 473240
rect 539966 637744 540022 637800
rect 539690 634616 539746 634672
rect 539782 624960 539838 625016
rect 539690 351056 539746 351112
rect 540242 637472 540298 637528
rect 540242 632168 540298 632224
rect 540150 628088 540206 628144
rect 540058 622376 540114 622432
rect 541070 657328 541126 657384
rect 543554 651208 543610 651264
rect 541162 645768 541218 645824
rect 541070 600480 541126 600536
rect 540426 476176 540482 476232
rect 540426 468424 540482 468480
rect 540242 385600 540298 385656
rect 540150 371864 540206 371920
rect 540058 362344 540114 362400
rect 541254 644408 541310 644464
rect 541346 641688 541402 641744
rect 542358 638968 542414 639024
rect 542726 637472 542782 637528
rect 542450 636248 542506 636304
rect 542542 633528 542598 633584
rect 542634 630808 542690 630864
rect 542726 629992 542782 630048
rect 542726 629448 542782 629504
rect 542634 385736 542690 385792
rect 542818 626728 542874 626784
rect 542910 617208 542966 617264
rect 542910 615848 542966 615904
rect 542910 389136 542966 389192
rect 542542 383016 542598 383072
rect 542450 382200 542506 382256
rect 542358 371320 542414 371376
rect 547878 699760 547934 699816
rect 545118 647128 545174 647184
rect 544382 629992 544438 630048
rect 544290 597896 544346 597952
rect 545118 601024 545174 601080
rect 544566 526496 544622 526552
rect 544566 476176 544622 476232
rect 544382 460128 544438 460184
rect 544290 388320 544346 388376
rect 546498 656920 546554 656976
rect 546682 657056 546738 657112
rect 546682 388728 546738 388784
rect 546498 386144 546554 386200
rect 529202 168952 529258 169008
rect 524326 166232 524382 166288
rect 500222 159704 500278 159760
rect 580262 697176 580318 697232
rect 548062 657192 548118 657248
rect 548062 388184 548118 388240
rect 580170 617516 580172 617536
rect 580172 617516 580224 617536
rect 580224 617516 580226 617536
rect 580170 617480 580226 617516
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 511264 580226 511320
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 378392 580226 378448
rect 580170 351872 580226 351928
rect 580354 644000 580410 644056
rect 580446 431568 580502 431624
rect 580262 325216 580318 325272
rect 580170 298696 580226 298752
rect 580262 272176 580318 272232
rect 580170 245520 580226 245576
rect 580170 205672 580226 205728
rect 580354 232328 580410 232384
rect 580446 219000 580502 219056
rect 580170 165824 580226 165880
rect 580538 192480 580594 192536
rect 580446 160656 580502 160712
rect 547878 158616 547934 158672
rect 580170 152632 580226 152688
rect 407210 139168 407266 139224
rect 407762 128016 407818 128072
rect 407210 116864 407266 116920
rect 407118 105712 407174 105768
rect 407210 100544 407266 100600
rect 382462 97824 382518 97880
rect 336278 85584 336334 85640
rect 332690 9016 332746 9072
rect 364614 85040 364670 85096
rect 357530 84904 357586 84960
rect 343362 84632 343418 84688
rect 339866 3304 339922 3360
rect 361118 84496 361174 84552
rect 368202 83408 368258 83464
rect 435362 83000 435418 83056
rect 432602 81640 432658 81696
rect 428554 80280 428610 80336
rect 421562 77560 421618 77616
rect 417422 76200 417478 76256
rect 414662 74840 414718 74896
rect 411902 57160 411958 57216
rect 389454 40704 389510 40760
rect 385958 15952 386014 16008
rect 378874 14592 378930 14648
rect 375286 11736 375342 11792
rect 382370 13096 382426 13152
rect 400126 39344 400182 39400
rect 396538 21392 396594 21448
rect 393042 18672 393098 18728
rect 407210 37984 407266 38040
rect 403622 17312 403678 17368
rect 410798 4800 410854 4856
rect 411902 4800 411958 4856
rect 414294 4800 414350 4856
rect 418802 61240 418858 61296
rect 417882 7656 417938 7712
rect 417422 3440 417478 3496
rect 414662 3032 414718 3088
rect 421378 53216 421434 53272
rect 418802 4800 418858 4856
rect 422942 68040 422998 68096
rect 425702 62600 425758 62656
rect 422942 7520 422998 7576
rect 424966 4800 425022 4856
rect 421562 3848 421618 3904
rect 425702 4120 425758 4176
rect 428462 4120 428518 4176
rect 431222 65320 431278 65376
rect 429842 63960 429898 64016
rect 431222 4936 431278 4992
rect 429842 4800 429898 4856
rect 432050 4800 432106 4856
rect 428554 3712 428610 3768
rect 450542 73480 450598 73536
rect 447782 72120 447838 72176
rect 443642 70760 443698 70816
rect 436742 66680 436798 66736
rect 435546 4936 435602 4992
rect 435362 3576 435418 3632
rect 432602 3168 432658 3224
rect 439502 47776 439558 47832
rect 436742 4120 436798 4176
rect 439134 4120 439190 4176
rect 442262 47640 442318 47696
rect 439502 3984 439558 4040
rect 442630 7520 442686 7576
rect 442262 3304 442318 3360
rect 446402 47504 446458 47560
rect 443642 4120 443698 4176
rect 446218 4120 446274 4176
rect 442906 3984 442962 4040
rect 467470 55800 467526 55856
rect 450542 4800 450598 4856
rect 453302 4800 453358 4856
rect 447782 4120 447838 4176
rect 449806 4120 449862 4176
rect 463974 3848 464030 3904
rect 460386 3440 460442 3496
rect 456890 3032 456946 3088
rect 517150 49000 517206 49056
rect 481730 46280 481786 46336
rect 471058 3712 471114 3768
rect 478142 3576 478198 3632
rect 474554 3168 474610 3224
rect 499394 43424 499450 43480
rect 495898 12960 495954 13016
rect 492310 11600 492366 11656
rect 488814 10240 488870 10296
rect 485226 8880 485282 8936
rect 506478 42064 506534 42120
rect 502982 14456 503038 14512
rect 512642 40568 512698 40624
rect 510066 15816 510122 15872
rect 512642 3440 512698 3496
rect 513562 3440 513618 3496
rect 580170 86128 580226 86184
rect 576122 48864 576178 48920
rect 549074 44784 549130 44840
rect 520738 39208 520794 39264
rect 524234 37848 524290 37904
rect 527822 36488 527878 36544
rect 534906 35128 534962 35184
rect 531318 17176 531374 17232
rect 538402 33768 538458 33824
rect 541990 30912 542046 30968
rect 545486 29552 545542 29608
rect 552662 28192 552718 28248
rect 559746 26832 559802 26888
rect 555422 18536 555478 18592
rect 562322 25472 562378 25528
rect 566830 24112 566886 24168
rect 562322 3440 562378 3496
rect 563242 3440 563298 3496
rect 570326 22616 570382 22672
rect 573914 21256 573970 21312
rect 580170 46280 580226 46336
rect 580170 6568 580226 6624
rect 576122 3984 576178 4040
rect 577410 3984 577466 4040
rect 582194 3304 582250 3360
<< metal3 >>
rect 163497 700498 163563 700501
rect 202781 700498 202847 700501
rect 163497 700496 202847 700498
rect 163497 700440 163502 700496
rect 163558 700440 202786 700496
rect 202842 700440 202847 700496
rect 163497 700438 202847 700440
rect 163497 700435 163563 700438
rect 202781 700435 202847 700438
rect 24301 700362 24367 700365
rect 31017 700362 31083 700365
rect 24301 700360 31083 700362
rect 24301 700304 24306 700360
rect 24362 700304 31022 700360
rect 31078 700304 31083 700360
rect 24301 700302 31083 700304
rect 24301 700299 24367 700302
rect 31017 700299 31083 700302
rect 43069 700362 43135 700365
rect 89161 700362 89227 700365
rect 43069 700360 89227 700362
rect 43069 700304 43074 700360
rect 43130 700304 89166 700360
rect 89222 700304 89227 700360
rect 43069 700302 89227 700304
rect 43069 700299 43135 700302
rect 89161 700299 89227 700302
rect 135897 700362 135963 700365
rect 154113 700362 154179 700365
rect 135897 700360 154179 700362
rect 135897 700304 135902 700360
rect 135958 700304 154118 700360
rect 154174 700304 154179 700360
rect 135897 700302 154179 700304
rect 135897 700299 135963 700302
rect 154113 700299 154179 700302
rect 176929 700362 176995 700365
rect 218973 700362 219039 700365
rect 176929 700360 219039 700362
rect 176929 700304 176934 700360
rect 176990 700304 218978 700360
rect 219034 700304 219039 700360
rect 176929 700302 219039 700304
rect 176929 700299 176995 700302
rect 218973 700299 219039 700302
rect 235165 700362 235231 700365
rect 323577 700362 323643 700365
rect 235165 700360 323643 700362
rect 235165 700304 235170 700360
rect 235226 700304 323582 700360
rect 323638 700304 323643 700360
rect 235165 700302 323643 700304
rect 235165 700299 235231 700302
rect 323577 700299 323643 700302
rect 543457 699818 543523 699821
rect 547873 699818 547939 699821
rect 543457 699816 547939 699818
rect 543457 699760 543462 699816
rect 543518 699760 547878 699816
rect 547934 699760 547939 699816
rect 543457 699758 547939 699760
rect 543457 699755 543523 699758
rect 547873 699755 547939 699758
rect 173157 698322 173223 698325
rect 176929 698322 176995 698325
rect 173157 698320 176995 698322
rect 173157 698264 173162 698320
rect 173218 698264 176934 698320
rect 176990 698264 176995 698320
rect 173157 698262 176995 698264
rect 173157 698259 173223 698262
rect 176929 698259 176995 698262
rect -960 697220 480 697460
rect 580257 697234 580323 697237
rect 583520 697234 584960 697324
rect 580257 697232 584960 697234
rect 580257 697176 580262 697232
rect 580318 697176 584960 697232
rect 580257 697174 584960 697176
rect 580257 697171 580323 697174
rect 583520 697084 584960 697174
rect 164417 688530 164483 688533
rect 173157 688530 173223 688533
rect 164417 688528 173223 688530
rect 164417 688472 164422 688528
rect 164478 688472 173162 688528
rect 173218 688472 173223 688528
rect 164417 688470 173223 688472
rect 164417 688467 164483 688470
rect 173157 688467 173223 688470
rect 160093 687170 160159 687173
rect 163497 687170 163563 687173
rect 160093 687168 163563 687170
rect 160093 687112 160098 687168
rect 160154 687112 163502 687168
rect 163558 687112 163563 687168
rect 160093 687110 163563 687112
rect 160093 687107 160159 687110
rect 163497 687107 163563 687110
rect 158713 685130 158779 685133
rect 160093 685130 160159 685133
rect 158713 685128 160159 685130
rect 158713 685072 158718 685128
rect 158774 685072 160098 685128
rect 160154 685072 160159 685128
rect 158713 685070 160159 685072
rect 158713 685067 158779 685070
rect 160093 685067 160159 685070
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 558126 683844 558132 683908
rect 558196 683906 558202 683908
rect 583520 683906 584960 683996
rect 558196 683846 584960 683906
rect 558196 683844 558202 683846
rect 583520 683756 584960 683846
rect 162117 677514 162183 677517
rect 163681 677514 163747 677517
rect 162117 677512 163747 677514
rect 162117 677456 162122 677512
rect 162178 677456 163686 677512
rect 163742 677456 163747 677512
rect 162117 677454 163747 677456
rect 162117 677451 162183 677454
rect 163681 677451 163747 677454
rect 153837 674794 153903 674797
rect 158621 674794 158687 674797
rect 153837 674792 158687 674794
rect 153837 674736 153842 674792
rect 153898 674736 158626 674792
rect 158682 674736 158687 674792
rect 153837 674734 158687 674736
rect 153837 674731 153903 674734
rect 158621 674731 158687 674734
rect -960 671258 480 671348
rect 30414 671258 30420 671260
rect -960 671198 30420 671258
rect -960 671108 480 671198
rect 30414 671196 30420 671198
rect 30484 671196 30490 671260
rect 507761 670714 507827 670717
rect 583520 670714 584960 670804
rect 507761 670712 584960 670714
rect 507761 670656 507766 670712
rect 507822 670656 584960 670712
rect 507761 670654 584960 670656
rect 507761 670651 507827 670654
rect 583520 670564 584960 670654
rect 158805 667858 158871 667861
rect 162117 667858 162183 667861
rect 158805 667856 162183 667858
rect 158805 667800 158810 667856
rect 158866 667800 162122 667856
rect 162178 667800 162183 667856
rect 158805 667798 162183 667800
rect 158805 667795 158871 667798
rect 162117 667795 162183 667798
rect 157333 665818 157399 665821
rect 158805 665818 158871 665821
rect 157333 665816 158871 665818
rect 157333 665760 157338 665816
rect 157394 665760 158810 665816
rect 158866 665760 158871 665816
rect 157333 665758 158871 665760
rect 157333 665755 157399 665758
rect 158805 665755 158871 665758
rect 151077 662554 151143 662557
rect 153837 662554 153903 662557
rect 151077 662552 153903 662554
rect 151077 662496 151082 662552
rect 151138 662496 153842 662552
rect 153898 662496 153903 662552
rect 151077 662494 153903 662496
rect 151077 662491 151143 662494
rect 153837 662491 153903 662494
rect -960 658202 480 658292
rect 15694 658202 15700 658204
rect -960 658142 15700 658202
rect -960 658052 480 658142
rect 15694 658140 15700 658142
rect 15764 658140 15770 658204
rect 489821 657930 489887 657933
rect 494697 657930 494763 657933
rect 489821 657928 494763 657930
rect 489821 657872 489826 657928
rect 489882 657872 494702 657928
rect 494758 657872 494763 657928
rect 489821 657870 494763 657872
rect 489821 657867 489887 657870
rect 494697 657867 494763 657870
rect 429837 657794 429903 657797
rect 491109 657794 491175 657797
rect 429837 657792 491175 657794
rect 429837 657736 429842 657792
rect 429898 657736 491114 657792
rect 491170 657736 491175 657792
rect 429837 657734 491175 657736
rect 429837 657731 429903 657734
rect 491109 657731 491175 657734
rect 151169 657658 151235 657661
rect 157333 657658 157399 657661
rect 151169 657656 157399 657658
rect 151169 657600 151174 657656
rect 151230 657600 157338 657656
rect 157394 657600 157399 657656
rect 151169 657598 157399 657600
rect 151169 657595 151235 657598
rect 157333 657595 157399 657598
rect 323577 657658 323643 657661
rect 515581 657658 515647 657661
rect 323577 657656 515647 657658
rect 323577 657600 323582 657656
rect 323638 657600 515586 657656
rect 515642 657600 515647 657656
rect 323577 657598 515647 657600
rect 323577 657595 323643 657598
rect 515581 657595 515647 657598
rect 87597 657522 87663 657525
rect 521101 657522 521167 657525
rect 87597 657520 521167 657522
rect 87597 657464 87602 657520
rect 87658 657464 521106 657520
rect 521162 657464 521167 657520
rect 87597 657462 521167 657464
rect 87597 657459 87663 657462
rect 521101 657459 521167 657462
rect 507761 657386 507827 657389
rect 541065 657386 541131 657389
rect 507761 657384 541131 657386
rect 507761 657328 507766 657384
rect 507822 657328 541070 657384
rect 541126 657328 541131 657384
rect 507761 657326 541131 657328
rect 507761 657323 507827 657326
rect 541065 657323 541131 657326
rect 537661 657250 537727 657253
rect 548057 657250 548123 657253
rect 537661 657248 548123 657250
rect 537661 657192 537666 657248
rect 537722 657192 548062 657248
rect 548118 657192 548123 657248
rect 583520 657236 584960 657476
rect 537661 657190 548123 657192
rect 537661 657187 537727 657190
rect 548057 657187 548123 657190
rect 515581 657114 515647 657117
rect 535453 657114 535519 657117
rect 515581 657112 535519 657114
rect 515581 657056 515586 657112
rect 515642 657056 535458 657112
rect 535514 657056 535519 657112
rect 515581 657054 535519 657056
rect 515581 657051 515647 657054
rect 535453 657051 535519 657054
rect 536281 657114 536347 657117
rect 546677 657114 546743 657117
rect 536281 657112 546743 657114
rect 536281 657056 536286 657112
rect 536342 657056 546682 657112
rect 546738 657056 546743 657112
rect 536281 657054 546743 657056
rect 536281 657051 536347 657054
rect 546677 657051 546743 657054
rect 539041 656978 539107 656981
rect 546493 656978 546559 656981
rect 539041 656976 546559 656978
rect 539041 656920 539046 656976
rect 539102 656920 546498 656976
rect 546554 656920 546559 656976
rect 539041 656918 546559 656920
rect 539041 656915 539107 656918
rect 546493 656915 546559 656918
rect 535453 655618 535519 655621
rect 535453 655616 538230 655618
rect 535453 655560 535458 655616
rect 535514 655560 538230 655616
rect 535453 655558 538230 655560
rect 535453 655555 535519 655558
rect 538170 655482 538230 655558
rect 540237 655482 540303 655485
rect 538170 655480 540303 655482
rect 538170 655424 540242 655480
rect 540298 655424 540303 655480
rect 538170 655422 540303 655424
rect 540237 655419 540303 655422
rect 27429 655074 27495 655077
rect 178033 655074 178099 655077
rect 27429 655072 178099 655074
rect 27429 655016 27434 655072
rect 27490 655016 178038 655072
rect 178094 655016 178099 655072
rect 27429 655014 178099 655016
rect 27429 655011 27495 655014
rect 178033 655011 178099 655014
rect 179270 655012 179276 655076
rect 179340 655074 179346 655076
rect 450486 655074 450492 655076
rect 179340 655014 450492 655074
rect 179340 655012 179346 655014
rect 450486 655012 450492 655014
rect 450556 655012 450562 655076
rect 177849 654938 177915 654941
rect 475377 654938 475443 654941
rect 177849 654936 475443 654938
rect 177849 654880 177854 654936
rect 177910 654880 475382 654936
rect 475438 654880 475443 654936
rect 177849 654878 475443 654880
rect 177849 654875 177915 654878
rect 475377 654875 475443 654878
rect 177665 654802 177731 654805
rect 482461 654802 482527 654805
rect 177665 654800 482527 654802
rect 177665 654744 177670 654800
rect 177726 654744 482466 654800
rect 482522 654744 482527 654800
rect 177665 654742 482527 654744
rect 177665 654739 177731 654742
rect 482461 654739 482527 654742
rect 33041 654666 33107 654669
rect 359365 654666 359431 654669
rect 33041 654664 359431 654666
rect 33041 654608 33046 654664
rect 33102 654608 359370 654664
rect 359426 654608 359431 654664
rect 33041 654606 359431 654608
rect 33041 654603 33107 654606
rect 359365 654603 359431 654606
rect 30189 654530 30255 654533
rect 356789 654530 356855 654533
rect 30189 654528 356855 654530
rect 30189 654472 30194 654528
rect 30250 654472 356794 654528
rect 356850 654472 356855 654528
rect 30189 654470 356855 654472
rect 30189 654467 30255 654470
rect 356789 654467 356855 654470
rect 488165 654530 488231 654533
rect 500401 654530 500467 654533
rect 488165 654528 500467 654530
rect 488165 654472 488170 654528
rect 488226 654472 500406 654528
rect 500462 654472 500467 654528
rect 488165 654470 500467 654472
rect 488165 654467 488231 654470
rect 500401 654467 500467 654470
rect 30281 654394 30347 654397
rect 358077 654394 358143 654397
rect 30281 654392 358143 654394
rect 30281 654336 30286 654392
rect 30342 654336 358082 654392
rect 358138 654336 358143 654392
rect 30281 654334 358143 654336
rect 30281 654331 30347 654334
rect 358077 654331 358143 654334
rect 26785 654258 26851 654261
rect 363229 654258 363295 654261
rect 26785 654256 363295 654258
rect 26785 654200 26790 654256
rect 26846 654200 363234 654256
rect 363290 654200 363295 654256
rect 26785 654198 363295 654200
rect 26785 654195 26851 654198
rect 363229 654195 363295 654198
rect 41321 653714 41387 653717
rect 305269 653714 305335 653717
rect 41321 653712 305335 653714
rect 41321 653656 41326 653712
rect 41382 653656 305274 653712
rect 305330 653656 305335 653712
rect 41321 653654 305335 653656
rect 41321 653651 41387 653654
rect 305269 653651 305335 653654
rect 189165 653578 189231 653581
rect 463141 653578 463207 653581
rect 189165 653576 463207 653578
rect 189165 653520 189170 653576
rect 189226 653520 463146 653576
rect 463202 653520 463207 653576
rect 189165 653518 463207 653520
rect 189165 653515 189231 653518
rect 463141 653515 463207 653518
rect 190453 653442 190519 653445
rect 465717 653442 465783 653445
rect 190453 653440 465783 653442
rect 190453 653384 190458 653440
rect 190514 653384 465722 653440
rect 465778 653384 465783 653440
rect 190453 653382 465783 653384
rect 190453 653379 190519 653382
rect 465717 653379 465783 653382
rect 194317 653306 194383 653309
rect 471329 653306 471395 653309
rect 194317 653304 471395 653306
rect 194317 653248 194322 653304
rect 194378 653248 471334 653304
rect 471390 653248 471395 653304
rect 194317 653246 471395 653248
rect 194317 653243 194383 653246
rect 471329 653243 471395 653246
rect 175038 653108 175044 653172
rect 175108 653170 175114 653172
rect 480294 653170 480300 653172
rect 175108 653110 480300 653170
rect 175108 653108 175114 653110
rect 480294 653108 480300 653110
rect 480364 653108 480370 653172
rect 33777 653034 33843 653037
rect 360653 653034 360719 653037
rect 33777 653032 360719 653034
rect 33777 652976 33782 653032
rect 33838 652976 360658 653032
rect 360714 652976 360719 653032
rect 33777 652974 360719 652976
rect 33777 652971 33843 652974
rect 360653 652971 360719 652974
rect 28257 652898 28323 652901
rect 364517 652898 364583 652901
rect 28257 652896 364583 652898
rect 28257 652840 28262 652896
rect 28318 652840 364522 652896
rect 364578 652840 364583 652896
rect 28257 652838 364583 652840
rect 28257 652835 28323 652838
rect 364517 652835 364583 652838
rect 184013 652354 184079 652357
rect 227713 652354 227779 652357
rect 184013 652352 227779 652354
rect 184013 652296 184018 652352
rect 184074 652296 227718 652352
rect 227774 652296 227779 652352
rect 184013 652294 227779 652296
rect 184013 652291 184079 652294
rect 227713 652291 227779 652294
rect 227805 652218 227871 652221
rect 461577 652218 461643 652221
rect 227805 652216 461643 652218
rect 227805 652160 227810 652216
rect 227866 652160 461582 652216
rect 461638 652160 461643 652216
rect 227805 652158 461643 652160
rect 227805 652155 227871 652158
rect 461577 652155 461643 652158
rect 185301 652082 185367 652085
rect 233141 652082 233207 652085
rect 185301 652080 233207 652082
rect 185301 652024 185306 652080
rect 185362 652024 233146 652080
rect 233202 652024 233207 652080
rect 185301 652022 233207 652024
rect 185301 652019 185367 652022
rect 233141 652019 233207 652022
rect 233417 652082 233483 652085
rect 479609 652082 479675 652085
rect 233417 652080 479675 652082
rect 233417 652024 233422 652080
rect 233478 652024 479614 652080
rect 479670 652024 479675 652080
rect 233417 652022 479675 652024
rect 233417 652019 233483 652022
rect 479609 652019 479675 652022
rect 211061 651946 211127 651949
rect 469857 651946 469923 651949
rect 211061 651944 469923 651946
rect 211061 651888 211066 651944
rect 211122 651888 469862 651944
rect 469918 651888 469923 651944
rect 211061 651886 469923 651888
rect 211061 651883 211127 651886
rect 469857 651883 469923 651886
rect 208485 651810 208551 651813
rect 468477 651810 468543 651813
rect 208485 651808 468543 651810
rect 208485 651752 208490 651808
rect 208546 651752 468482 651808
rect 468538 651752 468543 651808
rect 208485 651750 468543 651752
rect 208485 651747 208551 651750
rect 468477 651747 468543 651750
rect 31661 651674 31727 651677
rect 213821 651674 213887 651677
rect 31661 651672 213887 651674
rect 31661 651616 31666 651672
rect 31722 651616 213826 651672
rect 213882 651616 213887 651672
rect 31661 651614 213887 651616
rect 31661 651611 31727 651614
rect 213821 651611 213887 651614
rect 214097 651674 214163 651677
rect 487981 651674 488047 651677
rect 214097 651672 488047 651674
rect 214097 651616 214102 651672
rect 214158 651616 487986 651672
rect 488042 651616 488047 651672
rect 214097 651614 488047 651616
rect 214097 651611 214163 651614
rect 487981 651611 488047 651614
rect 207197 651538 207263 651541
rect 487797 651538 487863 651541
rect 207197 651536 487863 651538
rect 207197 651480 207202 651536
rect 207258 651480 487802 651536
rect 487858 651480 487863 651536
rect 207197 651478 487863 651480
rect 207197 651475 207263 651478
rect 487797 651475 487863 651478
rect 187877 651402 187943 651405
rect 478229 651402 478295 651405
rect 187877 651400 478295 651402
rect 187877 651344 187882 651400
rect 187938 651344 478234 651400
rect 478290 651344 478295 651400
rect 187877 651342 478295 651344
rect 187877 651339 187943 651342
rect 478229 651339 478295 651342
rect 543549 651266 543615 651269
rect 539948 651264 543615 651266
rect 539948 651208 543554 651264
rect 543610 651208 543615 651264
rect 539948 651206 543615 651208
rect 543549 651203 543615 651206
rect 39665 651130 39731 651133
rect 226333 651130 226399 651133
rect 39665 651128 226399 651130
rect 39665 651072 39670 651128
rect 39726 651072 226338 651128
rect 226394 651072 226399 651128
rect 39665 651070 226399 651072
rect 39665 651067 39731 651070
rect 226333 651067 226399 651070
rect 39757 650994 39823 650997
rect 214557 650994 214623 650997
rect 39757 650992 214623 650994
rect 39757 650936 39762 650992
rect 39818 650936 214562 650992
rect 214618 650936 214623 650992
rect 39757 650934 214623 650936
rect 39757 650931 39823 650934
rect 214557 650931 214623 650934
rect 226517 650858 226583 650861
rect 461761 650858 461827 650861
rect 226517 650856 461827 650858
rect 226517 650800 226522 650856
rect 226578 650800 461766 650856
rect 461822 650800 461827 650856
rect 226517 650798 461827 650800
rect 226517 650795 226583 650798
rect 461761 650795 461827 650798
rect 39849 650722 39915 650725
rect 212441 650722 212507 650725
rect 39849 650720 212507 650722
rect 39849 650664 39854 650720
rect 39910 650664 212446 650720
rect 212502 650664 212507 650720
rect 39849 650662 212507 650664
rect 39849 650659 39915 650662
rect 212441 650659 212507 650662
rect 214925 650722 214991 650725
rect 467373 650722 467439 650725
rect 214925 650720 467439 650722
rect 214925 650664 214930 650720
rect 214986 650664 467378 650720
rect 467434 650664 467439 650720
rect 214925 650662 467439 650664
rect 214925 650659 214991 650662
rect 467373 650659 467439 650662
rect 42149 650586 42215 650589
rect 231761 650586 231827 650589
rect 42149 650584 231827 650586
rect 42149 650528 42154 650584
rect 42210 650528 231766 650584
rect 231822 650528 231827 650584
rect 42149 650526 231827 650528
rect 42149 650523 42215 650526
rect 231761 650523 231827 650526
rect 232037 650586 232103 650589
rect 485037 650586 485103 650589
rect 232037 650584 485103 650586
rect 232037 650528 232042 650584
rect 232098 650528 485042 650584
rect 485098 650528 485103 650584
rect 232037 650526 485103 650528
rect 232037 650523 232103 650526
rect 485037 650523 485103 650526
rect 40769 650450 40835 650453
rect 186313 650450 186379 650453
rect 40769 650448 186379 650450
rect 40769 650392 40774 650448
rect 40830 650392 186318 650448
rect 186374 650392 186379 650448
rect 40769 650390 186379 650392
rect 40769 650387 40835 650390
rect 186313 650387 186379 650390
rect 212349 650450 212415 650453
rect 467189 650450 467255 650453
rect 212349 650448 467255 650450
rect 212349 650392 212354 650448
rect 212410 650392 467194 650448
rect 467250 650392 467255 650448
rect 212349 650390 467255 650392
rect 212349 650387 212415 650390
rect 467189 650387 467255 650390
rect 42701 650314 42767 650317
rect 324589 650314 324655 650317
rect 42701 650312 324655 650314
rect 42701 650256 42706 650312
rect 42762 650256 324594 650312
rect 324650 650256 324655 650312
rect 42701 650254 324655 650256
rect 42701 650251 42767 650254
rect 324589 650251 324655 650254
rect 186589 650178 186655 650181
rect 480989 650178 481055 650181
rect 186589 650176 481055 650178
rect 186589 650120 186594 650176
rect 186650 650120 480994 650176
rect 481050 650120 481055 650176
rect 186589 650118 481055 650120
rect 186589 650115 186655 650118
rect 480989 650115 481055 650118
rect 176510 649980 176516 650044
rect 176580 650042 176586 650044
rect 476614 650042 476620 650044
rect 176580 649982 476620 650042
rect 176580 649980 176586 649982
rect 476614 649980 476620 649982
rect 476684 649980 476690 650044
rect 550766 649906 550772 649908
rect 539948 649846 550772 649906
rect 550766 649844 550772 649846
rect 550836 649844 550842 649908
rect 205909 649770 205975 649773
rect 224217 649770 224283 649773
rect 205909 649768 224283 649770
rect 205909 649712 205914 649768
rect 205970 649712 224222 649768
rect 224278 649712 224283 649768
rect 205909 649710 224283 649712
rect 205909 649707 205975 649710
rect 224217 649707 224283 649710
rect 53557 649634 53623 649637
rect 345197 649634 345263 649637
rect 53557 649632 345263 649634
rect 53557 649576 53562 649632
rect 53618 649576 345202 649632
rect 345258 649576 345263 649632
rect 53557 649574 345263 649576
rect 53557 649571 53623 649574
rect 345197 649571 345263 649574
rect 149697 649498 149763 649501
rect 151169 649498 151235 649501
rect 149697 649496 151235 649498
rect 149697 649440 149702 649496
rect 149758 649440 151174 649496
rect 151230 649440 151235 649496
rect 149697 649438 151235 649440
rect 149697 649435 149763 649438
rect 151169 649435 151235 649438
rect 223941 649498 224007 649501
rect 467281 649498 467347 649501
rect 223941 649496 467347 649498
rect 223941 649440 223946 649496
rect 224002 649440 467286 649496
rect 467342 649440 467347 649496
rect 223941 649438 467347 649440
rect 223941 649435 224007 649438
rect 467281 649435 467347 649438
rect 51441 649362 51507 649365
rect 314285 649362 314351 649365
rect 51441 649360 314351 649362
rect 51441 649304 51446 649360
rect 51502 649304 314290 649360
rect 314346 649304 314351 649360
rect 51441 649302 314351 649304
rect 51441 649299 51507 649302
rect 314285 649299 314351 649302
rect 52269 649226 52335 649229
rect 334893 649226 334959 649229
rect 52269 649224 334959 649226
rect 52269 649168 52274 649224
rect 52330 649168 334898 649224
rect 334954 649168 334959 649224
rect 52269 649166 334959 649168
rect 52269 649163 52335 649166
rect 334893 649163 334959 649166
rect 54845 649090 54911 649093
rect 343909 649090 343975 649093
rect 54845 649088 343975 649090
rect 54845 649032 54850 649088
rect 54906 649032 343914 649088
rect 343970 649032 343975 649088
rect 54845 649030 343975 649032
rect 54845 649027 54911 649030
rect 343909 649027 343975 649030
rect 41229 648954 41295 648957
rect 332317 648954 332383 648957
rect 41229 648952 332383 648954
rect 41229 648896 41234 648952
rect 41290 648896 332322 648952
rect 332378 648896 332383 648952
rect 41229 648894 332383 648896
rect 41229 648891 41295 648894
rect 332317 648891 332383 648894
rect 56225 648818 56291 648821
rect 347773 648818 347839 648821
rect 56225 648816 347839 648818
rect 56225 648760 56230 648816
rect 56286 648760 347778 648816
rect 347834 648760 347839 648816
rect 56225 648758 347839 648760
rect 56225 648755 56291 648758
rect 347773 648755 347839 648758
rect 196893 648682 196959 648685
rect 198733 648682 198799 648685
rect 196893 648680 198799 648682
rect 196893 648624 196898 648680
rect 196954 648624 198738 648680
rect 198794 648624 198799 648680
rect 196893 648622 198799 648624
rect 196893 648619 196959 648622
rect 198733 648619 198799 648622
rect 200757 648682 200823 648685
rect 205633 648682 205699 648685
rect 200757 648680 205699 648682
rect 200757 648624 200762 648680
rect 200818 648624 205638 648680
rect 205694 648624 205699 648680
rect 200757 648622 205699 648624
rect 200757 648619 200823 648622
rect 205633 648619 205699 648622
rect 44030 648212 44036 648276
rect 44100 648274 44106 648276
rect 377622 648274 377628 648276
rect 44100 648214 377628 648274
rect 44100 648212 44106 648214
rect 377622 648212 377628 648214
rect 377692 648212 377698 648276
rect 51809 648138 51875 648141
rect 234613 648138 234679 648141
rect 51809 648136 234679 648138
rect 51809 648080 51814 648136
rect 51870 648080 234618 648136
rect 234674 648080 234679 648136
rect 51809 648078 234679 648080
rect 51809 648075 51875 648078
rect 234613 648075 234679 648078
rect 235533 648138 235599 648141
rect 461669 648138 461735 648141
rect 235533 648136 461735 648138
rect 235533 648080 235538 648136
rect 235594 648080 461674 648136
rect 461730 648080 461735 648136
rect 235533 648078 461735 648080
rect 235533 648075 235599 648078
rect 461669 648075 461735 648078
rect 54109 648002 54175 648005
rect 327165 648002 327231 648005
rect 54109 648000 327231 648002
rect 54109 647944 54114 648000
rect 54170 647944 327170 648000
rect 327226 647944 327231 648000
rect 54109 647942 327231 647944
rect 54109 647939 54175 647942
rect 327165 647939 327231 647942
rect 56409 647866 56475 647869
rect 333605 647866 333671 647869
rect 56409 647864 333671 647866
rect 56409 647808 56414 647864
rect 56470 647808 333610 647864
rect 333666 647808 333671 647864
rect 56409 647806 333671 647808
rect 539918 647866 539978 648516
rect 539918 647806 547706 647866
rect 56409 647803 56475 647806
rect 333605 647803 333671 647806
rect 52177 647730 52243 647733
rect 336181 647730 336247 647733
rect 52177 647728 336247 647730
rect 52177 647672 52182 647728
rect 52238 647672 336186 647728
rect 336242 647672 336247 647728
rect 52177 647670 336247 647672
rect 52177 647667 52243 647670
rect 336181 647667 336247 647670
rect 43989 647594 44055 647597
rect 329741 647594 329807 647597
rect 43989 647592 329807 647594
rect 43989 647536 43994 647592
rect 44050 647536 329746 647592
rect 329802 647536 329807 647592
rect 43989 647534 329807 647536
rect 43989 647531 44055 647534
rect 329741 647531 329807 647534
rect 52085 647458 52151 647461
rect 341333 647458 341399 647461
rect 52085 647456 341399 647458
rect 52085 647400 52090 647456
rect 52146 647400 341338 647456
rect 341394 647400 341399 647456
rect 52085 647398 341399 647400
rect 52085 647395 52151 647398
rect 341333 647395 341399 647398
rect 176326 647260 176332 647324
rect 176396 647322 176402 647324
rect 176561 647322 176627 647325
rect 547646 647324 547706 647806
rect 176396 647320 176627 647322
rect 176396 647264 176566 647320
rect 176622 647264 176627 647320
rect 176396 647262 176627 647264
rect 176396 647260 176402 647262
rect 176561 647259 176627 647262
rect 547638 647260 547644 647324
rect 547708 647260 547714 647324
rect 545113 647186 545179 647189
rect 539948 647184 545179 647186
rect 539948 647128 545118 647184
rect 545174 647128 545179 647184
rect 539948 647126 545179 647128
rect 545113 647123 545179 647126
rect 66529 646914 66595 646917
rect 387149 646914 387215 646917
rect 66529 646912 387215 646914
rect 66529 646856 66534 646912
rect 66590 646856 387154 646912
rect 387210 646856 387215 646912
rect 66529 646854 387215 646856
rect 66529 646851 66595 646854
rect 387149 646851 387215 646854
rect 53005 646778 53071 646781
rect 115841 646778 115907 646781
rect 425605 646778 425671 646781
rect 53005 646776 115907 646778
rect 53005 646720 53010 646776
rect 53066 646720 115846 646776
rect 115902 646720 115907 646776
rect 53005 646718 115907 646720
rect 53005 646715 53071 646718
rect 115841 646715 115907 646718
rect 115982 646776 425671 646778
rect 115982 646720 425610 646776
rect 425666 646720 425671 646776
rect 115982 646718 425671 646720
rect 115473 646642 115539 646645
rect 115982 646642 116042 646718
rect 425605 646715 425671 646718
rect 115473 646640 116042 646642
rect 115473 646584 115478 646640
rect 115534 646584 116042 646640
rect 115473 646582 116042 646584
rect 116117 646642 116183 646645
rect 424593 646642 424659 646645
rect 116117 646640 424659 646642
rect 116117 646584 116122 646640
rect 116178 646584 424598 646640
rect 424654 646584 424659 646640
rect 116117 646582 424659 646584
rect 115473 646579 115539 646582
rect 116117 646579 116183 646582
rect 424593 646579 424659 646582
rect 112897 646506 112963 646509
rect 423581 646506 423647 646509
rect 112897 646504 423647 646506
rect 112897 646448 112902 646504
rect 112958 646448 423586 646504
rect 423642 646448 423647 646504
rect 112897 646446 423647 646448
rect 112897 646443 112963 646446
rect 423581 646443 423647 646446
rect 73061 646370 73127 646373
rect 392209 646370 392275 646373
rect 73061 646368 392275 646370
rect 73061 646312 73066 646368
rect 73122 646312 392214 646368
rect 392270 646312 392275 646368
rect 73061 646310 392275 646312
rect 73061 646307 73127 646310
rect 392209 646307 392275 646310
rect 71681 646234 71747 646237
rect 391197 646234 391263 646237
rect 71681 646232 391263 646234
rect 71681 646176 71686 646232
rect 71742 646176 391202 646232
rect 391258 646176 391263 646232
rect 71681 646174 391263 646176
rect 71681 646171 71747 646174
rect 391197 646171 391263 646174
rect 67817 646098 67883 646101
rect 388161 646098 388227 646101
rect 67817 646096 388227 646098
rect 67817 646040 67822 646096
rect 67878 646040 388166 646096
rect 388222 646040 388227 646096
rect 67817 646038 388227 646040
rect 67817 646035 67883 646038
rect 388161 646035 388227 646038
rect 114185 645962 114251 645965
rect 116117 645962 116183 645965
rect 114185 645960 116183 645962
rect 114185 645904 114190 645960
rect 114246 645904 116122 645960
rect 116178 645904 116183 645960
rect 114185 645902 116183 645904
rect 114185 645899 114251 645902
rect 116117 645899 116183 645902
rect 176142 645900 176148 645964
rect 176212 645962 176218 645964
rect 176561 645962 176627 645965
rect 176212 645960 176627 645962
rect 176212 645904 176566 645960
rect 176622 645904 176627 645960
rect 176212 645902 176627 645904
rect 176212 645900 176218 645902
rect 176561 645899 176627 645902
rect 541157 645826 541223 645829
rect 539948 645824 541223 645826
rect 539948 645768 541162 645824
rect 541218 645768 541223 645824
rect 539948 645766 541223 645768
rect 541157 645763 541223 645766
rect 54886 645356 54892 645420
rect 54956 645418 54962 645420
rect 296846 645418 296852 645420
rect 54956 645358 296852 645418
rect 54956 645356 54962 645358
rect 296846 645356 296852 645358
rect 296916 645356 296922 645420
rect 62665 645282 62731 645285
rect 131113 645282 131179 645285
rect 62665 645280 131179 645282
rect -960 644996 480 645236
rect 62665 645224 62670 645280
rect 62726 645224 131118 645280
rect 131174 645224 131179 645280
rect 62665 645222 131179 645224
rect 62665 645219 62731 645222
rect 131113 645219 131179 645222
rect 132217 645282 132283 645285
rect 383101 645282 383167 645285
rect 132217 645280 383167 645282
rect 132217 645224 132222 645280
rect 132278 645224 383106 645280
rect 383162 645224 383167 645280
rect 132217 645222 383167 645224
rect 132217 645219 132283 645222
rect 383101 645219 383167 645222
rect 25681 645146 25747 645149
rect 91093 645146 91159 645149
rect 25681 645144 91159 645146
rect 25681 645088 25686 645144
rect 25742 645088 91098 645144
rect 91154 645088 91159 645144
rect 25681 645086 91159 645088
rect 25681 645083 25747 645086
rect 91093 645083 91159 645086
rect 92289 645146 92355 645149
rect 407389 645146 407455 645149
rect 92289 645144 407455 645146
rect 92289 645088 92294 645144
rect 92350 645088 407394 645144
rect 407450 645088 407455 645144
rect 92289 645086 407455 645088
rect 92289 645083 92355 645086
rect 407389 645083 407455 645086
rect 84561 645010 84627 645013
rect 401317 645010 401383 645013
rect 84561 645008 401383 645010
rect 84561 644952 84566 645008
rect 84622 644952 401322 645008
rect 401378 644952 401383 645008
rect 84561 644950 401383 644952
rect 84561 644947 84627 644950
rect 401317 644947 401383 644950
rect 80697 644874 80763 644877
rect 398281 644874 398347 644877
rect 80697 644872 398347 644874
rect 80697 644816 80702 644872
rect 80758 644816 398286 644872
rect 398342 644816 398347 644872
rect 80697 644814 398347 644816
rect 80697 644811 80763 644814
rect 398281 644811 398347 644814
rect 76833 644738 76899 644741
rect 395245 644738 395311 644741
rect 76833 644736 395311 644738
rect 76833 644680 76838 644736
rect 76894 644680 395250 644736
rect 395306 644680 395311 644736
rect 76833 644678 395311 644680
rect 76833 644675 76899 644678
rect 395245 644675 395311 644678
rect 75545 644602 75611 644605
rect 394233 644602 394299 644605
rect 75545 644600 394299 644602
rect 75545 644544 75550 644600
rect 75606 644544 394238 644600
rect 394294 644544 394299 644600
rect 75545 644542 394299 644544
rect 75545 644539 75611 644542
rect 394233 644539 394299 644542
rect 541249 644466 541315 644469
rect 539948 644464 541315 644466
rect 539948 644408 541254 644464
rect 541310 644408 541315 644464
rect 539948 644406 541315 644408
rect 541249 644403 541315 644406
rect 25865 644194 25931 644197
rect 126881 644194 126947 644197
rect 25865 644192 126947 644194
rect 25865 644136 25870 644192
rect 25926 644136 126886 644192
rect 126942 644136 126947 644192
rect 25865 644134 126947 644136
rect 25865 644131 25931 644134
rect 126881 644131 126947 644134
rect 46841 644058 46907 644061
rect 124121 644058 124187 644061
rect 46841 644056 124187 644058
rect 46841 644000 46846 644056
rect 46902 644000 124126 644056
rect 124182 644000 124187 644056
rect 46841 643998 124187 644000
rect 46841 643995 46907 643998
rect 124121 643995 124187 643998
rect 125777 644058 125843 644061
rect 261661 644058 261727 644061
rect 125777 644056 261727 644058
rect 125777 644000 125782 644056
rect 125838 644000 261666 644056
rect 261722 644000 261727 644056
rect 125777 643998 261727 644000
rect 125777 643995 125843 643998
rect 261661 643995 261727 643998
rect 580349 644058 580415 644061
rect 583520 644058 584960 644148
rect 580349 644056 584960 644058
rect 580349 644000 580354 644056
rect 580410 644000 584960 644056
rect 580349 643998 584960 644000
rect 580349 643995 580415 643998
rect 123201 643922 123267 643925
rect 259637 643922 259703 643925
rect 123201 643920 259703 643922
rect 123201 643864 123206 643920
rect 123262 643864 259642 643920
rect 259698 643864 259703 643920
rect 583520 643908 584960 643998
rect 123201 643862 259703 643864
rect 123201 643859 123267 643862
rect 259637 643859 259703 643862
rect 49601 643786 49667 643789
rect 297265 643786 297331 643789
rect 49601 643784 297331 643786
rect 49601 643728 49606 643784
rect 49662 643728 297270 643784
rect 297326 643728 297331 643784
rect 49601 643726 297331 643728
rect 49601 643723 49667 643726
rect 297265 643723 297331 643726
rect 48630 643588 48636 643652
rect 48700 643650 48706 643652
rect 297030 643650 297036 643652
rect 48700 643590 297036 643650
rect 48700 643588 48706 643590
rect 297030 643588 297036 643590
rect 297100 643588 297106 643652
rect 48037 643514 48103 643517
rect 297909 643514 297975 643517
rect 48037 643512 297975 643514
rect 48037 643456 48042 643512
rect 48098 643456 297914 643512
rect 297970 643456 297975 643512
rect 48037 643454 297975 643456
rect 48037 643451 48103 643454
rect 297909 643451 297975 643454
rect 46790 643316 46796 643380
rect 46860 643378 46866 643380
rect 297725 643378 297791 643381
rect 46860 643376 297791 643378
rect 46860 643320 297730 643376
rect 297786 643320 297791 643376
rect 46860 643318 297791 643320
rect 46860 643316 46866 643318
rect 297725 643315 297791 643318
rect 26049 643242 26115 643245
rect 328453 643242 328519 643245
rect 26049 643240 328519 643242
rect 26049 643184 26054 643240
rect 26110 643184 328458 643240
rect 328514 643184 328519 643240
rect 26049 643182 328519 643184
rect 26049 643179 26115 643182
rect 328453 643179 328519 643182
rect 550030 643106 550036 643108
rect 539948 643046 550036 643106
rect 550030 643044 550036 643046
rect 550100 643044 550106 643108
rect 51901 642970 51967 642973
rect 294045 642970 294111 642973
rect 51901 642968 294111 642970
rect 51901 642912 51906 642968
rect 51962 642912 294050 642968
rect 294106 642912 294111 642968
rect 51901 642910 294111 642912
rect 51901 642907 51967 642910
rect 294045 642907 294111 642910
rect 57881 642834 57947 642837
rect 380065 642834 380131 642837
rect 57881 642832 380131 642834
rect 57881 642776 57886 642832
rect 57942 642776 380070 642832
rect 380126 642776 380131 642832
rect 57881 642774 380131 642776
rect 57881 642771 57947 642774
rect 380065 642771 380131 642774
rect 48221 642698 48287 642701
rect 297541 642698 297607 642701
rect 48221 642696 297607 642698
rect 48221 642640 48226 642696
rect 48282 642640 297546 642696
rect 297602 642640 297607 642696
rect 48221 642638 297607 642640
rect 48221 642635 48287 642638
rect 297541 642635 297607 642638
rect 178677 642562 178743 642565
rect 298093 642562 298159 642565
rect 178677 642560 298159 642562
rect 178677 642504 178682 642560
rect 178738 642504 298098 642560
rect 298154 642504 298159 642560
rect 178677 642502 298159 642504
rect 178677 642499 178743 642502
rect 298093 642499 298159 642502
rect 31293 642426 31359 642429
rect 59261 642426 59327 642429
rect 293953 642426 294019 642429
rect 31293 642424 59327 642426
rect 31293 642368 31298 642424
rect 31354 642368 59266 642424
rect 59322 642368 59327 642424
rect 31293 642366 59327 642368
rect 31293 642363 31359 642366
rect 59261 642363 59327 642366
rect 64830 642424 294019 642426
rect 64830 642368 293958 642424
rect 294014 642368 294019 642424
rect 64830 642366 294019 642368
rect 59077 642290 59143 642293
rect 64830 642290 64890 642366
rect 293953 642363 294019 642366
rect 59077 642288 64890 642290
rect 59077 642232 59082 642288
rect 59138 642232 64890 642288
rect 59077 642230 64890 642232
rect 294781 642290 294847 642293
rect 475561 642290 475627 642293
rect 294781 642288 475627 642290
rect 294781 642232 294786 642288
rect 294842 642232 475566 642288
rect 475622 642232 475627 642288
rect 294781 642230 475627 642232
rect 59077 642227 59143 642230
rect 294781 642227 294847 642230
rect 475561 642227 475627 642230
rect 42517 642154 42583 642157
rect 178033 642154 178099 642157
rect 42517 642152 178099 642154
rect 42517 642096 42522 642152
rect 42578 642096 178038 642152
rect 178094 642096 178099 642152
rect 42517 642094 178099 642096
rect 42517 642091 42583 642094
rect 178033 642091 178099 642094
rect 294597 642154 294663 642157
rect 475745 642154 475811 642157
rect 294597 642152 475811 642154
rect 294597 642096 294602 642152
rect 294658 642096 475750 642152
rect 475806 642096 475811 642152
rect 294597 642094 475811 642096
rect 294597 642091 294663 642094
rect 475745 642091 475811 642094
rect 32857 642018 32923 642021
rect 323301 642018 323367 642021
rect 32857 642016 323367 642018
rect 32857 641960 32862 642016
rect 32918 641960 323306 642016
rect 323362 641960 323367 642016
rect 32857 641958 323367 641960
rect 32857 641955 32923 641958
rect 323301 641955 323367 641958
rect 50613 641882 50679 641885
rect 57881 641882 57947 641885
rect 50613 641880 57947 641882
rect 50613 641824 50618 641880
rect 50674 641824 57886 641880
rect 57942 641824 57947 641880
rect 50613 641822 57947 641824
rect 50613 641819 50679 641822
rect 57881 641819 57947 641822
rect 59169 641882 59235 641885
rect 381077 641882 381143 641885
rect 59169 641880 381143 641882
rect 59169 641824 59174 641880
rect 59230 641824 381082 641880
rect 381138 641824 381143 641880
rect 59169 641822 381143 641824
rect 59169 641819 59235 641822
rect 381077 641819 381143 641822
rect 54753 641746 54819 641749
rect 59261 641746 59327 641749
rect 54753 641744 59327 641746
rect 54753 641688 54758 641744
rect 54814 641688 59266 641744
rect 59322 641688 59327 641744
rect 54753 641686 59327 641688
rect 54753 641683 54819 641686
rect 59261 641683 59327 641686
rect 177062 641684 177068 641748
rect 177132 641746 177138 641748
rect 177941 641746 178007 641749
rect 541341 641746 541407 641749
rect 177132 641744 178007 641746
rect 177132 641688 177946 641744
rect 178002 641688 178007 641744
rect 177132 641686 178007 641688
rect 539948 641744 541407 641746
rect 539948 641688 541346 641744
rect 541402 641688 541407 641744
rect 539948 641686 541407 641688
rect 177132 641684 177138 641686
rect 177941 641683 178007 641686
rect 541341 641683 541407 641686
rect 51993 641474 52059 641477
rect 127617 641474 127683 641477
rect 51993 641472 127683 641474
rect 51993 641416 51998 641472
rect 52054 641416 127622 641472
rect 127678 641416 127683 641472
rect 51993 641414 127683 641416
rect 51993 641411 52059 641414
rect 127617 641411 127683 641414
rect 30005 641338 30071 641341
rect 251081 641338 251147 641341
rect 30005 641336 251147 641338
rect 30005 641280 30010 641336
rect 30066 641280 251086 641336
rect 251142 641280 251147 641336
rect 30005 641278 251147 641280
rect 30005 641275 30071 641278
rect 251081 641275 251147 641278
rect 127065 641202 127131 641205
rect 262673 641202 262739 641205
rect 127065 641200 262739 641202
rect 127065 641144 127070 641200
rect 127126 641144 262678 641200
rect 262734 641144 262739 641200
rect 127065 641142 262739 641144
rect 127065 641139 127131 641142
rect 262673 641139 262739 641142
rect 294822 641140 294828 641204
rect 294892 641202 294898 641204
rect 479374 641202 479380 641204
rect 294892 641142 479380 641202
rect 294892 641140 294898 641142
rect 479374 641140 479380 641142
rect 479444 641140 479450 641204
rect 488073 641202 488139 641205
rect 488073 641200 490084 641202
rect 488073 641144 488078 641200
rect 488134 641144 490084 641200
rect 488073 641142 490084 641144
rect 488073 641139 488139 641142
rect 56317 641066 56383 641069
rect 249701 641066 249767 641069
rect 56317 641064 249767 641066
rect 56317 641008 56322 641064
rect 56378 641008 249706 641064
rect 249762 641008 249767 641064
rect 56317 641006 249767 641008
rect 56317 641003 56383 641006
rect 249701 641003 249767 641006
rect 259361 641066 259427 641069
rect 370957 641066 371023 641069
rect 259361 641064 371023 641066
rect 259361 641008 259366 641064
rect 259422 641008 370962 641064
rect 371018 641008 371023 641064
rect 259361 641006 371023 641008
rect 259361 641003 259427 641006
rect 370957 641003 371023 641006
rect 48129 640930 48195 640933
rect 297633 640930 297699 640933
rect 48129 640928 297699 640930
rect 48129 640872 48134 640928
rect 48190 640872 297638 640928
rect 297694 640872 297699 640928
rect 48129 640870 297699 640872
rect 48129 640867 48195 640870
rect 297633 640867 297699 640870
rect 55581 640794 55647 640797
rect 316861 640794 316927 640797
rect 55581 640792 316927 640794
rect 55581 640736 55586 640792
rect 55642 640736 316866 640792
rect 316922 640736 316927 640792
rect 55581 640734 316927 640736
rect 55581 640731 55647 640734
rect 316861 640731 316927 640734
rect 54937 640658 55003 640661
rect 315573 640658 315639 640661
rect 54937 640656 315639 640658
rect 54937 640600 54942 640656
rect 54998 640600 315578 640656
rect 315634 640600 315639 640656
rect 54937 640598 315639 640600
rect 54937 640595 55003 640598
rect 315573 640595 315639 640598
rect 35709 640522 35775 640525
rect 56501 640522 56567 640525
rect 35709 640520 56567 640522
rect 35709 640464 35714 640520
rect 35770 640464 56506 640520
rect 56562 640464 56567 640520
rect 35709 640462 56567 640464
rect 35709 640459 35775 640462
rect 56501 640459 56567 640462
rect 59169 640522 59235 640525
rect 379053 640522 379119 640525
rect 539593 640522 539659 640525
rect 59169 640520 379119 640522
rect 59169 640464 59174 640520
rect 59230 640464 379058 640520
rect 379114 640464 379119 640520
rect 59169 640462 379119 640464
rect 59169 640459 59235 640462
rect 379053 640459 379119 640462
rect 539550 640520 539659 640522
rect 539550 640464 539598 640520
rect 539654 640464 539659 640520
rect 539550 640459 539659 640464
rect 53373 640386 53439 640389
rect 59261 640386 59327 640389
rect 53373 640384 59327 640386
rect 53373 640328 53378 640384
rect 53434 640328 59266 640384
rect 59322 640328 59327 640384
rect 53373 640326 59327 640328
rect 53373 640323 53439 640326
rect 59261 640323 59327 640326
rect 177246 640324 177252 640388
rect 177316 640386 177322 640388
rect 177573 640386 177639 640389
rect 177316 640384 177639 640386
rect 177316 640328 177578 640384
rect 177634 640328 177639 640384
rect 177316 640326 177639 640328
rect 177316 640324 177322 640326
rect 177573 640323 177639 640326
rect 177798 640324 177804 640388
rect 177868 640386 177874 640388
rect 177941 640386 178007 640389
rect 177868 640384 178007 640386
rect 177868 640328 177946 640384
rect 178002 640328 178007 640384
rect 177868 640326 178007 640328
rect 177868 640324 177874 640326
rect 177941 640323 178007 640326
rect 249701 640386 249767 640389
rect 369669 640386 369735 640389
rect 249701 640384 369735 640386
rect 249701 640328 249706 640384
rect 249762 640328 369674 640384
rect 369730 640328 369735 640384
rect 539550 640356 539610 640459
rect 249701 640326 369735 640328
rect 249701 640323 249767 640326
rect 369669 640323 369735 640326
rect 297030 640188 297036 640252
rect 297100 640250 297106 640252
rect 298001 640250 298067 640253
rect 297100 640248 298067 640250
rect 297100 640192 298006 640248
rect 298062 640192 298067 640248
rect 297100 640190 298067 640192
rect 297100 640188 297106 640190
rect 298001 640187 298067 640190
rect 34329 640114 34395 640117
rect 88977 640114 89043 640117
rect 34329 640112 89043 640114
rect 34329 640056 34334 640112
rect 34390 640056 88982 640112
rect 89038 640056 89043 640112
rect 34329 640054 89043 640056
rect 34329 640051 34395 640054
rect 88977 640051 89043 640054
rect 50061 639978 50127 639981
rect 109033 639978 109099 639981
rect 50061 639976 109099 639978
rect 50061 639920 50066 639976
rect 50122 639920 109038 639976
rect 109094 639920 109099 639976
rect 50061 639918 109099 639920
rect 50061 639915 50127 639918
rect 109033 639915 109099 639918
rect 110321 639978 110387 639981
rect 154481 639978 154547 639981
rect 110321 639976 154547 639978
rect 110321 639920 110326 639976
rect 110382 639920 154486 639976
rect 154542 639920 154547 639976
rect 110321 639918 154547 639920
rect 110321 639915 110387 639918
rect 154481 639915 154547 639918
rect 66069 639842 66135 639845
rect 88241 639842 88307 639845
rect 66069 639840 88307 639842
rect 66069 639784 66074 639840
rect 66130 639784 88246 639840
rect 88302 639784 88307 639840
rect 66069 639782 88307 639784
rect 66069 639779 66135 639782
rect 88241 639779 88307 639782
rect 89713 639842 89779 639845
rect 107561 639842 107627 639845
rect 89713 639840 107627 639842
rect 89713 639784 89718 639840
rect 89774 639784 107566 639840
rect 107622 639784 107627 639840
rect 89713 639782 107627 639784
rect 89713 639779 89779 639782
rect 107561 639779 107627 639782
rect 153837 639842 153903 639845
rect 375465 639842 375531 639845
rect 153837 639840 375531 639842
rect 153837 639784 153842 639840
rect 153898 639784 375470 639840
rect 375526 639784 375531 639840
rect 153837 639782 375531 639784
rect 153837 639779 153903 639782
rect 375465 639779 375531 639782
rect 47894 639644 47900 639708
rect 47964 639706 47970 639708
rect 296846 639706 296852 639708
rect 47964 639646 296852 639706
rect 47964 639644 47970 639646
rect 296846 639644 296852 639646
rect 296916 639644 296922 639708
rect 52913 639570 52979 639573
rect 310421 639570 310487 639573
rect 52913 639568 310487 639570
rect 52913 639512 52918 639568
rect 52974 639512 310426 639568
rect 310482 639512 310487 639568
rect 52913 639510 310487 639512
rect 52913 639507 52979 639510
rect 310421 639507 310487 639510
rect 31518 639372 31524 639436
rect 31588 639434 31594 639436
rect 291878 639434 291884 639436
rect 31588 639374 291884 639434
rect 31588 639372 31594 639374
rect 291878 639372 291884 639374
rect 291948 639372 291954 639436
rect 294638 639372 294644 639436
rect 294708 639434 294714 639436
rect 478086 639434 478092 639436
rect 294708 639374 478092 639434
rect 294708 639372 294714 639374
rect 478086 639372 478092 639374
rect 478156 639372 478162 639436
rect 37181 639298 37247 639301
rect 307845 639298 307911 639301
rect 37181 639296 307911 639298
rect 37181 639240 37186 639296
rect 37242 639240 307850 639296
rect 307906 639240 307911 639296
rect 37181 639238 307911 639240
rect 37181 639235 37247 639238
rect 307845 639235 307911 639238
rect 87137 639162 87203 639165
rect 106181 639162 106247 639165
rect 87137 639160 106247 639162
rect 87137 639104 87142 639160
rect 87198 639104 106186 639160
rect 106242 639104 106247 639160
rect 87137 639102 106247 639104
rect 87137 639099 87203 639102
rect 106181 639099 106247 639102
rect 106457 639162 106523 639165
rect 418521 639162 418587 639165
rect 106457 639160 418587 639162
rect 106457 639104 106462 639160
rect 106518 639104 418526 639160
rect 418582 639104 418587 639160
rect 106457 639102 418587 639104
rect 106457 639099 106523 639102
rect 418521 639099 418587 639102
rect 45001 639026 45067 639029
rect 66161 639026 66227 639029
rect 45001 639024 66227 639026
rect 45001 638968 45006 639024
rect 45062 638968 66166 639024
rect 66222 638968 66227 639024
rect 45001 638966 66227 638968
rect 45001 638963 45067 638966
rect 66161 638963 66227 638966
rect 105169 639026 105235 639029
rect 417509 639026 417575 639029
rect 542353 639026 542419 639029
rect 105169 639024 417575 639026
rect 105169 638968 105174 639024
rect 105230 638968 417514 639024
rect 417570 638968 417575 639024
rect 105169 638966 417575 638968
rect 539948 639024 542419 639026
rect 539948 638968 542358 639024
rect 542414 638968 542419 639024
rect 539948 638966 542419 638968
rect 105169 638963 105235 638966
rect 417509 638963 417575 638966
rect 542353 638963 542419 638966
rect 102593 638890 102659 638893
rect 227713 638890 227779 638893
rect 102593 638888 227779 638890
rect 102593 638832 102598 638888
rect 102654 638832 227718 638888
rect 227774 638832 227779 638888
rect 102593 638830 227779 638832
rect 102593 638827 102659 638830
rect 227713 638827 227779 638830
rect 79409 638754 79475 638757
rect 118693 638754 118759 638757
rect 79409 638752 118759 638754
rect 79409 638696 79414 638752
rect 79470 638696 118698 638752
rect 118754 638696 118759 638752
rect 79409 638694 118759 638696
rect 79409 638691 79475 638694
rect 118693 638691 118759 638694
rect 137277 638754 137343 638757
rect 295977 638754 296043 638757
rect 137277 638752 296043 638754
rect 137277 638696 137282 638752
rect 137338 638696 295982 638752
rect 296038 638696 296043 638752
rect 137277 638694 296043 638696
rect 137277 638691 137343 638694
rect 295977 638691 296043 638694
rect 28533 638618 28599 638621
rect 86861 638618 86927 638621
rect 28533 638616 86927 638618
rect 28533 638560 28538 638616
rect 28594 638560 86866 638616
rect 86922 638560 86927 638616
rect 28533 638558 86927 638560
rect 28533 638555 28599 638558
rect 86861 638555 86927 638558
rect 111609 638618 111675 638621
rect 422569 638618 422635 638621
rect 111609 638616 422635 638618
rect 111609 638560 111614 638616
rect 111670 638560 422574 638616
rect 422630 638560 422635 638616
rect 111609 638558 422635 638560
rect 111609 638555 111675 638558
rect 422569 638555 422635 638558
rect 85849 638482 85915 638485
rect 129733 638482 129799 638485
rect 85849 638480 129799 638482
rect 85849 638424 85854 638480
rect 85910 638424 129738 638480
rect 129794 638424 129799 638480
rect 85849 638422 129799 638424
rect 85849 638419 85915 638422
rect 129733 638419 129799 638422
rect 179137 638482 179203 638485
rect 258717 638482 258783 638485
rect 179137 638480 258783 638482
rect 179137 638424 179142 638480
rect 179198 638424 258722 638480
rect 258778 638424 258783 638480
rect 179137 638422 258783 638424
rect 179137 638419 179203 638422
rect 258717 638419 258783 638422
rect 78121 638346 78187 638349
rect 82813 638346 82879 638349
rect 78121 638344 82879 638346
rect 78121 638288 78126 638344
rect 78182 638288 82818 638344
rect 82874 638288 82879 638344
rect 78121 638286 82879 638288
rect 78121 638283 78187 638286
rect 82813 638283 82879 638286
rect 83273 638346 83339 638349
rect 102133 638346 102199 638349
rect 83273 638344 102199 638346
rect 83273 638288 83278 638344
rect 83334 638288 102138 638344
rect 102194 638288 102199 638344
rect 83273 638286 102199 638288
rect 83273 638283 83339 638286
rect 102133 638283 102199 638286
rect 227897 638346 227963 638349
rect 250897 638346 250963 638349
rect 258073 638346 258139 638349
rect 259361 638346 259427 638349
rect 227897 638344 259427 638346
rect 227897 638288 227902 638344
rect 227958 638288 250902 638344
rect 250958 638288 258078 638344
rect 258134 638288 259366 638344
rect 259422 638288 259427 638344
rect 227897 638286 259427 638288
rect 227897 638283 227963 638286
rect 250897 638283 250963 638286
rect 258073 638283 258139 638286
rect 259361 638283 259427 638286
rect 35801 638210 35867 638213
rect 81433 638210 81499 638213
rect 35801 638208 81499 638210
rect 35801 638152 35806 638208
rect 35862 638152 81438 638208
rect 81494 638152 81499 638208
rect 35801 638150 81499 638152
rect 35801 638147 35867 638150
rect 81433 638147 81499 638150
rect 119337 638210 119403 638213
rect 256601 638210 256667 638213
rect 119337 638208 256667 638210
rect 119337 638152 119342 638208
rect 119398 638152 256606 638208
rect 256662 638152 256667 638208
rect 119337 638150 256667 638152
rect 119337 638147 119403 638150
rect 256601 638147 256667 638150
rect 32949 638074 33015 638077
rect 137277 638074 137343 638077
rect 32949 638072 137343 638074
rect 32949 638016 32954 638072
rect 33010 638016 137282 638072
rect 137338 638016 137343 638072
rect 32949 638014 137343 638016
rect 32949 638011 33015 638014
rect 137277 638011 137343 638014
rect 294454 638012 294460 638076
rect 294524 638074 294530 638076
rect 482134 638074 482140 638076
rect 294524 638014 482140 638074
rect 294524 638012 294530 638014
rect 482134 638012 482140 638014
rect 482204 638012 482210 638076
rect 34278 637876 34284 637940
rect 34348 637938 34354 637940
rect 291694 637938 291700 637940
rect 34348 637878 291700 637938
rect 34348 637876 34354 637878
rect 291694 637876 291700 637878
rect 291764 637876 291770 637940
rect 292062 637876 292068 637940
rect 292132 637938 292138 637940
rect 483606 637938 483612 637940
rect 292132 637878 483612 637938
rect 292132 637876 292138 637878
rect 483606 637876 483612 637878
rect 483676 637876 483682 637940
rect 50705 637802 50771 637805
rect 311709 637802 311775 637805
rect 539961 637802 540027 637805
rect 50705 637800 311775 637802
rect 50705 637744 50710 637800
rect 50766 637744 311714 637800
rect 311770 637744 311775 637800
rect 50705 637742 311775 637744
rect 50705 637739 50771 637742
rect 311709 637739 311775 637742
rect 539918 637800 540027 637802
rect 539918 637744 539966 637800
rect 540022 637744 540027 637800
rect 539918 637739 540027 637744
rect 81985 637666 82051 637669
rect 110413 637666 110479 637669
rect 81985 637664 110479 637666
rect 81985 637608 81990 637664
rect 82046 637608 110418 637664
rect 110474 637608 110479 637664
rect 81985 637606 110479 637608
rect 81985 637603 82051 637606
rect 110413 637603 110479 637606
rect 130929 637666 130995 637669
rect 130929 637664 138122 637666
rect 130929 637608 130934 637664
rect 130990 637608 138122 637664
rect 130929 637606 138122 637608
rect 130929 637603 130995 637606
rect 50889 637530 50955 637533
rect 121453 637530 121519 637533
rect 50889 637528 121519 637530
rect 50889 637472 50894 637528
rect 50950 637472 121458 637528
rect 121514 637472 121519 637528
rect 50889 637470 121519 637472
rect 138062 637530 138122 637606
rect 177430 637604 177436 637668
rect 177500 637666 177506 637668
rect 179045 637666 179111 637669
rect 177500 637664 179111 637666
rect 177500 637608 179050 637664
rect 179106 637608 179111 637664
rect 539918 637636 539978 637739
rect 177500 637606 179111 637608
rect 177500 637604 177506 637606
rect 179045 637603 179111 637606
rect 227897 637530 227963 637533
rect 138062 637528 227963 637530
rect 138062 637472 227902 637528
rect 227958 637472 227963 637528
rect 138062 637470 227963 637472
rect 50889 637467 50955 637470
rect 121453 637467 121519 637470
rect 227897 637467 227963 637470
rect 540237 637530 540303 637533
rect 542721 637530 542787 637533
rect 540237 637528 542787 637530
rect 540237 637472 540242 637528
rect 540298 637472 542726 637528
rect 542782 637472 542787 637528
rect 540237 637470 542787 637472
rect 540237 637467 540303 637470
rect 542721 637467 542787 637470
rect 58525 637394 58591 637397
rect 237281 637394 237347 637397
rect 242801 637394 242867 637397
rect 58525 637392 161490 637394
rect 58525 637336 58530 637392
rect 58586 637336 161490 637392
rect 58525 637334 161490 637336
rect 58525 637331 58591 637334
rect 32990 637196 32996 637260
rect 33060 637258 33066 637260
rect 128353 637258 128419 637261
rect 33060 637256 128419 637258
rect 33060 637200 128358 637256
rect 128414 637200 128419 637256
rect 33060 637198 128419 637200
rect 161430 637258 161490 637334
rect 237281 637392 242867 637394
rect 237281 637336 237286 637392
rect 237342 637336 242806 637392
rect 242862 637336 242867 637392
rect 237281 637334 242867 637336
rect 237281 637331 237347 637334
rect 242801 637331 242867 637334
rect 175089 637258 175155 637261
rect 260189 637258 260255 637261
rect 161430 637256 260255 637258
rect 161430 637200 175094 637256
rect 175150 637200 260194 637256
rect 260250 637200 260255 637256
rect 161430 637198 260255 637200
rect 33060 637196 33066 637198
rect 128353 637195 128419 637198
rect 175089 637195 175155 637198
rect 260189 637195 260255 637198
rect 74257 637122 74323 637125
rect 108297 637122 108363 637125
rect 74257 637120 108363 637122
rect 74257 637064 74262 637120
rect 74318 637064 108302 637120
rect 108358 637064 108363 637120
rect 74257 637062 108363 637064
rect 74257 637059 74323 637062
rect 108297 637059 108363 637062
rect 178902 637060 178908 637124
rect 178972 637122 178978 637124
rect 191741 637122 191807 637125
rect 240041 637122 240107 637125
rect 178972 637062 190470 637122
rect 178972 637060 178978 637062
rect 70393 636986 70459 636989
rect 117221 636986 117287 636989
rect 135989 636986 136055 636989
rect 70393 636984 117287 636986
rect 70393 636928 70398 636984
rect 70454 636928 117226 636984
rect 117282 636928 117287 636984
rect 70393 636926 117287 636928
rect 70393 636923 70459 636926
rect 117221 636923 117287 636926
rect 117454 636984 136055 636986
rect 117454 636928 135994 636984
rect 136050 636928 136055 636984
rect 117454 636926 136055 636928
rect 116761 636850 116827 636853
rect 117454 636850 117514 636926
rect 135989 636923 136055 636926
rect 177757 636986 177823 636989
rect 190410 636986 190470 637062
rect 191741 637120 240107 637122
rect 191741 637064 191746 637120
rect 191802 637064 240046 637120
rect 240102 637064 240107 637120
rect 191741 637062 240107 637064
rect 191741 637059 191807 637062
rect 240041 637059 240107 637062
rect 245009 637122 245075 637125
rect 247125 637122 247191 637125
rect 245009 637120 247191 637122
rect 245009 637064 245014 637120
rect 245070 637064 247130 637120
rect 247186 637064 247191 637120
rect 245009 637062 247191 637064
rect 245009 637059 245075 637062
rect 247125 637059 247191 637062
rect 235993 636986 236059 636989
rect 177757 636984 180810 636986
rect 177757 636928 177762 636984
rect 177818 636928 180810 636984
rect 177757 636926 180810 636928
rect 190410 636984 236059 636986
rect 190410 636928 235998 636984
rect 236054 636928 236059 636984
rect 190410 636926 236059 636928
rect 177757 636923 177823 636926
rect 116761 636848 117514 636850
rect 116761 636792 116766 636848
rect 116822 636792 117514 636848
rect 116761 636790 117514 636792
rect 118049 636850 118115 636853
rect 176653 636850 176719 636853
rect 118049 636848 176719 636850
rect 118049 636792 118054 636848
rect 118110 636792 176658 636848
rect 176714 636792 176719 636848
rect 118049 636790 176719 636792
rect 180750 636850 180810 636926
rect 235993 636923 236059 636926
rect 242433 636986 242499 636989
rect 465901 636986 465967 636989
rect 242433 636984 465967 636986
rect 242433 636928 242438 636984
rect 242494 636928 465906 636984
rect 465962 636928 465967 636984
rect 242433 636926 465967 636928
rect 242433 636923 242499 636926
rect 465901 636923 465967 636926
rect 191741 636850 191807 636853
rect 180750 636848 191807 636850
rect 180750 636792 191746 636848
rect 191802 636792 191807 636848
rect 180750 636790 191807 636792
rect 116761 636787 116827 636790
rect 118049 636787 118115 636790
rect 176653 636787 176719 636790
rect 191741 636787 191807 636790
rect 229461 636850 229527 636853
rect 287697 636850 287763 636853
rect 229461 636848 287763 636850
rect 229461 636792 229466 636848
rect 229522 636792 287702 636848
rect 287758 636792 287763 636848
rect 229461 636790 287763 636792
rect 229461 636787 229527 636790
rect 287697 636787 287763 636790
rect 48078 636652 48084 636716
rect 48148 636714 48154 636716
rect 128445 636714 128511 636717
rect 48148 636712 128511 636714
rect 48148 636656 128450 636712
rect 128506 636656 128511 636712
rect 48148 636654 128511 636656
rect 48148 636652 48154 636654
rect 128445 636651 128511 636654
rect 128813 636714 128879 636717
rect 133873 636714 133939 636717
rect 128813 636712 133939 636714
rect 128813 636656 128818 636712
rect 128874 636656 133878 636712
rect 133934 636656 133939 636712
rect 128813 636654 133939 636656
rect 128813 636651 128879 636654
rect 133873 636651 133939 636654
rect 137369 636714 137435 636717
rect 296161 636714 296227 636717
rect 137369 636712 296227 636714
rect 137369 636656 137374 636712
rect 137430 636656 296166 636712
rect 296222 636656 296227 636712
rect 137369 636654 296227 636656
rect 137369 636651 137435 636654
rect 296161 636651 296227 636654
rect 48446 636516 48452 636580
rect 48516 636578 48522 636580
rect 125501 636578 125567 636581
rect 48516 636576 125567 636578
rect 48516 636520 125506 636576
rect 125562 636520 125567 636576
rect 48516 636518 125567 636520
rect 48516 636516 48522 636518
rect 125501 636515 125567 636518
rect 125685 636578 125751 636581
rect 237373 636578 237439 636581
rect 125685 636576 237439 636578
rect 125685 636520 125690 636576
rect 125746 636520 237378 636576
rect 237434 636520 237439 636576
rect 125685 636518 237439 636520
rect 125685 636515 125751 636518
rect 237373 636515 237439 636518
rect 239673 636578 239739 636581
rect 246941 636578 247007 636581
rect 239673 636576 247007 636578
rect 239673 636520 239678 636576
rect 239734 636520 246946 636576
rect 247002 636520 247007 636576
rect 239673 636518 247007 636520
rect 239673 636515 239739 636518
rect 246941 636515 247007 636518
rect 247125 636578 247191 636581
rect 468569 636578 468635 636581
rect 247125 636576 468635 636578
rect 247125 636520 247130 636576
rect 247186 636520 468574 636576
rect 468630 636520 468635 636576
rect 247125 636518 468635 636520
rect 247125 636515 247191 636518
rect 468569 636515 468635 636518
rect 121913 636442 121979 636445
rect 136173 636442 136239 636445
rect 121913 636440 136239 636442
rect 121913 636384 121918 636440
rect 121974 636384 136178 636440
rect 136234 636384 136239 636440
rect 121913 636382 136239 636384
rect 121913 636379 121979 636382
rect 136173 636379 136239 636382
rect 179086 636380 179092 636444
rect 179156 636442 179162 636444
rect 179321 636442 179387 636445
rect 179156 636440 179387 636442
rect 179156 636384 179326 636440
rect 179382 636384 179387 636440
rect 179156 636382 179387 636384
rect 179156 636380 179162 636382
rect 179321 636379 179387 636382
rect 238385 636442 238451 636445
rect 245561 636442 245627 636445
rect 238385 636440 245627 636442
rect 238385 636384 238390 636440
rect 238446 636384 245566 636440
rect 245622 636384 245627 636440
rect 238385 636382 245627 636384
rect 238385 636379 238451 636382
rect 245561 636379 245627 636382
rect 246113 636442 246179 636445
rect 470041 636442 470107 636445
rect 246113 636440 470107 636442
rect 246113 636384 246118 636440
rect 246174 636384 470046 636440
rect 470102 636384 470107 636440
rect 246113 636382 470107 636384
rect 246113 636379 246179 636382
rect 470041 636379 470107 636382
rect 63953 636306 64019 636309
rect 66069 636306 66135 636309
rect 63953 636304 66135 636306
rect 63953 636248 63958 636304
rect 64014 636248 66074 636304
rect 66130 636248 66135 636304
rect 63953 636246 66135 636248
rect 63953 636243 64019 636246
rect 66069 636243 66135 636246
rect 69105 636306 69171 636309
rect 73153 636306 73219 636309
rect 69105 636304 73219 636306
rect 69105 636248 69110 636304
rect 69166 636248 73158 636304
rect 73214 636248 73219 636304
rect 69105 636246 73219 636248
rect 69105 636243 69171 636246
rect 73153 636243 73219 636246
rect 107745 636306 107811 636309
rect 117957 636306 118023 636309
rect 107745 636304 118023 636306
rect 107745 636248 107750 636304
rect 107806 636248 117962 636304
rect 118018 636248 118023 636304
rect 107745 636246 118023 636248
rect 107745 636243 107811 636246
rect 117957 636243 118023 636246
rect 129641 636306 129707 636309
rect 249701 636306 249767 636309
rect 129641 636304 249767 636306
rect 129641 636248 129646 636304
rect 129702 636248 249706 636304
rect 249762 636248 249767 636304
rect 129641 636246 249767 636248
rect 129641 636243 129707 636246
rect 249701 636243 249767 636246
rect 369669 636306 369735 636309
rect 374453 636306 374519 636309
rect 542445 636306 542511 636309
rect 369669 636304 374519 636306
rect 369669 636248 369674 636304
rect 369730 636248 374458 636304
rect 374514 636248 374519 636304
rect 369669 636246 374519 636248
rect 539948 636304 542511 636306
rect 539948 636248 542450 636304
rect 542506 636248 542511 636304
rect 539948 636246 542511 636248
rect 369669 636243 369735 636246
rect 374453 636243 374519 636246
rect 542445 636243 542511 636246
rect 98729 636034 98795 636037
rect 109125 636034 109191 636037
rect 98729 636032 109191 636034
rect 98729 635976 98734 636032
rect 98790 635976 109130 636032
rect 109186 635976 109191 636032
rect 98729 635974 109191 635976
rect 98729 635971 98795 635974
rect 109125 635971 109191 635974
rect 55990 635836 55996 635900
rect 56060 635898 56066 635900
rect 377806 635898 377812 635900
rect 56060 635838 377812 635898
rect 56060 635836 56066 635838
rect 377806 635836 377812 635838
rect 377876 635836 377882 635900
rect 57697 635762 57763 635765
rect 176653 635762 176719 635765
rect 255589 635762 255655 635765
rect 57697 635760 175106 635762
rect 57697 635704 57702 635760
rect 57758 635704 175106 635760
rect 57697 635702 175106 635704
rect 57697 635699 57763 635702
rect 56041 635626 56107 635629
rect 173893 635626 173959 635629
rect 56041 635624 173959 635626
rect 56041 635568 56046 635624
rect 56102 635568 173898 635624
rect 173954 635568 173959 635624
rect 56041 635566 173959 635568
rect 175046 635626 175106 635702
rect 176653 635760 255655 635762
rect 176653 635704 176658 635760
rect 176714 635704 255594 635760
rect 255650 635704 255655 635760
rect 176653 635702 255655 635704
rect 176653 635699 176719 635702
rect 255589 635699 255655 635702
rect 178953 635626 179019 635629
rect 185669 635626 185735 635629
rect 258901 635626 258967 635629
rect 175046 635624 185594 635626
rect 175046 635568 178958 635624
rect 179014 635568 185594 635624
rect 175046 635566 185594 635568
rect 56041 635563 56107 635566
rect 173893 635563 173959 635566
rect 178953 635563 179019 635566
rect 54661 635490 54727 635493
rect 179229 635490 179295 635493
rect 185393 635490 185459 635493
rect 54661 635488 185459 635490
rect 54661 635432 54666 635488
rect 54722 635432 179234 635488
rect 179290 635432 185398 635488
rect 185454 635432 185459 635488
rect 54661 635430 185459 635432
rect 185534 635490 185594 635566
rect 185669 635624 258967 635626
rect 185669 635568 185674 635624
rect 185730 635568 258906 635624
rect 258962 635568 258967 635624
rect 185669 635566 258967 635568
rect 185669 635563 185735 635566
rect 258901 635563 258967 635566
rect 260281 635490 260347 635493
rect 185534 635488 260347 635490
rect 185534 635432 260286 635488
rect 260342 635432 260347 635488
rect 185534 635430 260347 635432
rect 54661 635427 54727 635430
rect 179229 635427 179295 635430
rect 185393 635427 185459 635430
rect 260281 635427 260347 635430
rect 296662 635428 296668 635492
rect 296732 635490 296738 635492
rect 297817 635490 297883 635493
rect 296732 635488 297883 635490
rect 296732 635432 297822 635488
rect 297878 635432 297883 635488
rect 296732 635430 297883 635432
rect 296732 635428 296738 635430
rect 297817 635427 297883 635430
rect 47710 635292 47716 635356
rect 47780 635354 47786 635356
rect 296478 635354 296484 635356
rect 47780 635294 296484 635354
rect 47780 635292 47786 635294
rect 296478 635292 296484 635294
rect 296548 635292 296554 635356
rect 65241 635218 65307 635221
rect 95141 635218 95207 635221
rect 65241 635216 95207 635218
rect 65241 635160 65246 635216
rect 65302 635160 95146 635216
rect 95202 635160 95207 635216
rect 65241 635158 95207 635160
rect 65241 635155 65307 635158
rect 95141 635155 95207 635158
rect 109033 635218 109099 635221
rect 393957 635218 394023 635221
rect 109033 635216 394023 635218
rect 109033 635160 109038 635216
rect 109094 635160 393962 635216
rect 394018 635160 394023 635216
rect 109033 635158 394023 635160
rect 109033 635155 109099 635158
rect 393957 635155 394023 635158
rect 38469 635082 38535 635085
rect 92473 635082 92539 635085
rect 38469 635080 92539 635082
rect 38469 635024 38474 635080
rect 38530 635024 92478 635080
rect 92534 635024 92539 635080
rect 38469 635022 92539 635024
rect 38469 635019 38535 635022
rect 92473 635019 92539 635022
rect 93761 635082 93827 635085
rect 99373 635082 99439 635085
rect 93761 635080 99439 635082
rect 93761 635024 93766 635080
rect 93822 635024 99378 635080
rect 99434 635024 99439 635080
rect 93761 635022 99439 635024
rect 93761 635019 93827 635022
rect 99373 635019 99439 635022
rect 104249 635082 104315 635085
rect 416497 635082 416563 635085
rect 104249 635080 416563 635082
rect 104249 635024 104254 635080
rect 104310 635024 416502 635080
rect 416558 635024 416563 635080
rect 104249 635022 416563 635024
rect 104249 635019 104315 635022
rect 416497 635019 416563 635022
rect 94865 634946 94931 634949
rect 98085 634946 98151 634949
rect 94865 634944 98151 634946
rect 94865 634888 94870 634944
rect 94926 634888 98090 634944
rect 98146 634888 98151 634944
rect 94865 634886 98151 634888
rect 94865 634883 94931 634886
rect 98085 634883 98151 634886
rect 100017 634946 100083 634949
rect 104801 634946 104867 634949
rect 100017 634944 104867 634946
rect 100017 634888 100022 634944
rect 100078 634888 104806 634944
rect 104862 634888 104867 634944
rect 100017 634886 104867 634888
rect 100017 634883 100083 634886
rect 104801 634883 104867 634886
rect 58341 634810 58407 634813
rect 174721 634810 174787 634813
rect 179137 634810 179203 634813
rect 58341 634808 179203 634810
rect 58341 634752 58346 634808
rect 58402 634752 174726 634808
rect 174782 634752 179142 634808
rect 179198 634752 179203 634808
rect 58341 634750 179203 634752
rect 58341 634747 58407 634750
rect 174721 634747 174787 634750
rect 179137 634747 179203 634750
rect 248367 634810 248433 634813
rect 285029 634810 285095 634813
rect 248367 634808 285095 634810
rect 248367 634752 248372 634808
rect 248428 634752 285034 634808
rect 285090 634752 285095 634808
rect 248367 634750 285095 634752
rect 248367 634747 248433 634750
rect 285029 634747 285095 634750
rect 539734 634677 539794 634916
rect 54569 634674 54635 634677
rect 175181 634674 175247 634677
rect 54569 634672 175247 634674
rect 54569 634616 54574 634672
rect 54630 634616 175186 634672
rect 175242 634616 175247 634672
rect 54569 634614 175247 634616
rect 54569 634611 54635 634614
rect 175181 634611 175247 634614
rect 237373 634674 237439 634677
rect 260649 634674 260715 634677
rect 237373 634672 260715 634674
rect 237373 634616 237378 634672
rect 237434 634616 260654 634672
rect 260710 634616 260715 634672
rect 237373 634614 260715 634616
rect 237373 634611 237439 634614
rect 260649 634611 260715 634614
rect 539685 634672 539794 634677
rect 539685 634616 539690 634672
rect 539746 634616 539794 634672
rect 539685 634614 539794 634616
rect 539685 634611 539751 634614
rect 133873 634538 133939 634541
rect 263685 634538 263751 634541
rect 133873 634536 263751 634538
rect 133873 634480 133878 634536
rect 133934 634480 263690 634536
rect 263746 634480 263751 634536
rect 133873 634478 263751 634480
rect 133873 634475 133939 634478
rect 263685 634475 263751 634478
rect 304257 634538 304323 634541
rect 392577 634538 392643 634541
rect 304257 634536 392643 634538
rect 304257 634480 304262 634536
rect 304318 634480 392582 634536
rect 392638 634480 392643 634536
rect 304257 634478 392643 634480
rect 304257 634475 304323 634478
rect 392577 634475 392643 634478
rect 299657 634402 299723 634405
rect 302693 634402 302759 634405
rect 299657 634400 302759 634402
rect 299657 634344 299662 634400
rect 299718 634344 302698 634400
rect 302754 634344 302759 634400
rect 299657 634342 302759 634344
rect 299657 634339 299723 634342
rect 302693 634339 302759 634342
rect 120625 634266 120691 634269
rect 243215 634266 243281 634269
rect 303981 634266 304047 634269
rect 120625 634264 122850 634266
rect 120625 634208 120630 634264
rect 120686 634208 122850 634264
rect 120625 634206 122850 634208
rect 120625 634203 120691 634206
rect 122790 634130 122850 634206
rect 243215 634264 244290 634266
rect 243215 634208 243220 634264
rect 243276 634208 244290 634264
rect 243215 634206 244290 634208
rect 243215 634203 243281 634206
rect 127566 634130 127572 634132
rect 122790 634070 127572 634130
rect 127566 634068 127572 634070
rect 127636 634068 127642 634132
rect 244230 634130 244290 634206
rect 296670 634264 304047 634266
rect 296670 634208 303986 634264
rect 304042 634208 304047 634264
rect 296670 634206 304047 634208
rect 249006 634130 249012 634132
rect 244230 634070 249012 634130
rect 249006 634068 249012 634070
rect 249076 634068 249082 634132
rect 28717 633994 28783 633997
rect 296670 633994 296730 634206
rect 303981 634203 304047 634206
rect 299657 633994 299723 633997
rect 28717 633992 296730 633994
rect 28717 633936 28722 633992
rect 28778 633936 296730 633992
rect 28717 633934 296730 633936
rect 299614 633992 299723 633994
rect 299614 633936 299662 633992
rect 299718 633936 299723 633992
rect 28717 633931 28783 633934
rect 299614 633931 299723 633936
rect 28809 633858 28875 633861
rect 299614 633858 299674 633931
rect 28809 633856 299674 633858
rect 28809 633800 28814 633856
rect 28870 633800 299674 633856
rect 28809 633798 299674 633800
rect 28809 633795 28875 633798
rect 127566 633660 127572 633724
rect 127636 633722 127642 633724
rect 178769 633722 178835 633725
rect 127636 633720 178835 633722
rect 127636 633664 178774 633720
rect 178830 633664 178835 633720
rect 127636 633662 178835 633664
rect 127636 633660 127642 633662
rect 178769 633659 178835 633662
rect 249006 633660 249012 633724
rect 249076 633722 249082 633724
rect 489269 633722 489335 633725
rect 249076 633720 489335 633722
rect 249076 633664 489274 633720
rect 489330 633664 489335 633720
rect 249076 633662 489335 633664
rect 249076 633660 249082 633662
rect 489269 633659 489335 633662
rect 175181 633586 175247 633589
rect 179137 633586 179203 633589
rect 542537 633586 542603 633589
rect 175181 633584 180810 633586
rect 175181 633528 175186 633584
rect 175242 633528 179142 633584
rect 179198 633528 180810 633584
rect 175181 633526 180810 633528
rect 539948 633584 542603 633586
rect 539948 633528 542542 633584
rect 542598 633528 542603 633584
rect 539948 633526 542603 633528
rect 175181 633523 175247 633526
rect 179137 633523 179203 633526
rect 179965 633450 180031 633453
rect 180750 633450 180810 633526
rect 542537 633523 542603 633526
rect 255957 633450 256023 633453
rect 179965 633448 180074 633450
rect 179965 633392 179970 633448
rect 180026 633392 180074 633448
rect 179965 633387 180074 633392
rect 180750 633448 256023 633450
rect 180750 633392 255962 633448
rect 256018 633392 256023 633448
rect 180750 633390 256023 633392
rect 255957 633387 256023 633390
rect 59077 633314 59143 633317
rect 59077 633312 60076 633314
rect 59077 633256 59082 633312
rect 59138 633256 60076 633312
rect 180014 633284 180074 633387
rect 297265 633314 297331 633317
rect 297265 633312 300196 633314
rect 59077 633254 60076 633256
rect 297265 633256 297270 633312
rect 297326 633256 300196 633312
rect 297265 633254 300196 633256
rect 59077 633251 59143 633254
rect 297265 633251 297331 633254
rect 374453 632634 374519 632637
rect 480897 632634 480963 632637
rect 374453 632632 480963 632634
rect 374453 632576 374458 632632
rect 374514 632576 480902 632632
rect 480958 632576 480963 632632
rect 374453 632574 480963 632576
rect 374453 632571 374519 632574
rect 480897 632571 480963 632574
rect 59261 632226 59327 632229
rect 59261 632224 59554 632226
rect -960 632090 480 632180
rect 59261 632168 59266 632224
rect 59322 632168 59554 632224
rect 59261 632166 59554 632168
rect 59261 632163 59327 632166
rect 59494 632158 59554 632166
rect 179270 632164 179276 632228
rect 179340 632226 179346 632228
rect 297909 632226 297975 632229
rect 540237 632226 540303 632229
rect 179340 632166 180044 632226
rect 297909 632224 299674 632226
rect 297909 632168 297914 632224
rect 297970 632168 299674 632224
rect 297909 632166 299674 632168
rect 539948 632224 540303 632226
rect 539948 632168 540242 632224
rect 540298 632168 540303 632224
rect 539948 632166 540303 632168
rect 179340 632164 179346 632166
rect 297909 632163 297975 632166
rect 299614 632158 299674 632166
rect 540237 632163 540303 632166
rect 59494 632098 60076 632158
rect 299614 632098 300196 632158
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 57789 631138 57855 631141
rect 57789 631136 59554 631138
rect 57789 631080 57794 631136
rect 57850 631080 59554 631136
rect 57789 631078 59554 631080
rect 57789 631075 57855 631078
rect 59494 631070 59554 631078
rect 179086 631076 179092 631140
rect 179156 631138 179162 631140
rect 297725 631138 297791 631141
rect 179156 631078 180044 631138
rect 297725 631136 299674 631138
rect 297725 631080 297730 631136
rect 297786 631080 299674 631136
rect 297725 631078 299674 631080
rect 179156 631076 179162 631078
rect 297725 631075 297791 631078
rect 299614 631070 299674 631078
rect 59494 631010 60076 631070
rect 299614 631010 300196 631070
rect 542629 630866 542695 630869
rect 539948 630864 542695 630866
rect 539948 630808 542634 630864
rect 542690 630808 542695 630864
rect 539948 630806 542695 630808
rect 542629 630803 542695 630806
rect 555366 630804 555372 630868
rect 555436 630866 555442 630868
rect 583520 630866 584960 630956
rect 555436 630806 584960 630866
rect 555436 630804 555442 630806
rect 583520 630716 584960 630806
rect 59169 630050 59235 630053
rect 177757 630050 177823 630053
rect 298001 630050 298067 630053
rect 542721 630050 542787 630053
rect 544377 630050 544443 630053
rect 59169 630048 59554 630050
rect 59169 629992 59174 630048
rect 59230 629992 59554 630048
rect 59169 629990 59554 629992
rect 59169 629987 59235 629990
rect 59494 629982 59554 629990
rect 177757 630048 180044 630050
rect 177757 629992 177762 630048
rect 177818 629992 180044 630048
rect 177757 629990 180044 629992
rect 298001 630048 299674 630050
rect 298001 629992 298006 630048
rect 298062 629992 299674 630048
rect 298001 629990 299674 629992
rect 177757 629987 177823 629990
rect 298001 629987 298067 629990
rect 299614 629982 299674 629990
rect 542721 630048 544443 630050
rect 542721 629992 542726 630048
rect 542782 629992 544382 630048
rect 544438 629992 544443 630048
rect 542721 629990 544443 629992
rect 542721 629987 542787 629990
rect 544377 629987 544443 629990
rect 59494 629922 60076 629982
rect 299614 629922 300196 629982
rect 542721 629506 542787 629509
rect 539948 629504 542787 629506
rect 539948 629448 542726 629504
rect 542782 629448 542787 629504
rect 539948 629446 542787 629448
rect 542721 629443 542787 629446
rect 178902 628900 178908 628964
rect 178972 628962 178978 628964
rect 297541 628962 297607 628965
rect 178972 628902 180044 628962
rect 297541 628960 299674 628962
rect 297541 628904 297546 628960
rect 297602 628904 299674 628960
rect 297541 628902 299674 628904
rect 178972 628900 178978 628902
rect 297541 628899 297607 628902
rect 299614 628894 299674 628902
rect 59494 628834 60076 628894
rect 299614 628834 300196 628894
rect 57646 628764 57652 628828
rect 57716 628826 57722 628828
rect 59494 628826 59554 628834
rect 57716 628766 59554 628826
rect 57716 628764 57722 628766
rect 540145 628146 540211 628149
rect 539948 628144 540211 628146
rect 539948 628088 540150 628144
rect 540206 628088 540211 628144
rect 539948 628086 540211 628088
rect 540145 628083 540211 628086
rect 177849 627874 177915 627877
rect 297633 627874 297699 627877
rect 177849 627872 180044 627874
rect 177849 627816 177854 627872
rect 177910 627816 180044 627872
rect 177849 627814 180044 627816
rect 297633 627872 299674 627874
rect 297633 627816 297638 627872
rect 297694 627816 299674 627872
rect 297633 627814 299674 627816
rect 177849 627811 177915 627814
rect 297633 627811 297699 627814
rect 299614 627806 299674 627814
rect 59494 627746 60076 627806
rect 299614 627746 300196 627806
rect 57830 627676 57836 627740
rect 57900 627738 57906 627740
rect 59494 627738 59554 627746
rect 57900 627678 59554 627738
rect 57900 627676 57906 627678
rect 177665 626786 177731 626789
rect 297817 626786 297883 626789
rect 542813 626786 542879 626789
rect 177665 626784 180044 626786
rect 177665 626728 177670 626784
rect 177726 626728 180044 626784
rect 177665 626726 180044 626728
rect 297817 626784 299674 626786
rect 297817 626728 297822 626784
rect 297878 626728 299674 626784
rect 297817 626726 299674 626728
rect 539948 626784 542879 626786
rect 539948 626728 542818 626784
rect 542874 626728 542879 626784
rect 539948 626726 542879 626728
rect 177665 626723 177731 626726
rect 297817 626723 297883 626726
rect 299614 626718 299674 626726
rect 542813 626723 542879 626726
rect 59494 626658 60076 626718
rect 299614 626658 300196 626718
rect 58934 626588 58940 626652
rect 59004 626650 59010 626652
rect 59494 626650 59554 626658
rect 59004 626590 59554 626650
rect 59004 626588 59010 626590
rect 166349 626514 166415 626517
rect 291142 626514 291148 626516
rect 142110 626512 166415 626514
rect 134934 626378 134994 626484
rect 142110 626456 166354 626512
rect 166410 626456 166415 626512
rect 142110 626454 166415 626456
rect 254932 626454 291148 626514
rect 142110 626378 142170 626454
rect 166349 626451 166415 626454
rect 291142 626452 291148 626454
rect 291212 626452 291218 626516
rect 377622 626514 377628 626516
rect 374900 626454 377628 626514
rect 377622 626452 377628 626454
rect 377692 626452 377698 626516
rect 134934 626318 142170 626378
rect 137369 626242 137435 626245
rect 374729 626242 374795 626245
rect 134934 626240 137435 626242
rect 134934 626184 137374 626240
rect 137430 626184 137435 626240
rect 134934 626182 137435 626184
rect 57881 625698 57947 625701
rect 57881 625696 60076 625698
rect 57881 625640 57886 625696
rect 57942 625640 60076 625696
rect 134934 625668 134994 626182
rect 137369 626179 137435 626182
rect 374686 626240 374795 626242
rect 374686 626184 374734 626240
rect 374790 626184 374795 626240
rect 374686 626179 374795 626184
rect 57881 625638 60076 625640
rect 57881 625635 57947 625638
rect 176142 625636 176148 625700
rect 176212 625698 176218 625700
rect 294781 625698 294847 625701
rect 176212 625638 180044 625698
rect 254932 625696 294847 625698
rect 254932 625640 294786 625696
rect 294842 625640 294847 625696
rect 254932 625638 294847 625640
rect 176212 625636 176218 625638
rect 294781 625635 294847 625638
rect 296846 625636 296852 625700
rect 296916 625698 296922 625700
rect 296916 625638 300196 625698
rect 374686 625668 374746 626179
rect 296916 625636 296922 625638
rect 539734 625021 539794 625396
rect 374545 625018 374611 625021
rect 374502 625016 374611 625018
rect 374502 624960 374550 625016
rect 374606 624960 374611 625016
rect 374502 624955 374611 624960
rect 539734 625016 539843 625021
rect 539734 624960 539782 625016
rect 539838 624960 539843 625016
rect 539734 624958 539843 624960
rect 539777 624955 539843 624958
rect 169017 624882 169083 624885
rect 294597 624882 294663 624885
rect 142110 624880 169083 624882
rect 134934 624746 134994 624852
rect 142110 624824 169022 624880
rect 169078 624824 169083 624880
rect 142110 624822 169083 624824
rect 254932 624880 294663 624882
rect 254932 624824 294602 624880
rect 294658 624824 294663 624880
rect 374502 624852 374562 624955
rect 254932 624822 294663 624824
rect 142110 624746 142170 624822
rect 169017 624819 169083 624822
rect 294597 624819 294663 624822
rect 134934 624686 142170 624746
rect 57605 624610 57671 624613
rect 57605 624608 60076 624610
rect 57605 624552 57610 624608
rect 57666 624552 60076 624608
rect 57605 624550 60076 624552
rect 57605 624547 57671 624550
rect 177246 624548 177252 624612
rect 177316 624610 177322 624612
rect 177316 624550 180044 624610
rect 177316 624548 177322 624550
rect 297030 624548 297036 624612
rect 297100 624610 297106 624612
rect 374821 624610 374887 624613
rect 297100 624550 300196 624610
rect 374821 624608 374930 624610
rect 374821 624552 374826 624608
rect 374882 624552 374930 624608
rect 297100 624548 297106 624550
rect 374821 624547 374930 624552
rect 167637 624066 167703 624069
rect 294822 624066 294828 624068
rect 142110 624064 167703 624066
rect 134934 623930 134994 624036
rect 142110 624008 167642 624064
rect 167698 624008 167703 624064
rect 142110 624006 167703 624008
rect 254932 624006 294828 624066
rect 142110 623930 142170 624006
rect 167637 624003 167703 624006
rect 294822 624004 294828 624006
rect 294892 624004 294898 624068
rect 374870 624036 374930 624547
rect 550766 624066 550772 624068
rect 539948 624006 550772 624066
rect 550766 624004 550772 624006
rect 550836 624004 550842 624068
rect 134934 623870 142170 623930
rect 374453 623658 374519 623661
rect 374453 623656 374562 623658
rect 374453 623600 374458 623656
rect 374514 623600 374562 623656
rect 374453 623595 374562 623600
rect 57789 623522 57855 623525
rect 177573 623522 177639 623525
rect 297357 623522 297423 623525
rect 57789 623520 60076 623522
rect 57789 623464 57794 623520
rect 57850 623464 60076 623520
rect 57789 623462 60076 623464
rect 177573 623520 180044 623522
rect 177573 623464 177578 623520
rect 177634 623464 180044 623520
rect 177573 623462 180044 623464
rect 297357 623520 300196 623522
rect 297357 623464 297362 623520
rect 297418 623464 300196 623520
rect 297357 623462 300196 623464
rect 57789 623459 57855 623462
rect 177573 623459 177639 623462
rect 297357 623459 297423 623462
rect 166257 623250 166323 623253
rect 294638 623250 294644 623252
rect 142110 623248 166323 623250
rect 134934 623114 134994 623220
rect 142110 623192 166262 623248
rect 166318 623192 166323 623248
rect 142110 623190 166323 623192
rect 254932 623190 294644 623250
rect 142110 623114 142170 623190
rect 166257 623187 166323 623190
rect 294638 623188 294644 623190
rect 294708 623188 294714 623252
rect 374502 623220 374562 623595
rect 134934 623054 142170 623114
rect 134934 622510 142170 622570
rect 56961 622434 57027 622437
rect 56961 622432 60076 622434
rect 56961 622376 56966 622432
rect 57022 622376 60076 622432
rect 134934 622404 134994 622510
rect 142110 622434 142170 622510
rect 167821 622434 167887 622437
rect 142110 622432 167887 622434
rect 56961 622374 60076 622376
rect 142110 622376 167826 622432
rect 167882 622376 167887 622432
rect 142110 622374 167887 622376
rect 56961 622371 57027 622374
rect 167821 622371 167887 622374
rect 177614 622372 177620 622436
rect 177684 622434 177690 622436
rect 288382 622434 288388 622436
rect 177684 622374 180044 622434
rect 254932 622374 288388 622434
rect 177684 622372 177690 622374
rect 288382 622372 288388 622374
rect 288452 622372 288458 622436
rect 291929 622434 291995 622437
rect 377213 622434 377279 622437
rect 291929 622432 300196 622434
rect 291929 622376 291934 622432
rect 291990 622376 300196 622432
rect 291929 622374 300196 622376
rect 374900 622432 377279 622434
rect 374900 622376 377218 622432
rect 377274 622376 377279 622432
rect 374900 622374 377279 622376
rect 539918 622434 539978 622676
rect 540053 622434 540119 622437
rect 539918 622432 540119 622434
rect 539918 622376 540058 622432
rect 540114 622376 540119 622432
rect 539918 622374 540119 622376
rect 291929 622371 291995 622374
rect 377213 622371 377279 622374
rect 540053 622371 540119 622374
rect 178677 621618 178743 621621
rect 292062 621618 292068 621620
rect 142110 621616 178743 621618
rect 134934 621482 134994 621588
rect 142110 621560 178682 621616
rect 178738 621560 178743 621616
rect 142110 621558 178743 621560
rect 254932 621558 292068 621618
rect 142110 621482 142170 621558
rect 178677 621555 178743 621558
rect 292062 621556 292068 621558
rect 292132 621556 292138 621620
rect 375649 621618 375715 621621
rect 374900 621616 375715 621618
rect 374900 621560 375654 621616
rect 375710 621560 375715 621616
rect 374900 621558 375715 621560
rect 375649 621555 375715 621558
rect 134934 621422 142170 621482
rect 57237 621346 57303 621349
rect 57237 621344 60076 621346
rect 57237 621288 57242 621344
rect 57298 621288 60076 621344
rect 57237 621286 60076 621288
rect 57237 621283 57303 621286
rect 177062 621284 177068 621348
rect 177132 621346 177138 621348
rect 297357 621346 297423 621349
rect 543774 621346 543780 621348
rect 177132 621286 180044 621346
rect 297357 621344 300196 621346
rect 297357 621288 297362 621344
rect 297418 621288 300196 621344
rect 297357 621286 300196 621288
rect 539948 621286 543780 621346
rect 177132 621284 177138 621286
rect 297357 621283 297423 621286
rect 543774 621284 543780 621286
rect 543844 621284 543850 621348
rect 137277 620938 137343 620941
rect 134934 620936 137343 620938
rect 134934 620880 137282 620936
rect 137338 620880 137343 620936
rect 134934 620878 137343 620880
rect 134934 620772 134994 620878
rect 137277 620875 137343 620878
rect 294454 620802 294460 620804
rect 254932 620742 294460 620802
rect 294454 620740 294460 620742
rect 294524 620740 294530 620804
rect 376845 620802 376911 620805
rect 374900 620800 376911 620802
rect 374900 620744 376850 620800
rect 376906 620744 376911 620800
rect 374900 620742 376911 620744
rect 376845 620739 376911 620742
rect 59118 620196 59124 620260
rect 59188 620258 59194 620260
rect 59188 620198 60076 620258
rect 59188 620196 59194 620198
rect 177246 620196 177252 620260
rect 177316 620258 177322 620260
rect 298001 620258 298067 620261
rect 177316 620198 180044 620258
rect 298001 620256 300196 620258
rect 298001 620200 298006 620256
rect 298062 620200 300196 620256
rect 298001 620198 300196 620200
rect 177316 620196 177322 620198
rect 298001 620195 298067 620198
rect 171777 619986 171843 619989
rect 298134 619986 298140 619988
rect 142110 619984 171843 619986
rect 134934 619850 134994 619956
rect 142110 619928 171782 619984
rect 171838 619928 171843 619984
rect 142110 619926 171843 619928
rect 254932 619926 298140 619986
rect 142110 619850 142170 619926
rect 171777 619923 171843 619926
rect 298134 619924 298140 619926
rect 298204 619924 298210 619988
rect 378593 619986 378659 619989
rect 546534 619986 546540 619988
rect 374900 619984 378659 619986
rect 374900 619928 378598 619984
rect 378654 619928 378659 619984
rect 374900 619926 378659 619928
rect 539948 619926 546540 619986
rect 378593 619923 378659 619926
rect 546534 619924 546540 619926
rect 546604 619924 546610 619988
rect 134934 619790 142170 619850
rect -960 619170 480 619260
rect 29126 619170 29132 619172
rect -960 619110 29132 619170
rect -960 619020 480 619110
rect 29126 619108 29132 619110
rect 29196 619108 29202 619172
rect 58750 619108 58756 619172
rect 58820 619170 58826 619172
rect 58820 619110 60076 619170
rect 58820 619108 58826 619110
rect 134934 618626 134994 619140
rect 175038 619108 175044 619172
rect 175108 619170 175114 619172
rect 290590 619170 290596 619172
rect 175108 619110 180044 619170
rect 254932 619110 290596 619170
rect 175108 619108 175114 619110
rect 290590 619108 290596 619110
rect 290660 619108 290666 619172
rect 298001 619170 298067 619173
rect 376201 619170 376267 619173
rect 298001 619168 300196 619170
rect 298001 619112 298006 619168
rect 298062 619112 300196 619168
rect 298001 619110 300196 619112
rect 374900 619168 376267 619170
rect 374900 619112 376206 619168
rect 376262 619112 376267 619168
rect 374900 619110 376267 619112
rect 298001 619107 298067 619110
rect 376201 619107 376267 619110
rect 137461 618626 137527 618629
rect 550950 618626 550956 618628
rect 134934 618624 137527 618626
rect 134934 618568 137466 618624
rect 137522 618568 137527 618624
rect 134934 618566 137527 618568
rect 539948 618566 550956 618626
rect 137461 618563 137527 618566
rect 550950 618564 550956 618566
rect 551020 618564 551026 618628
rect 374637 618490 374703 618493
rect 134934 618430 142170 618490
rect 134934 618324 134994 618430
rect 142110 618354 142170 618430
rect 374637 618488 374746 618490
rect 374637 618432 374642 618488
rect 374698 618432 374746 618488
rect 374637 618427 374746 618432
rect 172646 618354 172652 618356
rect 142110 618294 172652 618354
rect 172646 618292 172652 618294
rect 172716 618292 172722 618356
rect 295374 618354 295380 618356
rect 254932 618294 295380 618354
rect 295374 618292 295380 618294
rect 295444 618292 295450 618356
rect 374686 618324 374746 618427
rect 58801 618082 58867 618085
rect 58801 618080 60076 618082
rect 58801 618024 58806 618080
rect 58862 618024 60076 618080
rect 58801 618022 60076 618024
rect 58801 618019 58867 618022
rect 177430 618020 177436 618084
rect 177500 618082 177506 618084
rect 298001 618082 298067 618085
rect 177500 618022 180044 618082
rect 298001 618080 300196 618082
rect 298001 618024 298006 618080
rect 298062 618024 300196 618080
rect 298001 618022 300196 618024
rect 177500 618020 177506 618022
rect 298001 618019 298067 618022
rect 175222 617538 175228 617540
rect 134934 617402 134994 617508
rect 142110 617478 175228 617538
rect 142110 617402 142170 617478
rect 175222 617476 175228 617478
rect 175292 617476 175298 617540
rect 287094 617538 287100 617540
rect 254932 617478 287100 617538
rect 287094 617476 287100 617478
rect 287164 617476 287170 617540
rect 375741 617538 375807 617541
rect 374900 617536 375807 617538
rect 374900 617480 375746 617536
rect 375802 617480 375807 617536
rect 374900 617478 375807 617480
rect 375741 617475 375807 617478
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 134934 617342 142170 617402
rect 583520 617388 584960 617478
rect 542905 617266 542971 617269
rect 539948 617264 542971 617266
rect 539948 617208 542910 617264
rect 542966 617208 542971 617264
rect 539948 617206 542971 617208
rect 542905 617203 542971 617206
rect 58985 616994 59051 616997
rect 58985 616992 60076 616994
rect 58985 616936 58990 616992
rect 59046 616936 60076 616992
rect 58985 616934 60076 616936
rect 58985 616931 59051 616934
rect 176326 616932 176332 616996
rect 176396 616994 176402 616996
rect 297449 616994 297515 616997
rect 176396 616934 180044 616994
rect 297449 616992 300196 616994
rect 297449 616936 297454 616992
rect 297510 616936 300196 616992
rect 297449 616934 300196 616936
rect 176396 616932 176402 616934
rect 297449 616931 297515 616934
rect 173934 616722 173940 616724
rect 134934 616586 134994 616692
rect 142110 616662 173940 616722
rect 142110 616586 142170 616662
rect 173934 616660 173940 616662
rect 174004 616660 174010 616724
rect 295926 616722 295932 616724
rect 254932 616662 295932 616722
rect 295926 616660 295932 616662
rect 295996 616660 296002 616724
rect 378317 616722 378383 616725
rect 374900 616720 378383 616722
rect 374900 616664 378322 616720
rect 378378 616664 378383 616720
rect 374900 616662 378383 616664
rect 378317 616659 378383 616662
rect 134934 616526 142170 616586
rect 58249 615906 58315 615909
rect 173249 615906 173315 615909
rect 58249 615904 60076 615906
rect 58249 615848 58254 615904
rect 58310 615848 60076 615904
rect 142110 615904 173315 615906
rect 58249 615846 60076 615848
rect 58249 615843 58315 615846
rect 134934 615770 134994 615876
rect 142110 615848 173254 615904
rect 173310 615848 173315 615904
rect 142110 615846 173315 615848
rect 142110 615770 142170 615846
rect 173249 615843 173315 615846
rect 176510 615844 176516 615908
rect 176580 615906 176586 615908
rect 282126 615906 282132 615908
rect 176580 615846 180044 615906
rect 254932 615846 282132 615906
rect 176580 615844 176586 615846
rect 282126 615844 282132 615846
rect 282196 615844 282202 615908
rect 291878 615844 291884 615908
rect 291948 615906 291954 615908
rect 376293 615906 376359 615909
rect 542905 615906 542971 615909
rect 291948 615846 300196 615906
rect 374900 615904 376359 615906
rect 374900 615848 376298 615904
rect 376354 615848 376359 615904
rect 374900 615846 376359 615848
rect 539948 615904 542971 615906
rect 539948 615848 542910 615904
rect 542966 615848 542971 615904
rect 539948 615846 542971 615848
rect 291948 615844 291954 615846
rect 376293 615843 376359 615846
rect 542905 615843 542971 615846
rect 134934 615710 142170 615770
rect 134934 615166 142170 615226
rect 134934 615060 134994 615166
rect 142110 615090 142170 615166
rect 171869 615090 171935 615093
rect 288566 615090 288572 615092
rect 142110 615088 171935 615090
rect 142110 615032 171874 615088
rect 171930 615032 171935 615088
rect 142110 615030 171935 615032
rect 254932 615030 288572 615090
rect 171869 615027 171935 615030
rect 288566 615028 288572 615030
rect 288636 615028 288642 615092
rect 377806 615090 377812 615092
rect 374900 615030 377812 615090
rect 377806 615028 377812 615030
rect 377876 615028 377882 615092
rect 58433 614818 58499 614821
rect 58433 614816 60076 614818
rect 58433 614760 58438 614816
rect 58494 614760 60076 614816
rect 58433 614758 60076 614760
rect 58433 614755 58499 614758
rect 177798 614756 177804 614820
rect 177868 614818 177874 614820
rect 177868 614758 180044 614818
rect 177868 614756 177874 614758
rect 291694 614756 291700 614820
rect 291764 614818 291770 614820
rect 291764 614758 300196 614818
rect 291764 614756 291770 614758
rect 541014 614546 541020 614548
rect 539948 614486 541020 614546
rect 541014 614484 541020 614486
rect 541084 614484 541090 614548
rect 134934 614350 142170 614410
rect 134934 614244 134994 614350
rect 142110 614274 142170 614350
rect 173433 614274 173499 614277
rect 294822 614274 294828 614276
rect 142110 614272 173499 614274
rect 142110 614216 173438 614272
rect 173494 614216 173499 614272
rect 142110 614214 173499 614216
rect 254932 614214 294828 614274
rect 173433 614211 173499 614214
rect 294822 614212 294828 614214
rect 294892 614212 294898 614276
rect 374502 614005 374562 614244
rect 374502 614000 374611 614005
rect 374502 613944 374550 614000
rect 374606 613944 374611 614000
rect 374502 613942 374611 613944
rect 374545 613939 374611 613942
rect 58893 613730 58959 613733
rect 58893 613728 60076 613730
rect 58893 613672 58898 613728
rect 58954 613672 60076 613728
rect 58893 613670 60076 613672
rect 58893 613667 58959 613670
rect 177430 613668 177436 613732
rect 177500 613730 177506 613732
rect 298001 613730 298067 613733
rect 177500 613670 180044 613730
rect 298001 613728 300196 613730
rect 298001 613672 298006 613728
rect 298062 613672 300196 613728
rect 298001 613670 300196 613672
rect 177500 613668 177506 613670
rect 298001 613667 298067 613670
rect 134934 613534 142170 613594
rect 134934 613428 134994 613534
rect 142110 613458 142170 613534
rect 174629 613458 174695 613461
rect 280654 613458 280660 613460
rect 142110 613456 174695 613458
rect 142110 613400 174634 613456
rect 174690 613400 174695 613456
rect 142110 613398 174695 613400
rect 254932 613398 280660 613458
rect 174629 613395 174695 613398
rect 280654 613396 280660 613398
rect 280724 613396 280730 613460
rect 375833 613458 375899 613461
rect 374900 613456 375899 613458
rect 374900 613400 375838 613456
rect 375894 613400 375899 613456
rect 374900 613398 375899 613400
rect 375833 613395 375899 613398
rect 392577 613322 392643 613325
rect 397545 613322 397611 613325
rect 392577 613320 397611 613322
rect 392577 613264 392582 613320
rect 392638 613264 397550 613320
rect 397606 613264 397611 613320
rect 392577 613262 397611 613264
rect 392577 613259 392643 613262
rect 397545 613259 397611 613262
rect 480897 613322 480963 613325
rect 487061 613322 487127 613325
rect 490054 613322 490114 613700
rect 480897 613320 490114 613322
rect 480897 613264 480902 613320
rect 480958 613264 487066 613320
rect 487122 613264 490114 613320
rect 480897 613262 490114 613264
rect 480897 613259 480963 613262
rect 487061 613259 487127 613262
rect 542854 613186 542860 613188
rect 539948 613126 542860 613186
rect 542854 613124 542860 613126
rect 542924 613124 542930 613188
rect 56133 612642 56199 612645
rect 173157 612642 173223 612645
rect 56133 612640 60076 612642
rect 56133 612584 56138 612640
rect 56194 612584 60076 612640
rect 142110 612640 173223 612642
rect 56133 612582 60076 612584
rect 56133 612579 56199 612582
rect 134934 612506 134994 612612
rect 142110 612584 173162 612640
rect 173218 612584 173223 612640
rect 142110 612582 173223 612584
rect 142110 612506 142170 612582
rect 173157 612579 173223 612582
rect 177062 612580 177068 612644
rect 177132 612642 177138 612644
rect 294454 612642 294460 612644
rect 177132 612582 180044 612642
rect 254932 612582 294460 612642
rect 177132 612580 177138 612582
rect 294454 612580 294460 612582
rect 294524 612580 294530 612644
rect 298001 612642 298067 612645
rect 298001 612640 300196 612642
rect 298001 612584 298006 612640
rect 298062 612584 300196 612640
rect 298001 612582 300196 612584
rect 298001 612579 298067 612582
rect 134934 612446 142170 612506
rect 374502 612101 374562 612612
rect 374453 612096 374562 612101
rect 374453 612040 374458 612096
rect 374514 612040 374562 612096
rect 374453 612038 374562 612040
rect 374453 612035 374519 612038
rect 284886 611826 284892 611828
rect 57329 611554 57395 611557
rect 57329 611552 60076 611554
rect 57329 611496 57334 611552
rect 57390 611496 60076 611552
rect 57329 611494 60076 611496
rect 57329 611491 57395 611494
rect 134934 611418 134994 611796
rect 254932 611766 284892 611826
rect 284886 611764 284892 611766
rect 284956 611764 284962 611828
rect 378409 611826 378475 611829
rect 541198 611826 541204 611828
rect 374900 611824 378475 611826
rect 374900 611768 378414 611824
rect 378470 611768 378475 611824
rect 374900 611766 378475 611768
rect 539948 611766 541204 611826
rect 378409 611763 378475 611766
rect 541198 611764 541204 611766
rect 541268 611764 541274 611828
rect 177798 611492 177804 611556
rect 177868 611554 177874 611556
rect 284201 611554 284267 611557
rect 177868 611494 180044 611554
rect 284201 611552 300196 611554
rect 284201 611496 284206 611552
rect 284262 611496 300196 611552
rect 284201 611494 300196 611496
rect 177868 611492 177874 611494
rect 284201 611491 284267 611494
rect 137277 611418 137343 611421
rect 134934 611416 137343 611418
rect 134934 611360 137282 611416
rect 137338 611360 137343 611416
rect 134934 611358 137343 611360
rect 137277 611355 137343 611358
rect 177021 611418 177087 611421
rect 177614 611418 177620 611420
rect 177021 611416 177620 611418
rect 177021 611360 177026 611416
rect 177082 611360 177620 611416
rect 177021 611358 177620 611360
rect 177021 611355 177087 611358
rect 177614 611356 177620 611358
rect 177684 611356 177690 611420
rect 134934 611086 142170 611146
rect 134934 610980 134994 611086
rect 142110 611010 142170 611086
rect 174537 611010 174603 611013
rect 256734 611010 256740 611012
rect 142110 611008 174603 611010
rect 142110 610952 174542 611008
rect 174598 610952 174603 611008
rect 142110 610950 174603 610952
rect 254932 610950 256740 611010
rect 174537 610947 174603 610950
rect 256734 610948 256740 610950
rect 256804 610948 256810 611012
rect 375649 611010 375715 611013
rect 374900 611008 375715 611010
rect 374900 610952 375654 611008
rect 375710 610952 375715 611008
rect 374900 610950 375715 610952
rect 375649 610947 375715 610950
rect 177246 610676 177252 610740
rect 177316 610738 177322 610740
rect 177849 610738 177915 610741
rect 177316 610736 177915 610738
rect 177316 610680 177854 610736
rect 177910 610680 177915 610736
rect 177316 610678 177915 610680
rect 177316 610676 177322 610678
rect 177849 610675 177915 610678
rect 59670 610404 59676 610468
rect 59740 610466 59746 610468
rect 59740 610406 60076 610466
rect 59740 610404 59746 610406
rect 177982 610404 177988 610468
rect 178052 610466 178058 610468
rect 178052 610406 180044 610466
rect 178052 610404 178058 610406
rect 286174 610404 286180 610468
rect 286244 610466 286250 610468
rect 543406 610466 543412 610468
rect 286244 610406 300196 610466
rect 539948 610406 543412 610466
rect 286244 610404 286250 610406
rect 543406 610404 543412 610406
rect 543476 610404 543482 610468
rect 134934 610270 142170 610330
rect 134934 610164 134994 610270
rect 142110 610194 142170 610270
rect 175917 610194 175983 610197
rect 298318 610194 298324 610196
rect 142110 610192 175983 610194
rect 142110 610136 175922 610192
rect 175978 610136 175983 610192
rect 142110 610134 175983 610136
rect 254932 610134 298324 610194
rect 175917 610131 175983 610134
rect 298318 610132 298324 610134
rect 298388 610132 298394 610196
rect 378501 610194 378567 610197
rect 374900 610192 378567 610194
rect 374900 610136 378506 610192
rect 378562 610136 378567 610192
rect 374900 610134 378567 610136
rect 378501 610131 378567 610134
rect 177297 609786 177363 609789
rect 177430 609786 177436 609788
rect 177297 609784 177436 609786
rect 177297 609728 177302 609784
rect 177358 609728 177436 609784
rect 177297 609726 177436 609728
rect 177297 609723 177363 609726
rect 177430 609724 177436 609726
rect 177500 609724 177506 609788
rect 57421 609378 57487 609381
rect 57421 609376 60076 609378
rect 57421 609320 57426 609376
rect 57482 609320 60076 609376
rect 57421 609318 60076 609320
rect 57421 609315 57487 609318
rect 134934 609106 134994 609348
rect 176694 609316 176700 609380
rect 176764 609378 176770 609380
rect 294638 609378 294644 609380
rect 176764 609318 180044 609378
rect 254932 609318 294644 609378
rect 176764 609316 176770 609318
rect 294638 609316 294644 609318
rect 294708 609316 294714 609380
rect 297541 609378 297607 609381
rect 378869 609378 378935 609381
rect 297541 609376 300196 609378
rect 297541 609320 297546 609376
rect 297602 609320 300196 609376
rect 297541 609318 300196 609320
rect 374900 609376 378935 609378
rect 374900 609320 378874 609376
rect 378930 609320 378935 609376
rect 374900 609318 378935 609320
rect 297541 609315 297607 609318
rect 378869 609315 378935 609318
rect 178166 609106 178172 609108
rect 134934 609046 178172 609106
rect 178166 609044 178172 609046
rect 178236 609044 178242 609108
rect 539366 608701 539426 609076
rect 539366 608696 539475 608701
rect 539366 608640 539414 608696
rect 539470 608640 539475 608696
rect 539366 608638 539475 608640
rect 539409 608635 539475 608638
rect 177389 608562 177455 608565
rect 177798 608562 177804 608564
rect 177389 608560 177804 608562
rect 59721 608290 59787 608293
rect 59721 608288 60076 608290
rect 59721 608232 59726 608288
rect 59782 608232 60076 608288
rect 59721 608230 60076 608232
rect 59721 608227 59787 608230
rect 134934 608018 134994 608532
rect 177389 608504 177394 608560
rect 177450 608504 177804 608560
rect 177389 608502 177804 608504
rect 177389 608499 177455 608502
rect 177798 608500 177804 608502
rect 177868 608500 177874 608564
rect 290774 608562 290780 608564
rect 254932 608502 290780 608562
rect 290774 608500 290780 608502
rect 290844 608500 290850 608564
rect 375557 608562 375623 608565
rect 374900 608560 375623 608562
rect 374900 608504 375562 608560
rect 375618 608504 375623 608560
rect 374900 608502 375623 608504
rect 375557 608499 375623 608502
rect 177246 608228 177252 608292
rect 177316 608290 177322 608292
rect 297449 608290 297515 608293
rect 177316 608230 180044 608290
rect 297449 608288 300196 608290
rect 297449 608232 297454 608288
rect 297510 608232 300196 608288
rect 297449 608230 300196 608232
rect 177316 608228 177322 608230
rect 297449 608227 297515 608230
rect 137645 608018 137711 608021
rect 134934 608016 137711 608018
rect 134934 607960 137650 608016
rect 137706 607960 137711 608016
rect 134934 607958 137711 607960
rect 137645 607955 137711 607958
rect 134934 607822 142170 607882
rect 134934 607716 134994 607822
rect 142110 607746 142170 607822
rect 164877 607746 164943 607749
rect 299606 607746 299612 607748
rect 142110 607744 164943 607746
rect 142110 607688 164882 607744
rect 164938 607688 164943 607744
rect 142110 607686 164943 607688
rect 254932 607686 299612 607746
rect 164877 607683 164943 607686
rect 299606 607684 299612 607686
rect 299676 607684 299682 607748
rect 543038 607746 543044 607748
rect 374870 607341 374930 607716
rect 539948 607686 543044 607746
rect 543038 607684 543044 607686
rect 543108 607684 543114 607748
rect 374821 607336 374930 607341
rect 374821 607280 374826 607336
rect 374882 607280 374930 607336
rect 374821 607278 374930 607280
rect 374821 607275 374887 607278
rect 58709 607202 58775 607205
rect 58709 607200 60076 607202
rect 58709 607144 58714 607200
rect 58770 607144 60076 607200
rect 58709 607142 60076 607144
rect 58709 607139 58775 607142
rect 177062 607140 177068 607204
rect 177132 607202 177138 607204
rect 177205 607202 177271 607205
rect 177132 607200 177271 607202
rect 177132 607144 177210 607200
rect 177266 607144 177271 607200
rect 177132 607142 177271 607144
rect 177132 607140 177138 607142
rect 177205 607139 177271 607142
rect 177798 607140 177804 607204
rect 177868 607202 177874 607204
rect 177868 607142 180044 607202
rect 177868 607140 177874 607142
rect 296662 607140 296668 607204
rect 296732 607202 296738 607204
rect 397545 607202 397611 607205
rect 400949 607202 401015 607205
rect 296732 607142 300196 607202
rect 397545 607200 401015 607202
rect 397545 607144 397550 607200
rect 397606 607144 400954 607200
rect 401010 607144 401015 607200
rect 397545 607142 401015 607144
rect 296732 607140 296738 607142
rect 397545 607139 397611 607142
rect 400949 607139 401015 607142
rect 177665 607066 177731 607069
rect 177982 607066 177988 607068
rect 177665 607064 177988 607066
rect 177665 607008 177670 607064
rect 177726 607008 177988 607064
rect 177665 607006 177988 607008
rect 177665 607003 177731 607006
rect 177982 607004 177988 607006
rect 178052 607004 178058 607068
rect 298502 606930 298508 606932
rect 134934 606386 134994 606900
rect 254932 606870 298508 606930
rect 298502 606868 298508 606870
rect 298572 606868 298578 606932
rect 375465 606930 375531 606933
rect 374900 606928 375531 606930
rect 374900 606872 375470 606928
rect 375526 606872 375531 606928
rect 374900 606870 375531 606872
rect 375465 606867 375531 606870
rect 137369 606386 137435 606389
rect 543222 606386 543228 606388
rect 134934 606384 137435 606386
rect 134934 606328 137374 606384
rect 137430 606328 137435 606384
rect 134934 606326 137435 606328
rect 539948 606326 543228 606386
rect 137369 606323 137435 606326
rect 543222 606324 543228 606326
rect 543292 606324 543298 606388
rect -960 606114 480 606204
rect 134934 606190 142170 606250
rect 26734 606114 26740 606116
rect -960 606054 26740 606114
rect -960 605964 480 606054
rect 26734 606052 26740 606054
rect 26804 606052 26810 606116
rect 59813 606114 59879 606117
rect 59813 606112 60076 606114
rect 59813 606056 59818 606112
rect 59874 606056 60076 606112
rect 134934 606084 134994 606190
rect 142110 606114 142170 606190
rect 176009 606114 176075 606117
rect 142110 606112 176075 606114
rect 59813 606054 60076 606056
rect 142110 606056 176014 606112
rect 176070 606056 176075 606112
rect 142110 606054 176075 606056
rect 59813 606051 59879 606054
rect 176009 606051 176075 606054
rect 177062 606052 177068 606116
rect 177132 606114 177138 606116
rect 292614 606114 292620 606116
rect 177132 606054 180044 606114
rect 254932 606054 292620 606114
rect 177132 606052 177138 606054
rect 292614 606052 292620 606054
rect 292684 606052 292690 606116
rect 297633 606114 297699 606117
rect 378041 606114 378107 606117
rect 297633 606112 300196 606114
rect 297633 606056 297638 606112
rect 297694 606056 300196 606112
rect 297633 606054 300196 606056
rect 374900 606112 378107 606114
rect 374900 606056 378046 606112
rect 378102 606056 378107 606112
rect 374900 606054 378107 606056
rect 297633 606051 297699 606054
rect 378041 606051 378107 606054
rect 166441 605298 166507 605301
rect 299422 605298 299428 605300
rect 142110 605296 166507 605298
rect 134934 605162 134994 605268
rect 142110 605240 166446 605296
rect 166502 605240 166507 605296
rect 142110 605238 166507 605240
rect 254932 605238 299428 605298
rect 142110 605162 142170 605238
rect 166441 605235 166507 605238
rect 299422 605236 299428 605238
rect 299492 605236 299498 605300
rect 377029 605298 377095 605301
rect 374900 605296 377095 605298
rect 374900 605240 377034 605296
rect 377090 605240 377095 605296
rect 374900 605238 377095 605240
rect 377029 605235 377095 605238
rect 134934 605102 142170 605162
rect 57053 605026 57119 605029
rect 57053 605024 60076 605026
rect 57053 604968 57058 605024
rect 57114 604968 60076 605024
rect 57053 604966 60076 604968
rect 57053 604963 57119 604966
rect 177614 604964 177620 605028
rect 177684 605026 177690 605028
rect 177684 604966 180044 605026
rect 177684 604964 177690 604966
rect 297030 604964 297036 605028
rect 297100 605026 297106 605028
rect 297100 604966 300196 605026
rect 297100 604964 297106 604966
rect 539358 604964 539364 605028
rect 539428 604964 539434 605028
rect 134934 604558 135178 604618
rect 134934 604452 134994 604558
rect 135118 604482 135178 604558
rect 137553 604482 137619 604485
rect 135118 604480 137619 604482
rect 135118 604424 137558 604480
rect 137614 604424 137619 604480
rect 135118 604422 137619 604424
rect 137553 604419 137619 604422
rect 176694 604420 176700 604484
rect 176764 604482 176770 604484
rect 177757 604482 177823 604485
rect 299238 604482 299244 604484
rect 176764 604480 177823 604482
rect 176764 604424 177762 604480
rect 177818 604424 177823 604480
rect 176764 604422 177823 604424
rect 254932 604422 299244 604482
rect 176764 604420 176770 604422
rect 177757 604419 177823 604422
rect 299238 604420 299244 604422
rect 299308 604420 299314 604484
rect 299606 604420 299612 604484
rect 299676 604482 299682 604484
rect 299841 604482 299907 604485
rect 378041 604482 378107 604485
rect 299676 604480 299907 604482
rect 299676 604424 299846 604480
rect 299902 604424 299907 604480
rect 299676 604422 299907 604424
rect 374900 604480 378107 604482
rect 374900 604424 378046 604480
rect 378102 604424 378107 604480
rect 374900 604422 378107 604424
rect 299676 604420 299682 604422
rect 299841 604419 299907 604422
rect 378041 604419 378107 604422
rect 583520 604060 584960 604300
rect 58065 603938 58131 603941
rect 58065 603936 60076 603938
rect 58065 603880 58070 603936
rect 58126 603880 60076 603936
rect 58065 603878 60076 603880
rect 58065 603875 58131 603878
rect 166758 603876 166764 603940
rect 166828 603938 166834 603940
rect 297909 603938 297975 603941
rect 166828 603878 180044 603938
rect 297909 603936 300196 603938
rect 297909 603880 297914 603936
rect 297970 603880 300196 603936
rect 297909 603878 300196 603880
rect 166828 603876 166834 603878
rect 297909 603875 297975 603878
rect 163589 603666 163655 603669
rect 287646 603666 287652 603668
rect 142110 603664 163655 603666
rect 134934 603530 134994 603636
rect 142110 603608 163594 603664
rect 163650 603608 163655 603664
rect 142110 603606 163655 603608
rect 254932 603606 287652 603666
rect 142110 603530 142170 603606
rect 163589 603603 163655 603606
rect 287646 603604 287652 603606
rect 287716 603604 287722 603668
rect 375557 603666 375623 603669
rect 374900 603664 375623 603666
rect 374900 603608 375562 603664
rect 375618 603608 375623 603664
rect 374900 603606 375623 603608
rect 375557 603603 375623 603606
rect 539542 603604 539548 603668
rect 539612 603604 539618 603668
rect 134934 603470 142170 603530
rect 298686 602986 298692 602988
rect 296670 602926 298692 602986
rect 59813 602850 59879 602853
rect 173341 602850 173407 602853
rect 59813 602848 60076 602850
rect 59813 602792 59818 602848
rect 59874 602792 60076 602848
rect 142110 602848 173407 602850
rect 59813 602790 60076 602792
rect 59813 602787 59879 602790
rect 134934 602714 134994 602820
rect 142110 602792 173346 602848
rect 173402 602792 173407 602848
rect 142110 602790 173407 602792
rect 142110 602714 142170 602790
rect 173341 602787 173407 602790
rect 177430 602788 177436 602852
rect 177500 602850 177506 602852
rect 296670 602850 296730 602926
rect 298686 602924 298692 602926
rect 298756 602924 298762 602988
rect 299422 602924 299428 602988
rect 299492 602986 299498 602988
rect 299749 602986 299815 602989
rect 299492 602984 299815 602986
rect 299492 602928 299754 602984
rect 299810 602928 299815 602984
rect 299492 602926 299815 602928
rect 299492 602924 299498 602926
rect 299749 602923 299815 602926
rect 375373 602850 375439 602853
rect 177500 602790 180044 602850
rect 254932 602790 296730 602850
rect 298326 602790 300196 602850
rect 374900 602848 375439 602850
rect 374900 602792 375378 602848
rect 375434 602792 375439 602848
rect 374900 602790 375439 602792
rect 177500 602788 177506 602790
rect 134934 602654 142170 602714
rect 255262 602516 255268 602580
rect 255332 602578 255338 602580
rect 298326 602578 298386 602790
rect 375373 602787 375439 602790
rect 255332 602518 298386 602578
rect 255332 602516 255338 602518
rect 171961 602034 172027 602037
rect 299422 602034 299428 602036
rect 142110 602032 172027 602034
rect 134934 601898 134994 602004
rect 142110 601976 171966 602032
rect 172022 601976 172027 602032
rect 142110 601974 172027 601976
rect 254932 601974 299428 602034
rect 142110 601898 142170 601974
rect 171961 601971 172027 601974
rect 299422 601972 299428 601974
rect 299492 601972 299498 602036
rect 375925 602034 375991 602037
rect 374900 602032 375991 602034
rect 374900 601976 375930 602032
rect 375986 601976 375991 602032
rect 374900 601974 375991 601976
rect 375925 601971 375991 601974
rect 134934 601838 142170 601898
rect 298134 601836 298140 601900
rect 298204 601898 298210 601900
rect 299381 601898 299447 601901
rect 298204 601896 299447 601898
rect 298204 601840 299386 601896
rect 299442 601840 299447 601896
rect 298204 601838 299447 601840
rect 298204 601836 298210 601838
rect 299381 601835 299447 601838
rect 58525 601762 58591 601765
rect 58525 601760 60076 601762
rect 58525 601704 58530 601760
rect 58586 601704 60076 601760
rect 58525 601702 60076 601704
rect 58525 601699 58591 601702
rect 177246 601700 177252 601764
rect 177316 601762 177322 601764
rect 177481 601762 177547 601765
rect 177316 601760 177547 601762
rect 177316 601704 177486 601760
rect 177542 601704 177547 601760
rect 177316 601702 177547 601704
rect 177316 601700 177322 601702
rect 177481 601699 177547 601702
rect 179045 601762 179111 601765
rect 260189 601762 260255 601765
rect 179045 601760 180044 601762
rect 179045 601704 179050 601760
rect 179106 601704 180044 601760
rect 179045 601702 180044 601704
rect 260189 601760 300196 601762
rect 260189 601704 260194 601760
rect 260250 601704 300196 601760
rect 260189 601702 300196 601704
rect 179045 601699 179111 601702
rect 260189 601699 260255 601702
rect 538254 601700 538260 601764
rect 538324 601762 538330 601764
rect 539409 601762 539475 601765
rect 538324 601760 539475 601762
rect 538324 601704 539414 601760
rect 539470 601704 539475 601760
rect 538324 601702 539475 601704
rect 538324 601700 538330 601702
rect 539409 601699 539475 601702
rect 172053 601218 172119 601221
rect 295006 601218 295012 601220
rect 142110 601216 172119 601218
rect 134934 601082 134994 601188
rect 142110 601160 172058 601216
rect 172114 601160 172119 601216
rect 142110 601158 172119 601160
rect 254932 601158 295012 601218
rect 142110 601082 142170 601158
rect 172053 601155 172119 601158
rect 295006 601156 295012 601158
rect 295076 601156 295082 601220
rect 378685 601218 378751 601221
rect 374900 601216 378751 601218
rect 374900 601160 378690 601216
rect 378746 601160 378751 601216
rect 374900 601158 378751 601160
rect 378685 601155 378751 601158
rect 134934 601022 142170 601082
rect 294822 601020 294828 601084
rect 294892 601082 294898 601084
rect 295241 601082 295307 601085
rect 294892 601080 295307 601082
rect 294892 601024 295246 601080
rect 295302 601024 295307 601080
rect 294892 601022 295307 601024
rect 294892 601020 294898 601022
rect 295241 601019 295307 601022
rect 539501 601082 539567 601085
rect 545113 601082 545179 601085
rect 539501 601080 545179 601082
rect 539501 601024 539506 601080
rect 539562 601024 545118 601080
rect 545174 601024 545179 601080
rect 539501 601022 545179 601024
rect 539501 601019 539567 601022
rect 545113 601019 545179 601022
rect 57697 600674 57763 600677
rect 178953 600674 179019 600677
rect 260281 600674 260347 600677
rect 57697 600672 60076 600674
rect 57697 600616 57702 600672
rect 57758 600616 60076 600672
rect 57697 600614 60076 600616
rect 178953 600672 180044 600674
rect 178953 600616 178958 600672
rect 179014 600616 180044 600672
rect 178953 600614 180044 600616
rect 260281 600672 300196 600674
rect 260281 600616 260286 600672
rect 260342 600616 300196 600672
rect 260281 600614 300196 600616
rect 57697 600611 57763 600614
rect 178953 600611 179019 600614
rect 260281 600611 260347 600614
rect 537293 600538 537359 600541
rect 541065 600538 541131 600541
rect 134934 600478 142170 600538
rect 134934 600372 134994 600478
rect 142110 600402 142170 600478
rect 537293 600536 541131 600538
rect 537293 600480 537298 600536
rect 537354 600480 541070 600536
rect 541126 600480 541131 600536
rect 537293 600478 541131 600480
rect 537293 600475 537359 600478
rect 541065 600475 541131 600478
rect 170489 600402 170555 600405
rect 295742 600402 295748 600404
rect 142110 600400 170555 600402
rect 142110 600344 170494 600400
rect 170550 600344 170555 600400
rect 142110 600342 170555 600344
rect 254932 600342 295748 600402
rect 170489 600339 170555 600342
rect 295742 600340 295748 600342
rect 295812 600340 295818 600404
rect 376753 600402 376819 600405
rect 374900 600400 376819 600402
rect 374900 600344 376758 600400
rect 376814 600344 376819 600400
rect 374900 600342 376819 600344
rect 376753 600339 376819 600342
rect 538806 600340 538812 600404
rect 538876 600402 538882 600404
rect 539542 600402 539548 600404
rect 538876 600342 539548 600402
rect 538876 600340 538882 600342
rect 539542 600340 539548 600342
rect 539612 600340 539618 600404
rect 255957 600266 256023 600269
rect 255957 600264 258090 600266
rect 255957 600208 255962 600264
rect 256018 600208 258090 600264
rect 255957 600206 258090 600208
rect 255957 600203 256023 600206
rect 54569 599586 54635 599589
rect 170581 599586 170647 599589
rect 54569 599584 60076 599586
rect 54569 599528 54574 599584
rect 54630 599528 60076 599584
rect 142110 599584 170647 599586
rect 54569 599526 60076 599528
rect 54569 599523 54635 599526
rect 134934 599450 134994 599556
rect 142110 599528 170586 599584
rect 170642 599528 170647 599584
rect 142110 599526 170647 599528
rect 142110 599450 142170 599526
rect 170581 599523 170647 599526
rect 179137 599586 179203 599589
rect 258030 599586 258090 600206
rect 488073 600130 488139 600133
rect 504817 600130 504883 600133
rect 488073 600128 504883 600130
rect 488073 600072 488078 600128
rect 488134 600072 504822 600128
rect 504878 600072 504883 600128
rect 488073 600070 504883 600072
rect 488073 600067 488139 600070
rect 504817 600067 504883 600070
rect 489821 599994 489887 599997
rect 528737 599994 528803 599997
rect 489821 599992 528803 599994
rect 489821 599936 489826 599992
rect 489882 599936 528742 599992
rect 528798 599936 528803 599992
rect 489821 599934 528803 599936
rect 489821 599931 489887 599934
rect 528737 599931 528803 599934
rect 488165 599858 488231 599861
rect 532877 599858 532943 599861
rect 488165 599856 532943 599858
rect 488165 599800 488170 599856
rect 488226 599800 532882 599856
rect 532938 599800 532943 599856
rect 488165 599798 532943 599800
rect 488165 599795 488231 599798
rect 532877 599795 532943 599798
rect 397453 599722 397519 599725
rect 500166 599722 500172 599724
rect 397453 599720 500172 599722
rect 397453 599664 397458 599720
rect 397514 599664 500172 599720
rect 397453 599662 500172 599664
rect 397453 599659 397519 599662
rect 500166 599660 500172 599662
rect 500236 599660 500242 599724
rect 258165 599586 258231 599589
rect 386505 599586 386571 599589
rect 179137 599584 180044 599586
rect 179137 599528 179142 599584
rect 179198 599528 180044 599584
rect 258030 599584 300196 599586
rect 179137 599526 180044 599528
rect 179137 599523 179203 599526
rect 134934 599390 142170 599450
rect 254902 599450 254962 599556
rect 258030 599528 258170 599584
rect 258226 599528 300196 599584
rect 258030 599526 300196 599528
rect 374900 599584 386571 599586
rect 374900 599528 386510 599584
rect 386566 599528 386571 599584
rect 374900 599526 386571 599528
rect 258165 599523 258231 599526
rect 386505 599523 386571 599526
rect 487061 599586 487127 599589
rect 505093 599586 505159 599589
rect 487061 599584 505159 599586
rect 487061 599528 487066 599584
rect 487122 599528 505098 599584
rect 505154 599528 505159 599584
rect 487061 599526 505159 599528
rect 487061 599523 487127 599526
rect 505093 599523 505159 599526
rect 296294 599450 296300 599452
rect 254902 599390 296300 599450
rect 296294 599388 296300 599390
rect 296364 599388 296370 599452
rect 256734 598844 256740 598908
rect 256804 598906 256810 598908
rect 257981 598906 258047 598909
rect 256804 598904 258047 598906
rect 256804 598848 257986 598904
rect 258042 598848 258047 598904
rect 256804 598846 258047 598848
rect 256804 598844 256810 598846
rect 257981 598843 258047 598846
rect 503161 598906 503227 598909
rect 535453 598906 535519 598909
rect 503161 598904 535519 598906
rect 503161 598848 503166 598904
rect 503222 598848 535458 598904
rect 535514 598848 535519 598904
rect 503161 598846 535519 598848
rect 503161 598843 503227 598846
rect 535453 598843 535519 598846
rect 170397 598770 170463 598773
rect 256918 598770 256924 598772
rect 142110 598768 170463 598770
rect 134934 598634 134994 598740
rect 142110 598712 170402 598768
rect 170458 598712 170463 598768
rect 142110 598710 170463 598712
rect 254932 598710 256924 598770
rect 142110 598634 142170 598710
rect 170397 598707 170463 598710
rect 256918 598708 256924 598710
rect 256988 598708 256994 598772
rect 376845 598770 376911 598773
rect 374900 598768 376911 598770
rect 374900 598712 376850 598768
rect 376906 598712 376911 598768
rect 374900 598710 376911 598712
rect 376845 598707 376911 598710
rect 499021 598770 499087 598773
rect 532693 598770 532759 598773
rect 499021 598768 532759 598770
rect 499021 598712 499026 598768
rect 499082 598712 532698 598768
rect 532754 598712 532759 598768
rect 499021 598710 532759 598712
rect 499021 598707 499087 598710
rect 532693 598707 532759 598710
rect 134934 598574 142170 598634
rect 500401 598634 500467 598637
rect 534073 598634 534139 598637
rect 500401 598632 534139 598634
rect 500401 598576 500406 598632
rect 500462 598576 534078 598632
rect 534134 598576 534139 598632
rect 500401 598574 534139 598576
rect 500401 598571 500467 598574
rect 534073 598571 534139 598574
rect 58341 598498 58407 598501
rect 174721 598498 174787 598501
rect 258717 598498 258783 598501
rect 494881 598498 494947 598501
rect 528645 598498 528711 598501
rect 58341 598496 60076 598498
rect 58341 598440 58346 598496
rect 58402 598440 60076 598496
rect 58341 598438 60076 598440
rect 174721 598496 180044 598498
rect 174721 598440 174726 598496
rect 174782 598440 180044 598496
rect 174721 598438 180044 598440
rect 258717 598496 300196 598498
rect 258717 598440 258722 598496
rect 258778 598440 300196 598496
rect 258717 598438 300196 598440
rect 494881 598496 528711 598498
rect 494881 598440 494886 598496
rect 494942 598440 528650 598496
rect 528706 598440 528711 598496
rect 494881 598438 528711 598440
rect 58341 598435 58407 598438
rect 174721 598435 174787 598438
rect 258717 598435 258783 598438
rect 494881 598435 494947 598438
rect 528645 598435 528711 598438
rect 497641 598362 497707 598365
rect 531497 598362 531563 598365
rect 497641 598360 531563 598362
rect 497641 598304 497646 598360
rect 497702 598304 531502 598360
rect 531558 598304 531563 598360
rect 497641 598302 531563 598304
rect 497641 598299 497707 598302
rect 531497 598299 531563 598302
rect 532969 598362 533035 598365
rect 536925 598362 536991 598365
rect 532969 598360 536991 598362
rect 532969 598304 532974 598360
rect 533030 598304 536930 598360
rect 536986 598304 536991 598360
rect 532969 598302 536991 598304
rect 532969 598299 533035 598302
rect 536925 598299 536991 598302
rect 490741 598226 490807 598229
rect 538305 598226 538371 598229
rect 490741 598224 538371 598226
rect 490741 598168 490746 598224
rect 490802 598168 538310 598224
rect 538366 598168 538371 598224
rect 490741 598166 538371 598168
rect 490741 598163 490807 598166
rect 538305 598163 538371 598166
rect 504214 598028 504220 598092
rect 504284 598090 504290 598092
rect 504541 598090 504607 598093
rect 504284 598088 504607 598090
rect 504284 598032 504546 598088
rect 504602 598032 504607 598088
rect 504284 598030 504607 598032
rect 504284 598028 504290 598030
rect 504541 598027 504607 598030
rect 505921 598090 505987 598093
rect 505921 598088 506858 598090
rect 505921 598032 505926 598088
rect 505982 598032 506858 598088
rect 505921 598030 506858 598032
rect 505921 598027 505987 598030
rect 170765 597954 170831 597957
rect 256734 597954 256740 597956
rect 142110 597952 170831 597954
rect 134934 597818 134994 597924
rect 142110 597896 170770 597952
rect 170826 597896 170831 597952
rect 142110 597894 170831 597896
rect 254932 597894 256740 597954
rect 142110 597818 142170 597894
rect 170765 597891 170831 597894
rect 256734 597892 256740 597894
rect 256804 597892 256810 597956
rect 376753 597954 376819 597957
rect 374900 597952 376819 597954
rect 374900 597896 376758 597952
rect 376814 597896 376819 597952
rect 374900 597894 376819 597896
rect 506798 597954 506858 598030
rect 506974 598028 506980 598092
rect 507044 598090 507050 598092
rect 507301 598090 507367 598093
rect 507044 598088 507367 598090
rect 507044 598032 507306 598088
rect 507362 598032 507367 598088
rect 507044 598030 507367 598032
rect 507044 598028 507050 598030
rect 507301 598027 507367 598030
rect 509190 598030 528570 598090
rect 509190 597954 509250 598030
rect 506798 597894 509250 597954
rect 376753 597891 376819 597894
rect 134934 597758 142170 597818
rect 528510 597682 528570 598030
rect 533286 598028 533292 598092
rect 533356 598090 533362 598092
rect 533521 598090 533587 598093
rect 533356 598088 533587 598090
rect 533356 598032 533526 598088
rect 533582 598032 533587 598088
rect 533356 598030 533587 598032
rect 533356 598028 533362 598030
rect 533521 598027 533587 598030
rect 534574 598028 534580 598092
rect 534644 598090 534650 598092
rect 534901 598090 534967 598093
rect 534644 598088 534967 598090
rect 534644 598032 534906 598088
rect 534962 598032 534967 598088
rect 534644 598030 534967 598032
rect 534644 598028 534650 598030
rect 534901 598027 534967 598030
rect 529841 597954 529907 597957
rect 544285 597954 544351 597957
rect 529841 597952 544351 597954
rect 529841 597896 529846 597952
rect 529902 597896 544290 597952
rect 544346 597896 544351 597952
rect 529841 597894 544351 597896
rect 529841 597891 529907 597894
rect 544285 597891 544351 597894
rect 531313 597818 531379 597821
rect 534165 597818 534231 597821
rect 531313 597816 534231 597818
rect 531313 597760 531318 597816
rect 531374 597760 534170 597816
rect 534226 597760 534231 597816
rect 531313 597758 534231 597760
rect 531313 597755 531379 597758
rect 534165 597755 534231 597758
rect 535637 597682 535703 597685
rect 528510 597680 535703 597682
rect 528510 597624 535642 597680
rect 535698 597624 535703 597680
rect 528510 597622 535703 597624
rect 535637 597619 535703 597622
rect 295374 597484 295380 597548
rect 295444 597546 295450 597548
rect 296621 597546 296687 597549
rect 295444 597544 296687 597546
rect 295444 597488 296626 597544
rect 296682 597488 296687 597544
rect 295444 597486 296687 597488
rect 295444 597484 295450 597486
rect 296621 597483 296687 597486
rect 299422 597484 299428 597548
rect 299492 597546 299498 597548
rect 299933 597546 299999 597549
rect 299492 597544 299999 597546
rect 299492 597488 299938 597544
rect 299994 597488 299999 597544
rect 299492 597486 299999 597488
rect 299492 597484 299498 597486
rect 299933 597483 299999 597486
rect 54661 597410 54727 597413
rect 179229 597410 179295 597413
rect 258901 597410 258967 597413
rect 54661 597408 60076 597410
rect 54661 597352 54666 597408
rect 54722 597352 60076 597408
rect 54661 597350 60076 597352
rect 179229 597408 180044 597410
rect 179229 597352 179234 597408
rect 179290 597352 180044 597408
rect 179229 597350 180044 597352
rect 258901 597408 300196 597410
rect 258901 597352 258906 597408
rect 258962 597352 300196 597408
rect 258901 597350 300196 597352
rect 54661 597347 54727 597350
rect 179229 597347 179295 597350
rect 258901 597347 258967 597350
rect 174813 597138 174879 597141
rect 296110 597138 296116 597140
rect 142110 597136 174879 597138
rect 134934 597002 134994 597108
rect 142110 597080 174818 597136
rect 174874 597080 174879 597136
rect 142110 597078 174879 597080
rect 254932 597078 296116 597138
rect 142110 597002 142170 597078
rect 174813 597075 174879 597078
rect 296110 597076 296116 597078
rect 296180 597076 296186 597140
rect 376017 597138 376083 597141
rect 374900 597136 376083 597138
rect 374900 597080 376022 597136
rect 376078 597080 376083 597136
rect 374900 597078 376083 597080
rect 376017 597075 376083 597078
rect 134934 596942 142170 597002
rect 171041 596866 171107 596869
rect 173893 596866 173959 596869
rect 400949 596866 401015 596869
rect 416037 596866 416103 596869
rect 171041 596864 178786 596866
rect 171041 596808 171046 596864
rect 171102 596808 173898 596864
rect 173954 596808 178786 596864
rect 171041 596806 178786 596808
rect 171041 596803 171107 596806
rect 173893 596803 173959 596806
rect 178534 596458 178540 596460
rect 134934 596398 178540 596458
rect 56041 596322 56107 596325
rect 56041 596320 60076 596322
rect 56041 596264 56046 596320
rect 56102 596264 60076 596320
rect 134934 596292 134994 596398
rect 178534 596396 178540 596398
rect 178604 596396 178610 596460
rect 178726 596322 178786 596806
rect 400949 596864 416103 596866
rect 400949 596808 400954 596864
rect 401010 596808 416042 596864
rect 416098 596808 416103 596864
rect 400949 596806 416103 596808
rect 400949 596803 401015 596806
rect 416037 596803 416103 596806
rect 292205 596594 292271 596597
rect 292205 596592 300042 596594
rect 292205 596536 292210 596592
rect 292266 596536 300042 596592
rect 292205 596534 300042 596536
rect 292205 596531 292271 596534
rect 299790 596458 299796 596460
rect 254902 596398 299796 596458
rect 56041 596262 60076 596264
rect 178726 596262 180044 596322
rect 254902 596292 254962 596398
rect 299790 596396 299796 596398
rect 299860 596396 299866 596460
rect 56041 596259 56107 596262
rect 295742 596260 295748 596324
rect 295812 596322 295818 596324
rect 296294 596322 296300 596324
rect 295812 596262 296300 596322
rect 295812 596260 295818 596262
rect 296294 596260 296300 596262
rect 296364 596260 296370 596324
rect 299982 596322 300042 596534
rect 378777 596322 378843 596325
rect 299982 596262 300196 596322
rect 374900 596320 378843 596322
rect 374900 596264 378782 596320
rect 378838 596264 378843 596320
rect 374900 596262 378843 596264
rect 378777 596259 378843 596262
rect 296529 596186 296595 596189
rect 296662 596186 296668 596188
rect 296529 596184 296668 596186
rect 296529 596128 296534 596184
rect 296590 596128 296668 596184
rect 296529 596126 296668 596128
rect 296529 596123 296595 596126
rect 296662 596124 296668 596126
rect 296732 596124 296738 596188
rect 134934 595582 142170 595642
rect 134934 595476 134994 595582
rect 142110 595506 142170 595582
rect 176285 595506 176351 595509
rect 299054 595506 299060 595508
rect 142110 595504 176351 595506
rect 142110 595448 176290 595504
rect 176346 595448 176351 595504
rect 142110 595446 176351 595448
rect 254932 595446 299060 595506
rect 176285 595443 176351 595446
rect 299054 595444 299060 595446
rect 299124 595444 299130 595508
rect 376109 595506 376175 595509
rect 374900 595504 376175 595506
rect 374900 595448 376114 595504
rect 376170 595448 376175 595504
rect 374900 595446 376175 595448
rect 376109 595443 376175 595446
rect 49509 595234 49575 595237
rect 162393 595234 162459 595237
rect 259085 595234 259151 595237
rect 49509 595232 60076 595234
rect 49509 595176 49514 595232
rect 49570 595176 60076 595232
rect 49509 595174 60076 595176
rect 162393 595232 180044 595234
rect 162393 595176 162398 595232
rect 162454 595176 180044 595232
rect 162393 595174 180044 595176
rect 259085 595232 300196 595234
rect 259085 595176 259090 595232
rect 259146 595176 300196 595232
rect 259085 595174 300196 595176
rect 49509 595171 49575 595174
rect 162393 595171 162459 595174
rect 179830 594962 179890 595174
rect 259085 595171 259151 595174
rect 179965 594962 180031 594965
rect 179830 594960 180031 594962
rect 179830 594904 179970 594960
rect 180026 594904 180031 594960
rect 179830 594902 180031 594904
rect 179965 594899 180031 594902
rect 298318 594764 298324 594828
rect 298388 594826 298394 594828
rect 299197 594826 299263 594829
rect 298388 594824 299263 594826
rect 298388 594768 299202 594824
rect 299258 594768 299263 594824
rect 298388 594766 299263 594768
rect 298388 594764 298394 594766
rect 299197 594763 299263 594766
rect 162117 594690 162183 594693
rect 291694 594690 291700 594692
rect 142110 594688 162183 594690
rect 134934 594554 134994 594660
rect 142110 594632 162122 594688
rect 162178 594632 162183 594688
rect 142110 594630 162183 594632
rect 254932 594630 291700 594690
rect 142110 594554 142170 594630
rect 162117 594627 162183 594630
rect 291694 594628 291700 594630
rect 291764 594628 291770 594692
rect 377949 594690 378015 594693
rect 374900 594688 378015 594690
rect 374900 594632 377954 594688
rect 378010 594632 378015 594688
rect 374900 594630 378015 594632
rect 377949 594627 378015 594630
rect 134934 594494 142170 594554
rect 46749 594146 46815 594149
rect 170857 594146 170923 594149
rect 255957 594146 256023 594149
rect 46749 594144 60076 594146
rect 46749 594088 46754 594144
rect 46810 594088 60076 594144
rect 46749 594086 60076 594088
rect 170857 594144 180044 594146
rect 170857 594088 170862 594144
rect 170918 594088 180044 594144
rect 170857 594086 180044 594088
rect 255957 594144 300196 594146
rect 255957 594088 255962 594144
rect 256018 594088 300196 594144
rect 255957 594086 300196 594088
rect 46749 594083 46815 594086
rect 170857 594083 170923 594086
rect 255957 594083 256023 594086
rect 134934 593950 142170 594010
rect 134934 593844 134994 593950
rect 142110 593874 142170 593950
rect 174721 593874 174787 593877
rect 283966 593874 283972 593876
rect 142110 593872 174787 593874
rect 142110 593816 174726 593872
rect 174782 593816 174787 593872
rect 142110 593814 174787 593816
rect 254932 593814 283972 593874
rect 174721 593811 174787 593814
rect 283966 593812 283972 593814
rect 284036 593812 284042 593876
rect 378041 593874 378107 593877
rect 374900 593872 378107 593874
rect 374900 593816 378046 593872
rect 378102 593816 378107 593872
rect 374900 593814 378107 593816
rect 378041 593811 378107 593814
rect -960 592908 480 593148
rect 57513 593058 57579 593061
rect 178033 593058 178099 593061
rect 179045 593058 179111 593061
rect 294597 593058 294663 593061
rect 378041 593058 378107 593061
rect 57513 593056 60076 593058
rect 57513 593000 57518 593056
rect 57574 593000 60076 593056
rect 178033 593056 180044 593058
rect 57513 592998 60076 593000
rect 57513 592995 57579 592998
rect 134934 592514 134994 593028
rect 178033 593000 178038 593056
rect 178094 593000 179050 593056
rect 179106 593000 180044 593056
rect 294597 593056 300196 593058
rect 178033 592998 180044 593000
rect 178033 592995 178099 592998
rect 179045 592995 179111 592998
rect 254902 592922 254962 593028
rect 294597 593000 294602 593056
rect 294658 593000 300196 593056
rect 294597 592998 300196 593000
rect 374900 593056 378107 593058
rect 374900 593000 378046 593056
rect 378102 593000 378107 593056
rect 374900 592998 378107 593000
rect 294597 592995 294663 592998
rect 378041 592995 378107 592998
rect 298870 592922 298876 592924
rect 254902 592862 298876 592922
rect 298870 592860 298876 592862
rect 298940 592860 298946 592924
rect 137737 592514 137803 592517
rect 134934 592512 137803 592514
rect 134934 592456 137742 592512
rect 137798 592456 137803 592512
rect 134934 592454 137803 592456
rect 137737 592451 137803 592454
rect 134934 592318 142170 592378
rect 134934 592212 134994 592318
rect 142110 592242 142170 592318
rect 170673 592242 170739 592245
rect 281022 592242 281028 592244
rect 142110 592240 170739 592242
rect 142110 592184 170678 592240
rect 170734 592184 170739 592240
rect 142110 592182 170739 592184
rect 254932 592182 281028 592242
rect 170673 592179 170739 592182
rect 281022 592180 281028 592182
rect 281092 592180 281098 592244
rect 378041 592242 378107 592245
rect 374900 592240 378107 592242
rect 374900 592184 378046 592240
rect 378102 592184 378107 592240
rect 374900 592182 378107 592184
rect 378041 592179 378107 592182
rect 162485 592106 162551 592109
rect 178033 592106 178099 592109
rect 162485 592104 178099 592106
rect 162485 592048 162490 592104
rect 162546 592048 178038 592104
rect 178094 592048 178099 592104
rect 162485 592046 178099 592048
rect 162485 592043 162551 592046
rect 178033 592043 178099 592046
rect 298502 592044 298508 592108
rect 298572 592106 298578 592108
rect 299289 592106 299355 592109
rect 298572 592104 299355 592106
rect 298572 592048 299294 592104
rect 299350 592048 299355 592104
rect 298572 592046 299355 592048
rect 298572 592044 298578 592046
rect 299289 592043 299355 592046
rect 45093 591970 45159 591973
rect 169385 591970 169451 591973
rect 259361 591970 259427 591973
rect 45093 591968 60076 591970
rect 45093 591912 45098 591968
rect 45154 591912 60076 591968
rect 45093 591910 60076 591912
rect 169385 591968 180044 591970
rect 169385 591912 169390 591968
rect 169446 591912 180044 591968
rect 169385 591910 180044 591912
rect 259361 591968 300196 591970
rect 259361 591912 259366 591968
rect 259422 591912 300196 591968
rect 259361 591910 300196 591912
rect 45093 591907 45159 591910
rect 169385 591907 169451 591910
rect 259361 591907 259427 591910
rect 134934 591502 142170 591562
rect 134934 591396 134994 591502
rect 142110 591426 142170 591502
rect 163497 591426 163563 591429
rect 285254 591426 285260 591428
rect 142110 591424 163563 591426
rect 142110 591368 163502 591424
rect 163558 591368 163563 591424
rect 142110 591366 163563 591368
rect 254932 591366 285260 591426
rect 163497 591363 163563 591366
rect 285254 591364 285260 591366
rect 285324 591364 285330 591428
rect 378041 591426 378107 591429
rect 374900 591424 378107 591426
rect 374900 591368 378046 591424
rect 378102 591368 378107 591424
rect 374900 591366 378107 591368
rect 378041 591363 378107 591366
rect 580206 590956 580212 591020
rect 580276 591018 580282 591020
rect 583520 591018 584960 591108
rect 580276 590958 584960 591018
rect 580276 590956 580282 590958
rect 45369 590882 45435 590885
rect 169569 590882 169635 590885
rect 292021 590882 292087 590885
rect 45369 590880 60076 590882
rect 45369 590824 45374 590880
rect 45430 590824 60076 590880
rect 45369 590822 60076 590824
rect 169569 590880 180044 590882
rect 169569 590824 169574 590880
rect 169630 590824 180044 590880
rect 169569 590822 180044 590824
rect 292021 590880 300196 590882
rect 292021 590824 292026 590880
rect 292082 590824 300196 590880
rect 583520 590868 584960 590958
rect 292021 590822 300196 590824
rect 45369 590819 45435 590822
rect 169569 590819 169635 590822
rect 292021 590819 292087 590822
rect 166625 590610 166691 590613
rect 142110 590608 166691 590610
rect 134934 590474 134994 590580
rect 142110 590552 166630 590608
rect 166686 590552 166691 590608
rect 142110 590550 166691 590552
rect 254932 590550 277410 590610
rect 142110 590474 142170 590550
rect 166625 590547 166691 590550
rect 134934 590414 142170 590474
rect 277350 590338 277410 590550
rect 294454 590548 294460 590612
rect 294524 590610 294530 590612
rect 295149 590610 295215 590613
rect 378041 590610 378107 590613
rect 294524 590608 295215 590610
rect 294524 590552 295154 590608
rect 295210 590552 295215 590608
rect 294524 590550 295215 590552
rect 374900 590608 378107 590610
rect 374900 590552 378046 590608
rect 378102 590552 378107 590608
rect 374900 590550 378107 590552
rect 294524 590548 294530 590550
rect 295149 590547 295215 590550
rect 378041 590547 378107 590550
rect 294822 590338 294828 590340
rect 277350 590278 294828 590338
rect 294822 590276 294828 590278
rect 294892 590276 294898 590340
rect 134934 589870 142170 589930
rect 45185 589794 45251 589797
rect 45185 589792 60076 589794
rect 45185 589736 45190 589792
rect 45246 589736 60076 589792
rect 134934 589764 134994 589870
rect 142110 589794 142170 589870
rect 167729 589794 167795 589797
rect 256049 589794 256115 589797
rect 378041 589794 378107 589797
rect 142110 589792 167795 589794
rect 45185 589734 60076 589736
rect 142110 589736 167734 589792
rect 167790 589736 167795 589792
rect 142110 589734 167795 589736
rect 45185 589731 45251 589734
rect 167729 589731 167795 589734
rect 171090 589734 180044 589794
rect 256049 589792 300196 589794
rect 164969 589658 165035 589661
rect 171090 589658 171150 589734
rect 164969 589656 171150 589658
rect 164969 589600 164974 589656
rect 165030 589600 171150 589656
rect 164969 589598 171150 589600
rect 254902 589658 254962 589764
rect 256049 589736 256054 589792
rect 256110 589736 300196 589792
rect 256049 589734 300196 589736
rect 374900 589792 378107 589794
rect 374900 589736 378046 589792
rect 378102 589736 378107 589792
rect 374900 589734 378107 589736
rect 256049 589731 256115 589734
rect 378041 589731 378107 589734
rect 283782 589658 283788 589660
rect 254902 589598 283788 589658
rect 164969 589595 165035 589598
rect 283782 589596 283788 589598
rect 283852 589596 283858 589660
rect 294638 589188 294644 589252
rect 294708 589250 294714 589252
rect 295057 589250 295123 589253
rect 294708 589248 295123 589250
rect 294708 589192 295062 589248
rect 295118 589192 295123 589248
rect 294708 589190 295123 589192
rect 294708 589188 294714 589190
rect 295057 589187 295123 589190
rect 294454 588978 294460 588980
rect 54661 588706 54727 588709
rect 54661 588704 60076 588706
rect 54661 588648 54666 588704
rect 54722 588648 60076 588704
rect 54661 588646 60076 588648
rect 54661 588643 54727 588646
rect 134934 588434 134994 588948
rect 254932 588918 294460 588978
rect 294454 588916 294460 588918
rect 294524 588916 294530 588980
rect 376937 588978 377003 588981
rect 374900 588976 377003 588978
rect 374900 588920 376942 588976
rect 376998 588920 377003 588976
rect 374900 588918 377003 588920
rect 376937 588915 377003 588918
rect 176561 588706 176627 588709
rect 254577 588706 254643 588709
rect 176561 588704 180044 588706
rect 176561 588648 176566 588704
rect 176622 588648 180044 588704
rect 176561 588646 180044 588648
rect 254577 588704 300196 588706
rect 254577 588648 254582 588704
rect 254638 588648 300196 588704
rect 254577 588646 300196 588648
rect 176561 588643 176627 588646
rect 254577 588643 254643 588646
rect 137921 588434 137987 588437
rect 134934 588432 137987 588434
rect 134934 588376 137926 588432
rect 137982 588376 137987 588432
rect 134934 588374 137987 588376
rect 137921 588371 137987 588374
rect 134934 588238 142170 588298
rect 134934 588132 134994 588238
rect 142110 588162 142170 588238
rect 170305 588162 170371 588165
rect 289302 588162 289308 588164
rect 142110 588160 170371 588162
rect 142110 588104 170310 588160
rect 170366 588104 170371 588160
rect 142110 588102 170371 588104
rect 254932 588102 289308 588162
rect 170305 588099 170371 588102
rect 289302 588100 289308 588102
rect 289372 588100 289378 588164
rect 378041 588162 378107 588165
rect 374900 588160 378107 588162
rect 374900 588104 378046 588160
rect 378102 588104 378107 588160
rect 374900 588102 378107 588104
rect 378041 588099 378107 588102
rect 165153 588026 165219 588029
rect 176561 588026 176627 588029
rect 165153 588024 176627 588026
rect 165153 587968 165158 588024
rect 165214 587968 176566 588024
rect 176622 587968 176627 588024
rect 165153 587966 176627 587968
rect 165153 587963 165219 587966
rect 176561 587963 176627 587966
rect 49417 587618 49483 587621
rect 173709 587618 173775 587621
rect 256417 587618 256483 587621
rect 49417 587616 60076 587618
rect 49417 587560 49422 587616
rect 49478 587560 60076 587616
rect 49417 587558 60076 587560
rect 173709 587616 180044 587618
rect 173709 587560 173714 587616
rect 173770 587560 180044 587616
rect 173709 587558 180044 587560
rect 256417 587616 300196 587618
rect 256417 587560 256422 587616
rect 256478 587560 300196 587616
rect 256417 587558 300196 587560
rect 49417 587555 49483 587558
rect 173709 587555 173775 587558
rect 256417 587555 256483 587558
rect 134934 587422 142170 587482
rect 134934 587316 134994 587422
rect 142110 587346 142170 587422
rect 173525 587346 173591 587349
rect 294638 587346 294644 587348
rect 142110 587344 173591 587346
rect 142110 587288 173530 587344
rect 173586 587288 173591 587344
rect 142110 587286 173591 587288
rect 254932 587286 294644 587346
rect 173525 587283 173591 587286
rect 294638 587284 294644 587286
rect 294708 587284 294714 587348
rect 377765 587346 377831 587349
rect 374900 587344 377831 587346
rect 374900 587288 377770 587344
rect 377826 587288 377831 587344
rect 374900 587286 377831 587288
rect 377765 587283 377831 587286
rect 296529 587210 296595 587213
rect 296713 587210 296779 587213
rect 296529 587208 296779 587210
rect 296529 587152 296534 587208
rect 296590 587152 296718 587208
rect 296774 587152 296779 587208
rect 296529 587150 296779 587152
rect 296529 587147 296595 587150
rect 296713 587147 296779 587150
rect 178718 586802 178724 586804
rect 134934 586742 178724 586802
rect 59494 586470 60076 586530
rect 134934 586500 134994 586742
rect 178718 586740 178724 586742
rect 178788 586740 178794 586804
rect 296670 586742 299674 586802
rect 292113 586666 292179 586669
rect 296670 586666 296730 586742
rect 287010 586606 287898 586666
rect 179462 586470 180044 586530
rect 254932 586470 263610 586530
rect 49325 586394 49391 586397
rect 59494 586394 59554 586470
rect 49325 586392 59554 586394
rect 49325 586336 49330 586392
rect 49386 586336 59554 586392
rect 49325 586334 59554 586336
rect 172421 586394 172487 586397
rect 179462 586394 179522 586470
rect 172421 586392 179522 586394
rect 172421 586336 172426 586392
rect 172482 586336 179522 586392
rect 172421 586334 179522 586336
rect 263550 586394 263610 586470
rect 287010 586394 287070 586606
rect 287838 586532 287898 586606
rect 292113 586664 296730 586666
rect 292113 586608 292118 586664
rect 292174 586608 296730 586664
rect 292113 586606 296730 586608
rect 292113 586603 292179 586606
rect 294965 586532 295031 586533
rect 287830 586468 287836 586532
rect 287900 586468 287906 586532
rect 294965 586530 295012 586532
rect 294920 586528 295012 586530
rect 294920 586472 294970 586528
rect 294920 586470 295012 586472
rect 294965 586468 295012 586470
rect 295076 586468 295082 586532
rect 296713 586530 296779 586533
rect 296670 586528 296779 586530
rect 296670 586472 296718 586528
rect 296774 586472 296779 586528
rect 294965 586467 295031 586468
rect 296670 586467 296779 586472
rect 299614 586530 299674 586742
rect 378041 586530 378107 586533
rect 299614 586470 300196 586530
rect 374900 586470 375482 586530
rect 263550 586334 287070 586394
rect 296529 586394 296595 586397
rect 296670 586394 296730 586467
rect 296529 586392 296730 586394
rect 296529 586336 296534 586392
rect 296590 586336 296730 586392
rect 296529 586334 296730 586336
rect 375422 586394 375482 586470
rect 377814 586528 378107 586530
rect 377814 586472 378046 586528
rect 378102 586472 378107 586528
rect 377814 586470 378107 586472
rect 377814 586394 377874 586470
rect 378041 586467 378107 586470
rect 375422 586334 377874 586394
rect 49325 586331 49391 586334
rect 172421 586331 172487 586334
rect 296529 586331 296595 586334
rect 174905 585714 174971 585717
rect 290958 585714 290964 585716
rect 142110 585712 174971 585714
rect 134934 585578 134994 585684
rect 142110 585656 174910 585712
rect 174966 585656 174971 585712
rect 142110 585654 174971 585656
rect 254932 585654 290964 585714
rect 142110 585578 142170 585654
rect 174905 585651 174971 585654
rect 290958 585652 290964 585654
rect 291028 585652 291034 585716
rect 378041 585714 378107 585717
rect 374900 585712 378107 585714
rect 374900 585656 378046 585712
rect 378102 585656 378107 585712
rect 374900 585654 378107 585656
rect 378041 585651 378107 585654
rect 134934 585518 142170 585578
rect 49233 585442 49299 585445
rect 256325 585442 256391 585445
rect 49233 585440 60076 585442
rect 49233 585384 49238 585440
rect 49294 585384 60076 585440
rect 49233 585382 60076 585384
rect 175414 585382 180044 585442
rect 256325 585440 300196 585442
rect 256325 585384 256330 585440
rect 256386 585384 300196 585440
rect 256325 585382 300196 585384
rect 49233 585379 49299 585382
rect 168281 585306 168347 585309
rect 175181 585306 175247 585309
rect 168281 585304 175247 585306
rect 168281 585248 168286 585304
rect 168342 585248 175186 585304
rect 175242 585248 175247 585304
rect 168281 585246 175247 585248
rect 168281 585243 168347 585246
rect 175181 585243 175247 585246
rect 168097 585170 168163 585173
rect 175089 585170 175155 585173
rect 175414 585170 175474 585382
rect 256325 585379 256391 585382
rect 168097 585168 175474 585170
rect 168097 585112 168102 585168
rect 168158 585112 175094 585168
rect 175150 585112 175474 585168
rect 168097 585110 175474 585112
rect 168097 585107 168163 585110
rect 175089 585107 175155 585110
rect 290590 585108 290596 585172
rect 290660 585170 290666 585172
rect 291101 585170 291167 585173
rect 290660 585168 291167 585170
rect 290660 585112 291106 585168
rect 291162 585112 291167 585168
rect 290660 585110 291167 585112
rect 290660 585108 290666 585110
rect 291101 585107 291167 585110
rect 175825 584898 175891 584901
rect 288198 584898 288204 584900
rect 142110 584896 175891 584898
rect 134934 584762 134994 584868
rect 142110 584840 175830 584896
rect 175886 584840 175891 584896
rect 142110 584838 175891 584840
rect 254932 584838 288204 584898
rect 142110 584762 142170 584838
rect 175825 584835 175891 584838
rect 288198 584836 288204 584838
rect 288268 584836 288274 584900
rect 378041 584898 378107 584901
rect 374900 584896 378107 584898
rect 374900 584840 378046 584896
rect 378102 584840 378107 584896
rect 374900 584838 378107 584840
rect 378041 584835 378107 584838
rect 134934 584702 142170 584762
rect 54569 584354 54635 584357
rect 175181 584354 175247 584357
rect 176377 584354 176443 584357
rect 255865 584354 255931 584357
rect 54569 584352 60076 584354
rect 54569 584296 54574 584352
rect 54630 584296 60076 584352
rect 54569 584294 60076 584296
rect 175181 584352 180044 584354
rect 175181 584296 175186 584352
rect 175242 584296 176382 584352
rect 176438 584296 180044 584352
rect 175181 584294 180044 584296
rect 255865 584352 300196 584354
rect 255865 584296 255870 584352
rect 255926 584296 300196 584352
rect 255865 584294 300196 584296
rect 54569 584291 54635 584294
rect 175181 584291 175247 584294
rect 176377 584291 176443 584294
rect 255865 584291 255931 584294
rect 178585 584082 178651 584085
rect 286358 584082 286364 584084
rect 142110 584080 178651 584082
rect 134934 583946 134994 584052
rect 142110 584024 178590 584080
rect 178646 584024 178651 584080
rect 142110 584022 178651 584024
rect 254932 584022 286364 584082
rect 142110 583946 142170 584022
rect 178585 584019 178651 584022
rect 286358 584020 286364 584022
rect 286428 584020 286434 584084
rect 378041 584082 378107 584085
rect 374900 584080 378107 584082
rect 374900 584024 378046 584080
rect 378102 584024 378107 584080
rect 374900 584022 378107 584024
rect 378041 584019 378107 584022
rect 134934 583886 142170 583946
rect 55121 583266 55187 583269
rect 172145 583266 172211 583269
rect 285070 583266 285076 583268
rect 55121 583264 60076 583266
rect 55121 583208 55126 583264
rect 55182 583208 60076 583264
rect 172145 583264 180044 583266
rect 55121 583206 60076 583208
rect 55121 583203 55187 583206
rect 134934 583130 134994 583236
rect 172145 583208 172150 583264
rect 172206 583208 180044 583264
rect 172145 583206 180044 583208
rect 254932 583206 285076 583266
rect 172145 583203 172211 583206
rect 285070 583204 285076 583206
rect 285140 583204 285146 583268
rect 292389 583266 292455 583269
rect 378041 583266 378107 583269
rect 292389 583264 300196 583266
rect 292389 583208 292394 583264
rect 292450 583208 300196 583264
rect 292389 583206 300196 583208
rect 374900 583264 378107 583266
rect 374900 583208 378046 583264
rect 378102 583208 378107 583264
rect 374900 583206 378107 583208
rect 292389 583203 292455 583206
rect 378041 583203 378107 583206
rect 176193 583130 176259 583133
rect 134934 583128 176259 583130
rect 134934 583072 176198 583128
rect 176254 583072 176259 583128
rect 134934 583070 176259 583072
rect 176193 583067 176259 583070
rect 176469 582586 176535 582589
rect 134934 582584 176535 582586
rect 134934 582528 176474 582584
rect 176530 582528 176535 582584
rect 134934 582526 176535 582528
rect 134934 582420 134994 582526
rect 176469 582523 176535 582526
rect 283414 582450 283420 582452
rect 254932 582390 283420 582450
rect 283414 582388 283420 582390
rect 283484 582388 283490 582452
rect 378041 582450 378107 582453
rect 374900 582448 378107 582450
rect 374900 582392 378046 582448
rect 378102 582392 378107 582448
rect 374900 582390 378107 582392
rect 378041 582387 378107 582390
rect 43897 582178 43963 582181
rect 166901 582178 166967 582181
rect 256233 582178 256299 582181
rect 43897 582176 60076 582178
rect 43897 582120 43902 582176
rect 43958 582120 60076 582176
rect 43897 582118 60076 582120
rect 166901 582176 180044 582178
rect 166901 582120 166906 582176
rect 166962 582120 180044 582176
rect 166901 582118 180044 582120
rect 256233 582176 300196 582178
rect 256233 582120 256238 582176
rect 256294 582120 300196 582176
rect 256233 582118 300196 582120
rect 43897 582115 43963 582118
rect 166901 582115 166967 582118
rect 256233 582115 256299 582118
rect 159357 581634 159423 581637
rect 283598 581634 283604 581636
rect 142110 581632 159423 581634
rect 134934 581498 134994 581604
rect 142110 581576 159362 581632
rect 159418 581576 159423 581632
rect 142110 581574 159423 581576
rect 254932 581574 283604 581634
rect 142110 581498 142170 581574
rect 159357 581571 159423 581574
rect 283598 581572 283604 581574
rect 283668 581572 283674 581636
rect 377857 581634 377923 581637
rect 374900 581632 377923 581634
rect 374900 581576 377862 581632
rect 377918 581576 377923 581632
rect 374900 581574 377923 581576
rect 377857 581571 377923 581574
rect 134934 581438 142170 581498
rect 159541 581226 159607 581229
rect 166901 581226 166967 581229
rect 159541 581224 166967 581226
rect 159541 581168 159546 581224
rect 159602 581168 166906 581224
rect 166962 581168 166967 581224
rect 159541 581166 166967 581168
rect 159541 581163 159607 581166
rect 166901 581163 166967 581166
rect 289169 581226 289235 581229
rect 289169 581224 296730 581226
rect 289169 581168 289174 581224
rect 289230 581168 296730 581224
rect 289169 581166 296730 581168
rect 289169 581163 289235 581166
rect 47945 581090 48011 581093
rect 159725 581090 159791 581093
rect 169477 581090 169543 581093
rect 290917 581092 290983 581093
rect 47945 581088 60076 581090
rect 47945 581032 47950 581088
rect 48006 581032 60076 581088
rect 47945 581030 60076 581032
rect 159725 581088 180044 581090
rect 159725 581032 159730 581088
rect 159786 581032 169482 581088
rect 169538 581032 180044 581088
rect 159725 581030 180044 581032
rect 290917 581088 290964 581092
rect 291028 581090 291034 581092
rect 296670 581090 296730 581166
rect 290917 581032 290922 581088
rect 47945 581027 48011 581030
rect 159725 581027 159791 581030
rect 169477 581027 169543 581030
rect 290917 581028 290964 581032
rect 291028 581030 291074 581090
rect 296670 581030 300196 581090
rect 291028 581028 291034 581030
rect 290917 581027 290983 581028
rect 290774 580892 290780 580956
rect 290844 580954 290850 580956
rect 291009 580954 291075 580957
rect 290844 580952 291075 580954
rect 290844 580896 291014 580952
rect 291070 580896 291075 580952
rect 290844 580894 291075 580896
rect 290844 580892 290850 580894
rect 291009 580891 291075 580894
rect 178861 580818 178927 580821
rect 290958 580818 290964 580820
rect 142110 580816 178927 580818
rect 134934 580682 134994 580788
rect 142110 580760 178866 580816
rect 178922 580760 178927 580816
rect 142110 580758 178927 580760
rect 254932 580758 290964 580818
rect 142110 580682 142170 580758
rect 178861 580755 178927 580758
rect 290958 580756 290964 580758
rect 291028 580756 291034 580820
rect 377121 580818 377187 580821
rect 374900 580816 377187 580818
rect 374900 580760 377126 580816
rect 377182 580760 377187 580816
rect 374900 580758 377187 580760
rect 377121 580755 377187 580758
rect 134934 580622 142170 580682
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 46657 580002 46723 580005
rect 289261 580002 289327 580005
rect 377581 580002 377647 580005
rect 46657 580000 60076 580002
rect 46657 579944 46662 580000
rect 46718 579944 60076 580000
rect 46657 579942 60076 579944
rect 46657 579939 46723 579942
rect 134934 579866 134994 579972
rect 176334 579942 180044 580002
rect 289261 580000 300196 580002
rect 176101 579866 176167 579869
rect 134934 579864 176167 579866
rect 134934 579808 176106 579864
rect 176162 579808 176167 579864
rect 134934 579806 176167 579808
rect 176101 579803 176167 579806
rect 159449 579730 159515 579733
rect 172973 579730 173039 579733
rect 176334 579730 176394 579942
rect 254902 579866 254962 579972
rect 289261 579944 289266 580000
rect 289322 579944 300196 580000
rect 289261 579942 300196 579944
rect 374900 580000 377647 580002
rect 374900 579944 377586 580000
rect 377642 579944 377647 580000
rect 374900 579942 377647 579944
rect 289261 579939 289327 579942
rect 377581 579939 377647 579942
rect 289486 579866 289492 579868
rect 254902 579806 289492 579866
rect 289486 579804 289492 579806
rect 289556 579804 289562 579868
rect 159449 579728 176394 579730
rect 159449 579672 159454 579728
rect 159510 579672 172978 579728
rect 173034 579672 176394 579728
rect 159449 579670 176394 579672
rect 159449 579667 159515 579670
rect 172973 579667 173039 579670
rect 179229 579186 179295 579189
rect 293166 579186 293172 579188
rect 142110 579184 179295 579186
rect 134934 579050 134994 579156
rect 142110 579128 179234 579184
rect 179290 579128 179295 579184
rect 142110 579126 179295 579128
rect 254932 579126 293172 579186
rect 142110 579050 142170 579126
rect 179229 579123 179295 579126
rect 293166 579124 293172 579126
rect 293236 579124 293242 579188
rect 377029 579186 377095 579189
rect 374900 579184 377095 579186
rect 374900 579128 377034 579184
rect 377090 579128 377095 579184
rect 374900 579126 377095 579128
rect 377029 579123 377095 579126
rect 134934 578990 142170 579050
rect 44909 578914 44975 578917
rect 256141 578914 256207 578917
rect 44909 578912 60076 578914
rect 44909 578856 44914 578912
rect 44970 578856 60076 578912
rect 44909 578854 60076 578856
rect 171090 578854 180044 578914
rect 256141 578912 300196 578914
rect 256141 578856 256146 578912
rect 256202 578856 300196 578912
rect 256141 578854 300196 578856
rect 44909 578851 44975 578854
rect 159633 578506 159699 578509
rect 169937 578506 170003 578509
rect 171090 578506 171150 578854
rect 256141 578851 256207 578854
rect 134934 578446 142170 578506
rect 134934 578340 134994 578446
rect 142110 578370 142170 578446
rect 159633 578504 171150 578506
rect 159633 578448 159638 578504
rect 159694 578448 169942 578504
rect 169998 578448 171150 578504
rect 159633 578446 171150 578448
rect 159633 578443 159699 578446
rect 169937 578443 170003 578446
rect 178953 578370 179019 578373
rect 290590 578370 290596 578372
rect 142110 578368 179019 578370
rect 142110 578312 178958 578368
rect 179014 578312 179019 578368
rect 142110 578310 179019 578312
rect 254932 578310 290596 578370
rect 178953 578307 179019 578310
rect 290590 578308 290596 578310
rect 290660 578308 290666 578372
rect 377857 578370 377923 578373
rect 374900 578368 377923 578370
rect 374900 578312 377862 578368
rect 377918 578312 377923 578368
rect 374900 578310 377923 578312
rect 377857 578307 377923 578310
rect 287094 578172 287100 578236
rect 287164 578234 287170 578236
rect 288341 578234 288407 578237
rect 287164 578232 288407 578234
rect 287164 578176 288346 578232
rect 288402 578176 288407 578232
rect 287164 578174 288407 578176
rect 287164 578172 287170 578174
rect 288341 578171 288407 578174
rect 46565 577826 46631 577829
rect 169661 577826 169727 577829
rect 255037 577826 255103 577829
rect 46565 577824 60076 577826
rect 46565 577768 46570 577824
rect 46626 577768 60076 577824
rect 46565 577766 60076 577768
rect 169661 577824 180044 577826
rect 169661 577768 169666 577824
rect 169722 577768 180044 577824
rect 169661 577766 180044 577768
rect 255037 577824 300196 577826
rect 255037 577768 255042 577824
rect 255098 577768 300196 577824
rect 255037 577766 300196 577768
rect 46565 577763 46631 577766
rect 169661 577763 169727 577766
rect 255037 577763 255103 577766
rect 551134 577628 551140 577692
rect 551204 577690 551210 577692
rect 583520 577690 584960 577780
rect 551204 577630 584960 577690
rect 551204 577628 551210 577630
rect 179137 577554 179203 577557
rect 288014 577554 288020 577556
rect 142110 577552 179203 577554
rect 134934 577418 134994 577524
rect 142110 577496 179142 577552
rect 179198 577496 179203 577552
rect 142110 577494 179203 577496
rect 254932 577494 288020 577554
rect 142110 577418 142170 577494
rect 179137 577491 179203 577494
rect 288014 577492 288020 577494
rect 288084 577492 288090 577556
rect 379462 577554 379468 577556
rect 374900 577494 379468 577554
rect 379462 577492 379468 577494
rect 379532 577492 379538 577556
rect 583520 577540 584960 577630
rect 134934 577358 142170 577418
rect 296529 577418 296595 577421
rect 296662 577418 296668 577420
rect 296529 577416 296668 577418
rect 296529 577360 296534 577416
rect 296590 577360 296668 577416
rect 296529 577358 296668 577360
rect 296529 577355 296595 577358
rect 296662 577356 296668 577358
rect 296732 577356 296738 577420
rect 162761 576874 162827 576877
rect 169661 576874 169727 576877
rect 162761 576872 169727 576874
rect 162761 576816 162766 576872
rect 162822 576816 169666 576872
rect 169722 576816 169727 576872
rect 162761 576814 169727 576816
rect 162761 576811 162827 576814
rect 169661 576811 169727 576814
rect 44817 576738 44883 576741
rect 179321 576738 179387 576741
rect 179873 576738 179939 576741
rect 292062 576738 292068 576740
rect 44817 576736 60076 576738
rect 44817 576680 44822 576736
rect 44878 576680 60076 576736
rect 142110 576736 179387 576738
rect 44817 576678 60076 576680
rect 44817 576675 44883 576678
rect 134934 576602 134994 576708
rect 142110 576680 179326 576736
rect 179382 576680 179387 576736
rect 142110 576678 179387 576680
rect 142110 576602 142170 576678
rect 179321 576675 179387 576678
rect 179462 576736 180044 576738
rect 179462 576680 179878 576736
rect 179934 576680 180044 576736
rect 179462 576678 180044 576680
rect 254932 576678 292068 576738
rect 134934 576542 142170 576602
rect 162669 576602 162735 576605
rect 179462 576602 179522 576678
rect 179873 576675 179939 576678
rect 292062 576676 292068 576678
rect 292132 576676 292138 576740
rect 296529 576738 296595 576741
rect 296662 576738 296668 576740
rect 296529 576736 296668 576738
rect 296529 576680 296534 576736
rect 296590 576680 296668 576736
rect 296529 576678 296668 576680
rect 296529 576675 296595 576678
rect 296662 576676 296668 576678
rect 296732 576676 296738 576740
rect 380985 576738 381051 576741
rect 298326 576678 300196 576738
rect 374900 576736 381051 576738
rect 374900 576680 380990 576736
rect 381046 576680 381051 576736
rect 374900 576678 381051 576680
rect 298326 576602 298386 576678
rect 380985 576675 381051 576678
rect 162669 576600 179522 576602
rect 162669 576544 162674 576600
rect 162730 576544 179522 576600
rect 162669 576542 179522 576544
rect 258030 576542 298386 576602
rect 162669 576539 162735 576542
rect 254945 576466 255011 576469
rect 258030 576466 258090 576542
rect 254945 576464 258090 576466
rect 254945 576408 254950 576464
rect 255006 576408 258090 576464
rect 254945 576406 258090 576408
rect 254945 576403 255011 576406
rect 257102 575922 257108 575924
rect 47853 575650 47919 575653
rect 47853 575648 60076 575650
rect 47853 575592 47858 575648
rect 47914 575592 60076 575648
rect 47853 575590 60076 575592
rect 47853 575587 47919 575590
rect 134934 575514 134994 575892
rect 254932 575862 257108 575922
rect 257102 575860 257108 575862
rect 257172 575860 257178 575924
rect 377121 575922 377187 575925
rect 374900 575920 377187 575922
rect 374900 575864 377126 575920
rect 377182 575864 377187 575920
rect 374900 575862 377187 575864
rect 377121 575859 377187 575862
rect 173709 575650 173775 575653
rect 254761 575650 254827 575653
rect 173709 575648 180044 575650
rect 173709 575592 173714 575648
rect 173770 575592 180044 575648
rect 173709 575590 180044 575592
rect 254761 575648 300196 575650
rect 254761 575592 254766 575648
rect 254822 575592 300196 575648
rect 254761 575590 300196 575592
rect 173709 575587 173775 575590
rect 254761 575587 254827 575590
rect 137185 575514 137251 575517
rect 134934 575512 137251 575514
rect 134934 575456 137190 575512
rect 137246 575456 137251 575512
rect 134934 575454 137251 575456
rect 137185 575451 137251 575454
rect 256918 575452 256924 575516
rect 256988 575514 256994 575516
rect 257705 575514 257771 575517
rect 256988 575512 257771 575514
rect 256988 575456 257710 575512
rect 257766 575456 257771 575512
rect 256988 575454 257771 575456
rect 256988 575452 256994 575454
rect 257705 575451 257771 575454
rect 134934 575182 142170 575242
rect 134934 575076 134994 575182
rect 142110 575106 142170 575182
rect 173065 575106 173131 575109
rect 291878 575106 291884 575108
rect 142110 575104 173131 575106
rect 142110 575048 173070 575104
rect 173126 575048 173131 575104
rect 142110 575046 173131 575048
rect 254932 575046 291884 575106
rect 173065 575043 173131 575046
rect 291878 575044 291884 575046
rect 291948 575044 291954 575108
rect 376937 575106 377003 575109
rect 374900 575104 377003 575106
rect 374900 575048 376942 575104
rect 376998 575048 377003 575104
rect 374900 575046 377003 575048
rect 376937 575043 377003 575046
rect 53465 574562 53531 574565
rect 171133 574562 171199 574565
rect 255221 574562 255287 574565
rect 53465 574560 60076 574562
rect 53465 574504 53470 574560
rect 53526 574504 60076 574560
rect 53465 574502 60076 574504
rect 171133 574560 180044 574562
rect 171133 574504 171138 574560
rect 171194 574504 180044 574560
rect 171133 574502 180044 574504
rect 255221 574560 300196 574562
rect 255221 574504 255226 574560
rect 255282 574504 300196 574560
rect 255221 574502 300196 574504
rect 53465 574499 53531 574502
rect 171133 574499 171199 574502
rect 255221 574499 255287 574502
rect 134934 574366 142170 574426
rect 134934 574260 134994 574366
rect 142110 574290 142170 574366
rect 174445 574290 174511 574293
rect 285438 574290 285444 574292
rect 142110 574288 174511 574290
rect 142110 574232 174450 574288
rect 174506 574232 174511 574288
rect 142110 574230 174511 574232
rect 254932 574230 285444 574290
rect 174445 574227 174511 574230
rect 285438 574228 285444 574230
rect 285508 574228 285514 574292
rect 382222 574290 382228 574292
rect 374900 574230 382228 574290
rect 382222 574228 382228 574230
rect 382292 574228 382298 574292
rect 55029 573474 55095 573477
rect 169109 573474 169175 573477
rect 378041 573474 378107 573477
rect 55029 573472 60076 573474
rect 55029 573416 55034 573472
rect 55090 573416 60076 573472
rect 169109 573472 180044 573474
rect 55029 573414 60076 573416
rect 55029 573411 55095 573414
rect 134934 573338 134994 573444
rect 169109 573416 169114 573472
rect 169170 573416 180044 573472
rect 169109 573414 180044 573416
rect 169109 573411 169175 573414
rect 178493 573338 178559 573341
rect 134934 573336 178559 573338
rect 134934 573280 178498 573336
rect 178554 573280 178559 573336
rect 134934 573278 178559 573280
rect 178493 573275 178559 573278
rect 254902 572930 254962 573444
rect 296670 573414 300196 573474
rect 374900 573472 378107 573474
rect 374900 573416 378046 573472
rect 378102 573416 378107 573472
rect 374900 573414 378107 573416
rect 255129 573202 255195 573205
rect 296670 573202 296730 573414
rect 378041 573411 378107 573414
rect 255129 573200 296730 573202
rect 255129 573144 255134 573200
rect 255190 573144 296730 573200
rect 255129 573142 296730 573144
rect 255129 573139 255195 573142
rect 257521 572930 257587 572933
rect 254902 572928 257587 572930
rect 254902 572872 257526 572928
rect 257582 572872 257587 572928
rect 254902 572870 257587 572872
rect 257521 572867 257587 572870
rect 256734 572732 256740 572796
rect 256804 572794 256810 572796
rect 257797 572794 257863 572797
rect 256804 572792 257863 572794
rect 256804 572736 257802 572792
rect 257858 572736 257863 572792
rect 256804 572734 257863 572736
rect 256804 572732 256810 572734
rect 257797 572731 257863 572734
rect 54477 572386 54543 572389
rect 54477 572384 60076 572386
rect 54477 572328 54482 572384
rect 54538 572328 60076 572384
rect 54477 572326 60076 572328
rect 54477 572323 54543 572326
rect 134934 572114 134994 572628
rect 174905 572386 174971 572389
rect 174905 572384 180044 572386
rect 174905 572328 174910 572384
rect 174966 572328 180044 572384
rect 174905 572326 180044 572328
rect 174905 572323 174971 572326
rect 137093 572114 137159 572117
rect 134934 572112 137159 572114
rect 134934 572056 137098 572112
rect 137154 572056 137159 572112
rect 134934 572054 137159 572056
rect 137093 572051 137159 572054
rect 254902 571978 254962 572628
rect 257102 572596 257108 572660
rect 257172 572658 257178 572660
rect 257889 572658 257955 572661
rect 378041 572658 378107 572661
rect 257172 572656 257955 572658
rect 257172 572600 257894 572656
rect 257950 572600 257955 572656
rect 257172 572598 257955 572600
rect 374900 572656 378107 572658
rect 374900 572600 378046 572656
rect 378102 572600 378107 572656
rect 374900 572598 378107 572600
rect 257172 572596 257178 572598
rect 257889 572595 257955 572598
rect 378041 572595 378107 572598
rect 291745 572386 291811 572389
rect 291745 572384 300196 572386
rect 291745 572328 291750 572384
rect 291806 572328 300196 572384
rect 291745 572326 300196 572328
rect 291745 572323 291811 572326
rect 134934 571918 142170 571978
rect 254902 571918 257354 571978
rect 134934 571812 134994 571918
rect 142110 571842 142170 571918
rect 162209 571842 162275 571845
rect 257102 571842 257108 571844
rect 142110 571840 162275 571842
rect 142110 571784 162214 571840
rect 162270 571784 162275 571840
rect 142110 571782 162275 571784
rect 254932 571782 257108 571842
rect 162209 571779 162275 571782
rect 257102 571780 257108 571782
rect 257172 571780 257178 571844
rect 257294 571842 257354 571918
rect 257613 571842 257679 571845
rect 378041 571842 378107 571845
rect 257294 571840 257679 571842
rect 257294 571784 257618 571840
rect 257674 571784 257679 571840
rect 257294 571782 257679 571784
rect 374900 571840 378107 571842
rect 374900 571784 378046 571840
rect 378102 571784 378107 571840
rect 374900 571782 378107 571784
rect 257613 571779 257679 571782
rect 378041 571779 378107 571782
rect 58617 571298 58683 571301
rect 58617 571296 60076 571298
rect 58617 571240 58622 571296
rect 58678 571240 60076 571296
rect 58617 571238 60076 571240
rect 58617 571235 58683 571238
rect 166574 571236 166580 571300
rect 166644 571298 166650 571300
rect 166644 571238 180044 571298
rect 166644 571236 166650 571238
rect 286542 571236 286548 571300
rect 286612 571298 286618 571300
rect 286612 571238 300196 571298
rect 286612 571236 286618 571238
rect 299105 571162 299171 571165
rect 299238 571162 299244 571164
rect 134934 571102 142170 571162
rect 134934 570996 134994 571102
rect 142110 571026 142170 571102
rect 299105 571160 299244 571162
rect 299105 571104 299110 571160
rect 299166 571104 299244 571160
rect 299105 571102 299244 571104
rect 299105 571099 299171 571102
rect 299238 571100 299244 571102
rect 299308 571100 299314 571164
rect 175549 571026 175615 571029
rect 256918 571026 256924 571028
rect 142110 571024 175615 571026
rect 142110 570968 175554 571024
rect 175610 570968 175615 571024
rect 142110 570966 175615 570968
rect 254932 570966 256924 571026
rect 175549 570963 175615 570966
rect 256918 570964 256924 570966
rect 256988 570964 256994 571028
rect 374870 570346 374930 570996
rect 378041 570346 378107 570349
rect 134934 570286 142170 570346
rect 374870 570344 378107 570346
rect 374870 570288 378046 570344
rect 378102 570288 378107 570344
rect 374870 570286 378107 570288
rect 55949 570210 56015 570213
rect 55949 570208 60076 570210
rect 55949 570152 55954 570208
rect 56010 570152 60076 570208
rect 134934 570180 134994 570286
rect 142110 570210 142170 570286
rect 378041 570283 378107 570286
rect 174997 570210 175063 570213
rect 289721 570210 289787 570213
rect 142110 570208 175063 570210
rect 55949 570150 60076 570152
rect 142110 570152 175002 570208
rect 175058 570152 175063 570208
rect 142110 570150 175063 570152
rect 55949 570147 56015 570150
rect 174997 570147 175063 570150
rect 175230 570150 180044 570210
rect 289721 570208 300196 570210
rect 171542 570012 171548 570076
rect 171612 570074 171618 570076
rect 175230 570074 175290 570150
rect 171612 570014 175290 570074
rect 254902 570074 254962 570180
rect 289721 570152 289726 570208
rect 289782 570152 300196 570208
rect 289721 570150 300196 570152
rect 289721 570147 289787 570150
rect 299238 570074 299244 570076
rect 254902 570014 299244 570074
rect 171612 570012 171618 570014
rect 299238 570012 299244 570014
rect 299308 570012 299314 570076
rect 374686 569941 374746 570180
rect 165061 569938 165127 569941
rect 173801 569938 173867 569941
rect 165061 569936 173867 569938
rect 165061 569880 165066 569936
rect 165122 569880 173806 569936
rect 173862 569880 173867 569936
rect 165061 569878 173867 569880
rect 165061 569875 165127 569878
rect 173801 569875 173867 569878
rect 177113 569938 177179 569941
rect 294873 569940 294939 569941
rect 177246 569938 177252 569940
rect 177113 569936 177252 569938
rect 177113 569880 177118 569936
rect 177174 569880 177252 569936
rect 177113 569878 177252 569880
rect 177113 569875 177179 569878
rect 177246 569876 177252 569878
rect 177316 569876 177322 569940
rect 294822 569938 294828 569940
rect 294782 569878 294828 569938
rect 294892 569936 294939 569940
rect 294934 569880 294939 569936
rect 294822 569876 294828 569878
rect 294892 569876 294939 569880
rect 374686 569936 374795 569941
rect 374686 569880 374734 569936
rect 374790 569880 374795 569936
rect 374686 569878 374795 569880
rect 294873 569875 294939 569876
rect 374729 569875 374795 569878
rect 134934 569470 142170 569530
rect 134934 569364 134994 569470
rect 142110 569394 142170 569470
rect 166165 569394 166231 569397
rect 295006 569394 295012 569396
rect 142110 569392 166231 569394
rect 142110 569336 166170 569392
rect 166226 569336 166231 569392
rect 142110 569334 166231 569336
rect 254932 569334 295012 569394
rect 166165 569331 166231 569334
rect 295006 569332 295012 569334
rect 295076 569332 295082 569396
rect 377029 569394 377095 569397
rect 374900 569392 377095 569394
rect 374900 569336 377034 569392
rect 377090 569336 377095 569392
rect 374900 569334 377095 569336
rect 377029 569331 377095 569334
rect 256509 569258 256575 569261
rect 292205 569258 292271 569261
rect 256509 569256 292271 569258
rect 256509 569200 256514 569256
rect 256570 569200 292210 569256
rect 292266 569200 292271 569256
rect 256509 569198 292271 569200
rect 256509 569195 256575 569198
rect 292205 569195 292271 569198
rect 59629 569122 59695 569125
rect 59629 569120 60076 569122
rect 59629 569064 59634 569120
rect 59690 569064 60076 569120
rect 59629 569062 60076 569064
rect 59629 569059 59695 569062
rect 177246 569060 177252 569124
rect 177316 569122 177322 569124
rect 297725 569122 297791 569125
rect 177316 569062 180044 569122
rect 297725 569120 300196 569122
rect 297725 569064 297730 569120
rect 297786 569064 300196 569120
rect 297725 569062 300196 569064
rect 177316 569060 177322 569062
rect 297725 569059 297791 569062
rect 178401 568578 178467 568581
rect 142110 568576 178467 568578
rect 134934 568442 134994 568548
rect 142110 568520 178406 568576
rect 178462 568520 178467 568576
rect 142110 568518 178467 568520
rect 254932 568518 277410 568578
rect 142110 568442 142170 568518
rect 178401 568515 178467 568518
rect 134934 568382 142170 568442
rect 277350 568306 277410 568518
rect 292614 568516 292620 568580
rect 292684 568578 292690 568580
rect 293769 568578 293835 568581
rect 377765 568578 377831 568581
rect 292684 568576 293835 568578
rect 292684 568520 293774 568576
rect 293830 568520 293835 568576
rect 292684 568518 293835 568520
rect 374900 568576 377831 568578
rect 374900 568520 377770 568576
rect 377826 568520 377831 568576
rect 374900 568518 377831 568520
rect 292684 568516 292690 568518
rect 293769 568515 293835 568518
rect 377765 568515 377831 568518
rect 292982 568306 292988 568308
rect 277350 568246 292988 568306
rect 292982 568244 292988 568246
rect 293052 568244 293058 568308
rect 56501 568034 56567 568037
rect 56501 568032 60076 568034
rect 56501 567976 56506 568032
rect 56562 567976 60076 568032
rect 56501 567974 60076 567976
rect 56501 567971 56567 567974
rect 175038 567972 175044 568036
rect 175108 568034 175114 568036
rect 289445 568034 289511 568037
rect 175108 567974 180044 568034
rect 289445 568032 300196 568034
rect 289445 567976 289450 568032
rect 289506 567976 300196 568032
rect 289445 567974 300196 567976
rect 175108 567972 175114 567974
rect 289445 567971 289511 567974
rect 296529 567490 296595 567493
rect 296662 567490 296668 567492
rect 296529 567488 296668 567490
rect 296529 567432 296534 567488
rect 296590 567432 296668 567488
rect 296529 567430 296668 567432
rect 296529 567427 296595 567430
rect 296662 567428 296668 567430
rect 296732 567428 296738 567492
rect 296529 567082 296595 567085
rect 296662 567082 296668 567084
rect 296529 567080 296668 567082
rect -960 566946 480 567036
rect 296529 567024 296534 567080
rect 296590 567024 296668 567080
rect 296529 567022 296668 567024
rect 296529 567019 296595 567022
rect 296662 567020 296668 567022
rect 296732 567020 296738 567084
rect 2814 566946 2820 566948
rect -960 566886 2820 566946
rect -960 566796 480 566886
rect 2814 566884 2820 566886
rect 2884 566884 2890 566948
rect 292297 566946 292363 566949
rect 292297 566944 299674 566946
rect 292297 566888 292302 566944
rect 292358 566888 299674 566944
rect 292297 566886 299674 566888
rect 292297 566883 292363 566886
rect 59494 566818 60076 566878
rect 55765 566810 55831 566813
rect 59494 566810 59554 566818
rect 179822 566816 179828 566880
rect 179892 566878 179898 566880
rect 299614 566878 299674 566886
rect 179892 566818 180044 566878
rect 299614 566818 300196 566878
rect 179892 566816 179898 566818
rect 55765 566808 59554 566810
rect 55765 566752 55770 566808
rect 55826 566752 59554 566808
rect 55765 566750 59554 566752
rect 55765 566747 55831 566750
rect 59261 565858 59327 565861
rect 59261 565856 59922 565858
rect 59261 565800 59266 565856
rect 59322 565800 59922 565856
rect 59261 565798 59922 565800
rect 59261 565795 59327 565798
rect 59862 565790 59922 565798
rect 179454 565796 179460 565860
rect 179524 565858 179530 565860
rect 293861 565858 293927 565861
rect 179524 565798 180044 565858
rect 293861 565856 300042 565858
rect 293861 565800 293866 565856
rect 293922 565800 300042 565856
rect 293861 565798 300042 565800
rect 179524 565796 179530 565798
rect 293861 565795 293927 565798
rect 299982 565790 300042 565798
rect 59862 565730 60076 565790
rect 299982 565730 300196 565790
rect 176510 564708 176516 564772
rect 176580 564770 176586 564772
rect 176580 564710 180044 564770
rect 176580 564708 176586 564710
rect 289118 564708 289124 564772
rect 289188 564770 289194 564772
rect 289188 564710 299674 564770
rect 289188 564708 289194 564710
rect 299614 564702 299674 564710
rect 59494 564642 60076 564702
rect 299614 564642 300196 564702
rect 58341 564634 58407 564637
rect 59494 564634 59554 564642
rect 58341 564632 59554 564634
rect 58341 564576 58346 564632
rect 58402 564576 59554 564632
rect 58341 564574 59554 564576
rect 58341 564571 58407 564574
rect 288382 564436 288388 564500
rect 288452 564498 288458 564500
rect 289629 564498 289695 564501
rect 288452 564496 289695 564498
rect 288452 564440 289634 564496
rect 289690 564440 289695 564496
rect 288452 564438 289695 564440
rect 288452 564436 288458 564438
rect 289629 564435 289695 564438
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect 288934 563620 288940 563684
rect 289004 563682 289010 563684
rect 289004 563622 299674 563682
rect 289004 563620 289010 563622
rect 179689 563614 179755 563617
rect 299614 563614 299674 563622
rect 59494 563554 60076 563614
rect 179689 563612 180044 563614
rect 179689 563556 179694 563612
rect 179750 563556 180044 563612
rect 179689 563554 180044 563556
rect 299614 563554 300196 563614
rect 57697 563546 57763 563549
rect 59494 563546 59554 563554
rect 179689 563551 179755 563554
rect 57697 563544 59554 563546
rect 57697 563488 57702 563544
rect 57758 563488 59554 563544
rect 57697 563486 59554 563488
rect 57697 563483 57763 563486
rect 179597 563138 179663 563141
rect 179822 563138 179828 563140
rect 179597 563136 179828 563138
rect 179597 563080 179602 563136
rect 179658 563080 179828 563136
rect 179597 563078 179828 563080
rect 179597 563075 179663 563078
rect 179822 563076 179828 563078
rect 179892 563076 179898 563140
rect 288566 563076 288572 563140
rect 288636 563138 288642 563140
rect 289537 563138 289603 563141
rect 288636 563136 289603 563138
rect 288636 563080 289542 563136
rect 289598 563080 289603 563136
rect 288636 563078 289603 563080
rect 288636 563076 288642 563078
rect 289537 563075 289603 563078
rect 292246 562532 292252 562596
rect 292316 562594 292322 562596
rect 292316 562534 299674 562594
rect 292316 562532 292322 562534
rect 59494 562466 60076 562526
rect 57145 562458 57211 562461
rect 59494 562458 59554 562466
rect 180374 562464 180380 562528
rect 180444 562464 180450 562528
rect 299614 562526 299674 562534
rect 299614 562466 300196 562526
rect 57145 562456 59554 562458
rect 57145 562400 57150 562456
rect 57206 562400 59554 562456
rect 57145 562398 59554 562400
rect 57145 562395 57211 562398
rect 291142 562260 291148 562324
rect 291212 562322 291218 562324
rect 292481 562322 292547 562325
rect 291212 562320 292547 562322
rect 291212 562264 292486 562320
rect 292542 562264 292547 562320
rect 291212 562262 292547 562264
rect 291212 562260 291218 562262
rect 292481 562259 292547 562262
rect 259085 561778 259151 561781
rect 299013 561778 299079 561781
rect 259085 561776 299079 561778
rect 259085 561720 259090 561776
rect 259146 561720 299018 561776
rect 299074 561720 299079 561776
rect 259085 561718 299079 561720
rect 259085 561715 259151 561718
rect 299013 561715 299079 561718
rect 172646 561580 172652 561644
rect 172716 561642 172722 561644
rect 172881 561642 172947 561645
rect 172716 561640 172947 561642
rect 172716 561584 172886 561640
rect 172942 561584 172947 561640
rect 172716 561582 172947 561584
rect 172716 561580 172722 561582
rect 172881 561579 172947 561582
rect 59537 561438 59603 561441
rect 59537 561436 60076 561438
rect 59537 561380 59542 561436
rect 59598 561380 60076 561436
rect 59537 561378 60076 561380
rect 59537 561375 59603 561378
rect 180558 561376 180564 561440
rect 180628 561376 180634 561440
rect 299614 561378 300196 561438
rect 297909 561370 297975 561373
rect 299614 561370 299674 561378
rect 297909 561368 299674 561370
rect 297909 561312 297914 561368
rect 297970 561312 299674 561368
rect 297909 561310 299674 561312
rect 297909 561307 297975 561310
rect 255814 560628 255820 560692
rect 255884 560690 255890 560692
rect 255884 560630 299674 560690
rect 255884 560628 255890 560630
rect 49509 560554 49575 560557
rect 162393 560554 162459 560557
rect 49509 560552 162459 560554
rect 49509 560496 49514 560552
rect 49570 560496 162398 560552
rect 162454 560496 162459 560552
rect 49509 560494 162459 560496
rect 49509 560491 49575 560494
rect 162393 560491 162459 560494
rect 172973 560554 173039 560557
rect 172973 560552 233434 560554
rect 172973 560496 172978 560552
rect 173034 560496 233434 560552
rect 172973 560494 233434 560496
rect 172973 560491 173039 560494
rect 177982 560356 177988 560420
rect 178052 560418 178058 560420
rect 178052 560358 178970 560418
rect 178052 560356 178058 560358
rect 57605 560284 57671 560285
rect 57605 560282 57652 560284
rect 57560 560280 57652 560282
rect 57560 560224 57610 560280
rect 57560 560222 57652 560224
rect 57605 560220 57652 560222
rect 57716 560220 57722 560284
rect 59118 560220 59124 560284
rect 59188 560282 59194 560284
rect 60641 560282 60707 560285
rect 166809 560284 166875 560285
rect 166758 560282 166764 560284
rect 59188 560280 60707 560282
rect 59188 560224 60646 560280
rect 60702 560224 60707 560280
rect 59188 560222 60707 560224
rect 166718 560222 166764 560282
rect 166828 560280 166875 560284
rect 166870 560224 166875 560280
rect 59188 560220 59194 560222
rect 57605 560219 57671 560220
rect 60641 560219 60707 560222
rect 166758 560220 166764 560222
rect 166828 560220 166875 560224
rect 175222 560220 175228 560284
rect 175292 560282 175298 560284
rect 175457 560282 175523 560285
rect 175292 560280 175523 560282
rect 175292 560224 175462 560280
rect 175518 560224 175523 560280
rect 175292 560222 175523 560224
rect 175292 560220 175298 560222
rect 166809 560219 166875 560220
rect 175457 560219 175523 560222
rect 45093 560146 45159 560149
rect 178910 560146 178970 560358
rect 233374 560285 233434 560494
rect 255078 560492 255084 560556
rect 255148 560554 255154 560556
rect 298737 560554 298803 560557
rect 255148 560552 298803 560554
rect 255148 560496 298742 560552
rect 298798 560496 298803 560552
rect 255148 560494 298803 560496
rect 299614 560554 299674 560630
rect 302233 560554 302299 560557
rect 299614 560552 302299 560554
rect 299614 560496 302238 560552
rect 302294 560496 302299 560552
rect 299614 560494 302299 560496
rect 255148 560492 255154 560494
rect 298737 560491 298803 560494
rect 302233 560491 302299 560494
rect 253013 560418 253079 560421
rect 529933 560418 529999 560421
rect 253013 560416 529999 560418
rect 253013 560360 253018 560416
rect 253074 560360 529938 560416
rect 529994 560360 529999 560416
rect 253013 560358 529999 560360
rect 253013 560355 253079 560358
rect 529933 560355 529999 560358
rect 233374 560282 233483 560285
rect 289261 560282 289327 560285
rect 233374 560280 289327 560282
rect 233374 560224 233422 560280
rect 233478 560224 289266 560280
rect 289322 560224 289327 560280
rect 233374 560222 289327 560224
rect 233417 560219 233483 560222
rect 289261 560219 289327 560222
rect 299013 560282 299079 560285
rect 305545 560282 305611 560285
rect 299013 560280 305611 560282
rect 299013 560224 299018 560280
rect 299074 560224 305550 560280
rect 305606 560224 305611 560280
rect 299013 560222 305611 560224
rect 299013 560219 299079 560222
rect 305545 560219 305611 560222
rect 179045 560146 179111 560149
rect 45093 560144 157350 560146
rect 45093 560088 45098 560144
rect 45154 560088 157350 560144
rect 45093 560086 157350 560088
rect 178910 560144 179111 560146
rect 178910 560088 179050 560144
rect 179106 560088 179111 560144
rect 178910 560086 179111 560088
rect 45093 560083 45159 560086
rect 157290 560010 157350 560086
rect 179045 560083 179111 560086
rect 216903 560146 216969 560149
rect 233693 560146 233759 560149
rect 248597 560146 248663 560149
rect 294597 560146 294663 560149
rect 216903 560144 233759 560146
rect 216903 560088 216908 560144
rect 216964 560088 233698 560144
rect 233754 560088 233759 560144
rect 216903 560086 233759 560088
rect 216903 560083 216969 560086
rect 233693 560083 233759 560086
rect 238710 560144 248663 560146
rect 238710 560088 248602 560144
rect 248658 560088 248663 560144
rect 238710 560086 248663 560088
rect 171041 560010 171107 560013
rect 238710 560010 238770 560086
rect 248597 560083 248663 560086
rect 258030 560144 294663 560146
rect 258030 560088 294602 560144
rect 294658 560088 294663 560144
rect 258030 560086 294663 560088
rect 157290 559950 167378 560010
rect 46749 559874 46815 559877
rect 162301 559874 162367 559877
rect 46749 559872 162367 559874
rect 46749 559816 46754 559872
rect 46810 559816 162306 559872
rect 162362 559816 162367 559872
rect 46749 559814 162367 559816
rect 167318 559874 167378 559950
rect 171041 560008 238770 560010
rect 171041 559952 171046 560008
rect 171102 559952 238770 560008
rect 171041 559950 238770 559952
rect 245469 560010 245535 560013
rect 258030 560010 258090 560086
rect 294597 560083 294663 560086
rect 245469 560008 258090 560010
rect 245469 559952 245474 560008
rect 245530 559952 258090 560008
rect 245469 559950 258090 559952
rect 171041 559947 171107 559950
rect 245469 559947 245535 559950
rect 169385 559874 169451 559877
rect 244457 559874 244523 559877
rect 258993 559874 259059 559877
rect 167318 559872 259059 559874
rect 167318 559816 169390 559872
rect 169446 559816 244462 559872
rect 244518 559816 258998 559872
rect 259054 559816 259059 559872
rect 167318 559814 259059 559816
rect 46749 559811 46815 559814
rect 162301 559811 162367 559814
rect 169385 559811 169451 559814
rect 244457 559811 244523 559814
rect 258993 559811 259059 559814
rect 294965 559874 295031 559877
rect 534257 559874 534323 559877
rect 294965 559872 534323 559874
rect 294965 559816 294970 559872
rect 295026 559816 534262 559872
rect 534318 559816 534323 559872
rect 294965 559814 534323 559816
rect 294965 559811 295031 559814
rect 534257 559811 534323 559814
rect 58801 559738 58867 559741
rect 169845 559738 169911 559741
rect 58801 559736 169911 559738
rect 58801 559680 58806 559736
rect 58862 559680 169850 559736
rect 169906 559680 169911 559736
rect 58801 559678 169911 559680
rect 58801 559675 58867 559678
rect 169845 559675 169911 559678
rect 170949 559738 171015 559741
rect 246389 559738 246455 559741
rect 170949 559736 246455 559738
rect 170949 559680 170954 559736
rect 171010 559680 246394 559736
rect 246450 559680 246455 559736
rect 170949 559678 246455 559680
rect 170949 559675 171015 559678
rect 246389 559675 246455 559678
rect 257705 559738 257771 559741
rect 501413 559738 501479 559741
rect 257705 559736 501479 559738
rect 257705 559680 257710 559736
rect 257766 559680 501418 559736
rect 501474 559680 501479 559736
rect 257705 559678 501479 559680
rect 257705 559675 257771 559678
rect 501413 559675 501479 559678
rect 166165 559602 166231 559605
rect 427629 559602 427695 559605
rect 166165 559600 427695 559602
rect 166165 559544 166170 559600
rect 166226 559544 427634 559600
rect 427690 559544 427695 559600
rect 166165 559542 427695 559544
rect 166165 559539 166231 559542
rect 427629 559539 427695 559542
rect 58750 559404 58756 559468
rect 58820 559466 58826 559468
rect 169753 559466 169819 559469
rect 58820 559464 169819 559466
rect 58820 559408 169758 559464
rect 169814 559408 169819 559464
rect 58820 559406 169819 559408
rect 58820 559404 58826 559406
rect 169753 559403 169819 559406
rect 176561 559466 176627 559469
rect 240133 559466 240199 559469
rect 176561 559464 240199 559466
rect 176561 559408 176566 559464
rect 176622 559408 240138 559464
rect 240194 559408 240199 559464
rect 176561 559406 240199 559408
rect 176561 559403 176627 559406
rect 240133 559403 240199 559406
rect 55121 559330 55187 559333
rect 172145 559330 172211 559333
rect 172973 559330 173039 559333
rect 55121 559328 173039 559330
rect 55121 559272 55126 559328
rect 55182 559272 172150 559328
rect 172206 559272 172978 559328
rect 173034 559272 173039 559328
rect 55121 559270 173039 559272
rect 55121 559267 55187 559270
rect 172145 559267 172211 559270
rect 172973 559267 173039 559270
rect 176377 559330 176443 559333
rect 237373 559330 237439 559333
rect 255865 559330 255931 559333
rect 176377 559328 255931 559330
rect 176377 559272 176382 559328
rect 176438 559272 237378 559328
rect 237434 559272 255870 559328
rect 255926 559272 255931 559328
rect 176377 559270 255931 559272
rect 176377 559267 176443 559270
rect 237373 559267 237439 559270
rect 255865 559267 255931 559270
rect 58709 559194 58775 559197
rect 216673 559194 216739 559197
rect 58709 559192 216739 559194
rect 58709 559136 58714 559192
rect 58770 559136 216678 559192
rect 216734 559136 216739 559192
rect 58709 559134 216739 559136
rect 58709 559131 58775 559134
rect 216673 559131 216739 559134
rect 240409 559194 240475 559197
rect 256417 559194 256483 559197
rect 240409 559192 256483 559194
rect 240409 559136 240414 559192
rect 240470 559136 256422 559192
rect 256478 559136 256483 559192
rect 240409 559134 256483 559136
rect 240409 559131 240475 559134
rect 256417 559131 256483 559134
rect 59854 558996 59860 559060
rect 59924 559058 59930 559060
rect 175733 559058 175799 559061
rect 59924 559056 175799 559058
rect 59924 559000 175738 559056
rect 175794 559000 175799 559056
rect 59924 558998 175799 559000
rect 59924 558996 59930 558998
rect 175733 558995 175799 558998
rect 252553 559058 252619 559061
rect 260281 559058 260347 559061
rect 252553 559056 260347 559058
rect 252553 559000 252558 559056
rect 252614 559000 260286 559056
rect 260342 559000 260347 559056
rect 252553 558998 260347 559000
rect 252553 558995 252619 558998
rect 260281 558995 260347 558998
rect 511993 559058 512059 559061
rect 512126 559058 512132 559060
rect 511993 559056 512132 559058
rect 511993 559000 511998 559056
rect 512054 559000 512132 559056
rect 511993 558998 512132 559000
rect 511993 558995 512059 558998
rect 512126 558996 512132 558998
rect 512196 558996 512202 559060
rect 173934 558860 173940 558924
rect 174004 558922 174010 558924
rect 174261 558922 174327 558925
rect 180609 558924 180675 558925
rect 180558 558922 180564 558924
rect 174004 558920 174327 558922
rect 174004 558864 174266 558920
rect 174322 558864 174327 558920
rect 174004 558862 174327 558864
rect 180518 558862 180564 558922
rect 180628 558920 180675 558924
rect 180670 558864 180675 558920
rect 174004 558860 174010 558862
rect 174261 558859 174327 558862
rect 180558 558860 180564 558862
rect 180628 558860 180675 558864
rect 180609 558859 180675 558860
rect 246389 558922 246455 558925
rect 255957 558922 256023 558925
rect 246389 558920 256023 558922
rect 246389 558864 246394 558920
rect 246450 558864 255962 558920
rect 256018 558864 256023 558920
rect 246389 558862 256023 558864
rect 246389 558859 246455 558862
rect 255957 558859 256023 558862
rect 54477 558786 54543 558789
rect 54477 558784 171150 558786
rect 54477 558728 54482 558784
rect 54538 558728 171150 558784
rect 54477 558726 171150 558728
rect 54477 558723 54543 558726
rect 45369 558650 45435 558653
rect 162577 558650 162643 558653
rect 45369 558648 162643 558650
rect 45369 558592 45374 558648
rect 45430 558592 162582 558648
rect 162638 558592 162643 558648
rect 45369 558590 162643 558592
rect 45369 558587 45435 558590
rect 162577 558587 162643 558590
rect 54569 558514 54635 558517
rect 168281 558514 168347 558517
rect 54569 558512 168347 558514
rect 54569 558456 54574 558512
rect 54630 558456 168286 558512
rect 168342 558456 168347 558512
rect 54569 558454 168347 558456
rect 171090 558514 171150 558726
rect 180374 558724 180380 558788
rect 180444 558786 180450 558788
rect 180701 558786 180767 558789
rect 180444 558784 180767 558786
rect 180444 558728 180706 558784
rect 180762 558728 180767 558784
rect 180444 558726 180767 558728
rect 180444 558724 180450 558726
rect 180701 558723 180767 558726
rect 243445 558786 243511 558789
rect 292021 558786 292087 558789
rect 243445 558784 292087 558786
rect 243445 558728 243450 558784
rect 243506 558728 292026 558784
rect 292082 558728 292087 558784
rect 243445 558726 292087 558728
rect 243445 558723 243511 558726
rect 292021 558723 292087 558726
rect 292205 558786 292271 558789
rect 322749 558786 322815 558789
rect 292205 558784 322815 558786
rect 292205 558728 292210 558784
rect 292266 558728 322754 558784
rect 322810 558728 322815 558784
rect 292205 558726 322815 558728
rect 292205 558723 292271 558726
rect 322749 558723 322815 558726
rect 172973 558650 173039 558653
rect 236361 558650 236427 558653
rect 292389 558650 292455 558653
rect 172973 558648 292455 558650
rect 172973 558592 172978 558648
rect 173034 558592 236366 558648
rect 236422 558592 292394 558648
rect 292450 558592 292455 558648
rect 172973 558590 292455 558592
rect 172973 558587 173039 558590
rect 236361 558587 236427 558590
rect 292389 558587 292455 558590
rect 174905 558514 174971 558517
rect 226241 558514 226307 558517
rect 291745 558514 291811 558517
rect 171090 558512 291811 558514
rect 171090 558456 174910 558512
rect 174966 558456 226246 558512
rect 226302 558456 291750 558512
rect 291806 558456 291811 558512
rect 171090 558454 291811 558456
rect 54569 558451 54635 558454
rect 168281 558451 168347 558454
rect 174905 558451 174971 558454
rect 226241 558451 226307 558454
rect 291745 558451 291811 558454
rect 295006 558452 295012 558516
rect 295076 558514 295082 558516
rect 523166 558514 523172 558516
rect 295076 558454 523172 558514
rect 295076 558452 295082 558454
rect 523166 558452 523172 558454
rect 523236 558452 523242 558516
rect 175181 558378 175247 558381
rect 238385 558378 238451 558381
rect 256325 558378 256391 558381
rect 175181 558376 256391 558378
rect 175181 558320 175186 558376
rect 175242 558320 238390 558376
rect 238446 558320 256330 558376
rect 256386 558320 256391 558376
rect 175181 558318 256391 558320
rect 175181 558315 175247 558318
rect 238385 558315 238451 558318
rect 256325 558315 256391 558318
rect 257521 558378 257587 558381
rect 515397 558378 515463 558381
rect 257521 558376 515463 558378
rect 257521 558320 257526 558376
rect 257582 558320 515402 558376
rect 515458 558320 515463 558376
rect 257521 558318 515463 558320
rect 257521 558315 257587 558318
rect 515397 558315 515463 558318
rect 39481 558242 39547 558245
rect 56041 558242 56107 558245
rect 39481 558240 56107 558242
rect 39481 558184 39486 558240
rect 39542 558184 56046 558240
rect 56102 558184 56107 558240
rect 39481 558182 56107 558184
rect 39481 558179 39547 558182
rect 56041 558179 56107 558182
rect 64505 558242 64571 558245
rect 68277 558242 68343 558245
rect 64505 558240 68343 558242
rect 64505 558184 64510 558240
rect 64566 558184 68282 558240
rect 68338 558184 68343 558240
rect 64505 558182 68343 558184
rect 64505 558179 64571 558182
rect 68277 558179 68343 558182
rect 169569 558242 169635 558245
rect 243445 558242 243511 558245
rect 169569 558240 243511 558242
rect 169569 558184 169574 558240
rect 169630 558184 243450 558240
rect 243506 558184 243511 558240
rect 169569 558182 243511 558184
rect 169569 558179 169635 558182
rect 243445 558179 243511 558182
rect 256918 558180 256924 558244
rect 256988 558242 256994 558244
rect 515254 558242 515260 558244
rect 256988 558182 515260 558242
rect 256988 558180 256994 558182
rect 515254 558180 515260 558182
rect 515324 558180 515330 558244
rect 43437 558106 43503 558109
rect 53833 558106 53899 558109
rect 43437 558104 53899 558106
rect 43437 558048 43442 558104
rect 43498 558048 53838 558104
rect 53894 558048 53899 558104
rect 43437 558046 53899 558048
rect 43437 558043 43503 558046
rect 53833 558043 53899 558046
rect 58801 558106 58867 558109
rect 63585 558106 63651 558109
rect 58801 558104 63651 558106
rect 58801 558048 58806 558104
rect 58862 558048 63590 558104
rect 63646 558048 63651 558104
rect 58801 558046 63651 558048
rect 58801 558043 58867 558046
rect 63585 558043 63651 558046
rect 231209 558106 231275 558109
rect 255037 558106 255103 558109
rect 231209 558104 255103 558106
rect 231209 558048 231214 558104
rect 231270 558048 255042 558104
rect 255098 558048 255103 558104
rect 231209 558046 255103 558048
rect 231209 558043 231275 558046
rect 255037 558043 255103 558046
rect 42057 557970 42123 557973
rect 53925 557970 53991 557973
rect 42057 557968 53991 557970
rect 42057 557912 42062 557968
rect 42118 557912 53930 557968
rect 53986 557912 53991 557968
rect 42057 557910 53991 557912
rect 42057 557907 42123 557910
rect 53925 557907 53991 557910
rect 56041 557970 56107 557973
rect 252461 557970 252527 557973
rect 56041 557968 252527 557970
rect 56041 557912 56046 557968
rect 56102 557912 252466 557968
rect 252522 557912 252527 557968
rect 56041 557910 252527 557912
rect 56041 557907 56107 557910
rect 252461 557907 252527 557910
rect 36629 557834 36695 557837
rect 59261 557834 59327 557837
rect 36629 557832 59327 557834
rect 36629 557776 36634 557832
rect 36690 557776 59266 557832
rect 59322 557776 59327 557832
rect 36629 557774 59327 557776
rect 36629 557771 36695 557774
rect 59261 557771 59327 557774
rect 296529 557834 296595 557837
rect 296662 557834 296668 557836
rect 296529 557832 296668 557834
rect 296529 557776 296534 557832
rect 296590 557776 296668 557832
rect 296529 557774 296668 557776
rect 296529 557771 296595 557774
rect 296662 557772 296668 557774
rect 296732 557772 296738 557836
rect 53598 557636 53604 557700
rect 53668 557698 53674 557700
rect 231761 557698 231827 557701
rect 53668 557696 231827 557698
rect 53668 557640 231766 557696
rect 231822 557640 231827 557696
rect 53668 557638 231827 557640
rect 53668 557636 53674 557638
rect 231761 557635 231827 557638
rect 32806 557500 32812 557564
rect 32876 557562 32882 557564
rect 245653 557562 245719 557565
rect 32876 557560 245719 557562
rect 32876 557504 245658 557560
rect 245714 557504 245719 557560
rect 32876 557502 245719 557504
rect 32876 557500 32882 557502
rect 245653 557499 245719 557502
rect 251541 557562 251607 557565
rect 258165 557562 258231 557565
rect 251541 557560 258231 557562
rect 251541 557504 251546 557560
rect 251602 557504 258170 557560
rect 258226 557504 258231 557560
rect 251541 557502 258231 557504
rect 251541 557499 251607 557502
rect 258165 557499 258231 557502
rect 45185 557426 45251 557429
rect 164969 557426 165035 557429
rect 45185 557424 165035 557426
rect 45185 557368 45190 557424
rect 45246 557368 164974 557424
rect 165030 557368 165035 557424
rect 45185 557366 165035 557368
rect 45185 557363 45251 557366
rect 164969 557363 165035 557366
rect 173525 557426 173591 557429
rect 227713 557426 227779 557429
rect 173525 557424 227779 557426
rect 173525 557368 173530 557424
rect 173586 557368 227718 557424
rect 227774 557368 227779 557424
rect 173525 557366 227779 557368
rect 173525 557363 173591 557366
rect 227713 557363 227779 557366
rect 230197 557426 230263 557429
rect 254945 557426 255011 557429
rect 230197 557424 255011 557426
rect 230197 557368 230202 557424
rect 230258 557368 254950 557424
rect 255006 557368 255011 557424
rect 230197 557366 255011 557368
rect 230197 557363 230263 557366
rect 254945 557363 255011 557366
rect 294638 557364 294644 557428
rect 294708 557426 294714 557428
rect 499062 557426 499068 557428
rect 294708 557366 499068 557426
rect 294708 557364 294714 557366
rect 499062 557364 499068 557366
rect 499132 557364 499138 557428
rect 49233 557290 49299 557293
rect 168097 557290 168163 557293
rect 49233 557288 168163 557290
rect 49233 557232 49238 557288
rect 49294 557232 168102 557288
rect 168158 557232 168163 557288
rect 49233 557230 168163 557232
rect 49233 557227 49299 557230
rect 168097 557227 168163 557230
rect 179965 557290 180031 557293
rect 247125 557290 247191 557293
rect 179965 557288 247191 557290
rect 179965 557232 179970 557288
rect 180026 557232 247130 557288
rect 247186 557232 247191 557288
rect 179965 557230 247191 557232
rect 179965 557227 180031 557230
rect 247125 557227 247191 557230
rect 250529 557290 250595 557293
rect 258809 557290 258875 557293
rect 250529 557288 258875 557290
rect 250529 557232 250534 557288
rect 250590 557232 258814 557288
rect 258870 557232 258875 557288
rect 250529 557230 258875 557232
rect 250529 557227 250595 557230
rect 258809 557227 258875 557230
rect 296529 557290 296595 557293
rect 296662 557290 296668 557292
rect 296529 557288 296668 557290
rect 296529 557232 296534 557288
rect 296590 557232 296668 557288
rect 296529 557230 296668 557232
rect 296529 557227 296595 557230
rect 296662 557228 296668 557230
rect 296732 557228 296738 557292
rect 299054 557228 299060 557292
rect 299124 557290 299130 557292
rect 505134 557290 505140 557292
rect 299124 557230 505140 557290
rect 299124 557228 299130 557230
rect 505134 557228 505140 557230
rect 505204 557228 505210 557292
rect 49325 557154 49391 557157
rect 168005 557154 168071 557157
rect 49325 557152 168071 557154
rect 49325 557096 49330 557152
rect 49386 557096 168010 557152
rect 168066 557096 168071 557152
rect 49325 557094 168071 557096
rect 49325 557091 49391 557094
rect 168005 557091 168071 557094
rect 172421 557154 172487 557157
rect 242433 557154 242499 557157
rect 256049 557154 256115 557157
rect 172421 557152 256115 557154
rect 172421 557096 172426 557152
rect 172482 557096 242438 557152
rect 242494 557096 256054 557152
rect 256110 557096 256115 557152
rect 172421 557094 256115 557096
rect 172421 557091 172487 557094
rect 242433 557091 242499 557094
rect 256049 557091 256115 557094
rect 289302 557092 289308 557156
rect 289372 557154 289378 557156
rect 525374 557154 525380 557156
rect 289372 557094 525380 557154
rect 289372 557092 289378 557094
rect 525374 557092 525380 557094
rect 525444 557092 525450 557156
rect 46565 557018 46631 557021
rect 162761 557018 162827 557021
rect 46565 557016 162827 557018
rect 46565 556960 46570 557016
rect 46626 556960 162766 557016
rect 162822 556960 162827 557016
rect 46565 556958 162827 556960
rect 46565 556955 46631 556958
rect 162761 556955 162827 556958
rect 167729 557018 167795 557021
rect 178125 557018 178191 557021
rect 167729 557016 178191 557018
rect 167729 556960 167734 557016
rect 167790 556960 178130 557016
rect 178186 556960 178191 557016
rect 167729 556958 178191 556960
rect 167729 556955 167795 556958
rect 178125 556955 178191 556958
rect 178585 557018 178651 557021
rect 445845 557018 445911 557021
rect 178585 557016 445911 557018
rect 178585 556960 178590 557016
rect 178646 556960 445850 557016
rect 445906 556960 445911 557016
rect 178585 556958 445911 556960
rect 178585 556955 178651 556958
rect 445845 556955 445911 556958
rect 53465 556882 53531 556885
rect 169201 556882 169267 556885
rect 53465 556880 169267 556882
rect 53465 556824 53470 556880
rect 53526 556824 169206 556880
rect 169262 556824 169267 556880
rect 53465 556822 169267 556824
rect 53465 556819 53531 556822
rect 169201 556819 169267 556822
rect 175825 556882 175891 556885
rect 446857 556882 446923 556885
rect 175825 556880 446923 556882
rect 175825 556824 175830 556880
rect 175886 556824 446862 556880
rect 446918 556824 446923 556880
rect 175825 556822 446923 556824
rect 175825 556819 175891 556822
rect 446857 556819 446923 556822
rect 47945 556746 48011 556749
rect 159725 556746 159791 556749
rect 47945 556744 159791 556746
rect 47945 556688 47950 556744
rect 48006 556688 159730 556744
rect 159786 556688 159791 556744
rect 47945 556686 159791 556688
rect 47945 556683 48011 556686
rect 159725 556683 159791 556686
rect 175089 556746 175155 556749
rect 447869 556746 447935 556749
rect 175089 556744 447935 556746
rect 175089 556688 175094 556744
rect 175150 556688 447874 556744
rect 447930 556688 447935 556744
rect 175089 556686 447935 556688
rect 175089 556683 175155 556686
rect 447869 556683 447935 556686
rect 54661 556610 54727 556613
rect 165245 556610 165311 556613
rect 54661 556608 165311 556610
rect 54661 556552 54666 556608
rect 54722 556552 165250 556608
rect 165306 556552 165311 556608
rect 54661 556550 165311 556552
rect 54661 556547 54727 556550
rect 165245 556547 165311 556550
rect 166625 556610 166691 556613
rect 178033 556610 178099 556613
rect 166625 556608 178099 556610
rect 166625 556552 166630 556608
rect 166686 556552 178038 556608
rect 178094 556552 178099 556608
rect 166625 556550 178099 556552
rect 166625 556547 166691 556550
rect 178033 556547 178099 556550
rect 178718 556548 178724 556612
rect 178788 556610 178794 556612
rect 230381 556610 230447 556613
rect 178788 556608 230447 556610
rect 178788 556552 230386 556608
rect 230442 556552 230447 556608
rect 178788 556550 230447 556552
rect 178788 556548 178794 556550
rect 230381 556547 230447 556550
rect 163497 556474 163563 556477
rect 175825 556474 175891 556477
rect 163497 556472 175891 556474
rect 163497 556416 163502 556472
rect 163558 556416 175830 556472
rect 175886 556416 175891 556472
rect 163497 556414 175891 556416
rect 163497 556411 163563 556414
rect 175825 556411 175891 556414
rect 228265 556474 228331 556477
rect 255221 556474 255287 556477
rect 228265 556472 255287 556474
rect 228265 556416 228270 556472
rect 228326 556416 255226 556472
rect 255282 556416 255287 556472
rect 228265 556414 255287 556416
rect 228265 556411 228331 556414
rect 255221 556411 255287 556414
rect 170305 556338 170371 556341
rect 179413 556338 179479 556341
rect 170305 556336 179479 556338
rect 170305 556280 170310 556336
rect 170366 556280 179418 556336
rect 179474 556280 179479 556336
rect 170305 556278 179479 556280
rect 170305 556275 170371 556278
rect 179413 556275 179479 556278
rect 47526 556140 47532 556204
rect 47596 556202 47602 556204
rect 53833 556202 53899 556205
rect 47596 556200 53899 556202
rect 47596 556144 53838 556200
rect 53894 556144 53899 556200
rect 47596 556142 53899 556144
rect 47596 556140 47602 556142
rect 53833 556139 53899 556142
rect 165521 556202 165587 556205
rect 175181 556202 175247 556205
rect 165521 556200 175247 556202
rect 165521 556144 165526 556200
rect 165582 556144 175186 556200
rect 175242 556144 175247 556200
rect 165521 556142 175247 556144
rect 165521 556139 165587 556142
rect 175181 556139 175247 556142
rect 288382 556140 288388 556204
rect 288452 556202 288458 556204
rect 289445 556202 289511 556205
rect 288452 556200 289511 556202
rect 288452 556144 289450 556200
rect 289506 556144 289511 556200
rect 288452 556142 289511 556144
rect 288452 556140 288458 556142
rect 289445 556139 289511 556142
rect 47853 556066 47919 556069
rect 165429 556066 165495 556069
rect 47853 556064 165495 556066
rect 47853 556008 47858 556064
rect 47914 556008 165434 556064
rect 165490 556008 165495 556064
rect 47853 556006 165495 556008
rect 47853 556003 47919 556006
rect 165429 556003 165495 556006
rect 176009 556066 176075 556069
rect 179413 556066 179479 556069
rect 176009 556064 179479 556066
rect 176009 556008 176014 556064
rect 176070 556008 179418 556064
rect 179474 556008 179479 556064
rect 176009 556006 179479 556008
rect 176009 556003 176075 556006
rect 179413 556003 179479 556006
rect 241421 556066 241487 556069
rect 254577 556066 254643 556069
rect 241421 556064 254643 556066
rect 241421 556008 241426 556064
rect 241482 556008 254582 556064
rect 254638 556008 254643 556064
rect 241421 556006 254643 556008
rect 241421 556003 241487 556006
rect 254577 556003 254643 556006
rect 137093 555930 137159 555933
rect 313917 555930 313983 555933
rect 137093 555928 313983 555930
rect 137093 555872 137098 555928
rect 137154 555872 313922 555928
rect 313978 555872 313983 555928
rect 137093 555870 313983 555872
rect 137093 555867 137159 555870
rect 313917 555867 313983 555870
rect 44817 555794 44883 555797
rect 162669 555794 162735 555797
rect 44817 555792 162735 555794
rect 44817 555736 44822 555792
rect 44878 555736 162674 555792
rect 162730 555736 162735 555792
rect 44817 555734 162735 555736
rect 44817 555731 44883 555734
rect 162669 555731 162735 555734
rect 176285 555794 176351 555797
rect 226333 555794 226399 555797
rect 176285 555792 226399 555794
rect 176285 555736 176290 555792
rect 176346 555736 226338 555792
rect 226394 555736 226399 555792
rect 176285 555734 226399 555736
rect 176285 555731 176351 555734
rect 226333 555731 226399 555734
rect 234337 555794 234403 555797
rect 289169 555794 289235 555797
rect 234337 555792 289235 555794
rect 234337 555736 234342 555792
rect 234398 555736 289174 555792
rect 289230 555736 289235 555792
rect 234337 555734 289235 555736
rect 234337 555731 234403 555734
rect 289169 555731 289235 555734
rect 293769 555794 293835 555797
rect 500033 555794 500099 555797
rect 293769 555792 500099 555794
rect 293769 555736 293774 555792
rect 293830 555736 500038 555792
rect 500094 555736 500099 555792
rect 293769 555734 500099 555736
rect 293769 555731 293835 555734
rect 500033 555731 500099 555734
rect 49417 555658 49483 555661
rect 165061 555658 165127 555661
rect 49417 555656 165127 555658
rect 49417 555600 49422 555656
rect 49478 555600 165066 555656
rect 165122 555600 165127 555656
rect 49417 555598 165127 555600
rect 49417 555595 49483 555598
rect 165061 555595 165127 555598
rect 178493 555658 178559 555661
rect 432689 555658 432755 555661
rect 178493 555656 432755 555658
rect 178493 555600 178498 555656
rect 178554 555600 432694 555656
rect 432750 555600 432755 555656
rect 178493 555598 432755 555600
rect 178493 555595 178559 555598
rect 432689 555595 432755 555598
rect 44909 555522 44975 555525
rect 159633 555522 159699 555525
rect 44909 555520 159699 555522
rect 44909 555464 44914 555520
rect 44970 555464 159638 555520
rect 159694 555464 159699 555520
rect 44909 555462 159699 555464
rect 44909 555459 44975 555462
rect 159633 555459 159699 555462
rect 172329 555522 172395 555525
rect 240041 555522 240107 555525
rect 172329 555520 240107 555522
rect 172329 555464 172334 555520
rect 172390 555464 240046 555520
rect 240102 555464 240107 555520
rect 172329 555462 240107 555464
rect 172329 555459 172395 555462
rect 240041 555459 240107 555462
rect 257613 555522 257679 555525
rect 515489 555522 515555 555525
rect 257613 555520 515555 555522
rect 257613 555464 257618 555520
rect 257674 555464 515494 555520
rect 515550 555464 515555 555520
rect 257613 555462 515555 555464
rect 257613 555459 257679 555462
rect 515489 555459 515555 555462
rect 55029 555386 55095 555389
rect 170029 555386 170095 555389
rect 55029 555384 170095 555386
rect 55029 555328 55034 555384
rect 55090 555328 170034 555384
rect 170090 555328 170095 555384
rect 55029 555326 170095 555328
rect 55029 555323 55095 555326
rect 170029 555323 170095 555326
rect 174445 555386 174511 555389
rect 433701 555386 433767 555389
rect 174445 555384 433767 555386
rect 174445 555328 174450 555384
rect 174506 555328 433706 555384
rect 433762 555328 433767 555384
rect 174445 555326 433767 555328
rect 174445 555323 174511 555326
rect 433701 555323 433767 555326
rect 46657 555250 46723 555253
rect 159449 555250 159515 555253
rect 46657 555248 159515 555250
rect 46657 555192 46662 555248
rect 46718 555192 159454 555248
rect 159510 555192 159515 555248
rect 46657 555190 159515 555192
rect 46657 555187 46723 555190
rect 159449 555187 159515 555190
rect 164877 555250 164943 555253
rect 178033 555250 178099 555253
rect 164877 555248 178099 555250
rect 164877 555192 164882 555248
rect 164938 555192 178038 555248
rect 178094 555192 178099 555248
rect 164877 555190 178099 555192
rect 164877 555187 164943 555190
rect 178033 555187 178099 555190
rect 179873 555250 179939 555253
rect 230197 555250 230263 555253
rect 179873 555248 230263 555250
rect 179873 555192 179878 555248
rect 179934 555192 230202 555248
rect 230258 555192 230263 555248
rect 179873 555190 230263 555192
rect 179873 555187 179939 555190
rect 230197 555187 230263 555190
rect 247125 555250 247191 555253
rect 247493 555250 247559 555253
rect 258901 555250 258967 555253
rect 247125 555248 258967 555250
rect 247125 555192 247130 555248
rect 247186 555192 247498 555248
rect 247554 555192 258906 555248
rect 258962 555192 258967 555248
rect 247125 555190 258967 555192
rect 247125 555187 247191 555190
rect 247493 555187 247559 555190
rect 258901 555187 258967 555190
rect 227253 555114 227319 555117
rect 255129 555114 255195 555117
rect 227253 555112 255195 555114
rect 227253 555056 227258 555112
rect 227314 555056 255134 555112
rect 255190 555056 255195 555112
rect 227253 555054 255195 555056
rect 227253 555051 227319 555054
rect 255129 555051 255195 555054
rect 35750 554916 35756 554980
rect 35820 554978 35826 554980
rect 53833 554978 53899 554981
rect 35820 554976 53899 554978
rect 35820 554920 53838 554976
rect 53894 554920 53899 554976
rect 35820 554918 53899 554920
rect 35820 554916 35826 554918
rect 53833 554915 53899 554918
rect 55806 554916 55812 554980
rect 55876 554978 55882 554980
rect 137185 554978 137251 554981
rect 55876 554976 137251 554978
rect 55876 554920 137190 554976
rect 137246 554920 137251 554976
rect 55876 554918 137251 554920
rect 55876 554916 55882 554918
rect 137185 554915 137251 554918
rect 173065 554978 173131 554981
rect 247033 554978 247099 554981
rect 173065 554976 247099 554978
rect 173065 554920 173070 554976
rect 173126 554920 247038 554976
rect 247094 554920 247099 554976
rect 173065 554918 247099 554920
rect 173065 554915 173131 554918
rect 247033 554915 247099 554918
rect 30966 554780 30972 554844
rect 31036 554842 31042 554844
rect 56501 554842 56567 554845
rect 31036 554840 56567 554842
rect 31036 554784 56506 554840
rect 56562 554784 56567 554840
rect 31036 554782 56567 554784
rect 31036 554780 31042 554782
rect 56501 554779 56567 554782
rect 162485 554842 162551 554845
rect 175825 554842 175891 554845
rect 162485 554840 175891 554842
rect 162485 554784 162490 554840
rect 162546 554784 175830 554840
rect 175886 554784 175891 554840
rect 162485 554782 175891 554784
rect 162485 554779 162551 554782
rect 175825 554779 175891 554782
rect 240133 554842 240199 554845
rect 241421 554842 241487 554845
rect 507853 554844 507919 554845
rect 523033 554844 523099 554845
rect 507853 554842 507900 554844
rect 240133 554840 241487 554842
rect 240133 554784 240138 554840
rect 240194 554784 241426 554840
rect 241482 554784 241487 554840
rect 240133 554782 241487 554784
rect 507808 554840 507900 554842
rect 507808 554784 507858 554840
rect 507808 554782 507900 554784
rect 240133 554779 240199 554782
rect 241421 554779 241487 554782
rect 507853 554780 507900 554782
rect 507964 554780 507970 554844
rect 522982 554780 522988 554844
rect 523052 554842 523099 554844
rect 523052 554840 523144 554842
rect 523094 554784 523144 554840
rect 523052 554782 523144 554784
rect 523052 554780 523099 554782
rect 507853 554779 507919 554780
rect 523033 554779 523099 554780
rect 177246 554644 177252 554708
rect 177316 554706 177322 554708
rect 177941 554706 178007 554709
rect 177316 554704 178007 554706
rect 177316 554648 177946 554704
rect 178002 554648 178007 554704
rect 177316 554646 178007 554648
rect 177316 554644 177322 554646
rect 177941 554643 178007 554646
rect 239397 554706 239463 554709
rect 240041 554706 240107 554709
rect 292113 554706 292179 554709
rect 239397 554704 292179 554706
rect 239397 554648 239402 554704
rect 239458 554648 240046 554704
rect 240102 554648 292118 554704
rect 292174 554648 292179 554704
rect 239397 554646 292179 554648
rect 239397 554643 239463 554646
rect 240041 554643 240107 554646
rect 292113 554643 292179 554646
rect 173709 554570 173775 554573
rect 240409 554570 240475 554573
rect 173709 554568 240475 554570
rect 173709 554512 173714 554568
rect 173770 554512 240414 554568
rect 240470 554512 240475 554568
rect 173709 554510 240475 554512
rect 173709 554507 173775 554510
rect 240409 554507 240475 554510
rect 257981 554570 258047 554573
rect 501597 554570 501663 554573
rect 257981 554568 501663 554570
rect 257981 554512 257986 554568
rect 258042 554512 501602 554568
rect 501658 554512 501663 554568
rect 257981 554510 501663 554512
rect 257981 554507 258047 554510
rect 501597 554507 501663 554510
rect 58566 554372 58572 554436
rect 58636 554434 58642 554436
rect 230381 554434 230447 554437
rect 58636 554432 230447 554434
rect 58636 554376 230386 554432
rect 230442 554376 230447 554432
rect 58636 554374 230447 554376
rect 58636 554372 58642 554374
rect 230381 554371 230447 554374
rect 257797 554434 257863 554437
rect 504449 554434 504515 554437
rect 257797 554432 504515 554434
rect 257797 554376 257802 554432
rect 257858 554376 504454 554432
rect 504510 554376 504515 554432
rect 257797 554374 504515 554376
rect 257797 554371 257863 554374
rect 504449 554371 504515 554374
rect 33910 554236 33916 554300
rect 33980 554298 33986 554300
rect 291929 554298 291995 554301
rect 33980 554296 291995 554298
rect 33980 554240 291934 554296
rect 291990 554240 291995 554296
rect 33980 554238 291995 554240
rect 33980 554236 33986 554238
rect 291929 554235 291995 554238
rect 54518 554100 54524 554164
rect 54588 554162 54594 554164
rect 178033 554162 178099 554165
rect 54588 554160 178099 554162
rect 54588 554104 178038 554160
rect 178094 554104 178099 554160
rect 54588 554102 178099 554104
rect 54588 554100 54594 554102
rect 178033 554099 178099 554102
rect 178534 554100 178540 554164
rect 178604 554162 178610 554164
rect 461025 554162 461091 554165
rect 178604 554160 461091 554162
rect 178604 554104 461030 554160
rect 461086 554104 461091 554160
rect 178604 554102 461091 554104
rect 178604 554100 178610 554102
rect 461025 554099 461091 554102
rect 59629 554026 59695 554029
rect 345657 554026 345723 554029
rect 59629 554024 345723 554026
rect -960 553890 480 553980
rect 59629 553968 59634 554024
rect 59690 553968 345662 554024
rect 345718 553968 345723 554024
rect 59629 553966 345723 553968
rect 59629 553963 59695 553966
rect 345657 553963 345723 553966
rect 18454 553890 18460 553892
rect -960 553830 18460 553890
rect -960 553740 480 553830
rect 18454 553828 18460 553830
rect 18524 553828 18530 553892
rect 35566 553828 35572 553892
rect 35636 553890 35642 553892
rect 173801 553890 173867 553893
rect 35636 553888 173867 553890
rect 35636 553832 173806 553888
rect 173862 553832 173867 553888
rect 35636 553830 173867 553832
rect 35636 553828 35642 553830
rect 173801 553827 173867 553830
rect 249517 553890 249583 553893
rect 258717 553890 258783 553893
rect 249517 553888 258783 553890
rect 249517 553832 249522 553888
rect 249578 553832 258722 553888
rect 258778 553832 258783 553888
rect 249517 553830 258783 553832
rect 249517 553827 249583 553830
rect 258717 553827 258783 553830
rect 34237 553754 34303 553757
rect 59997 553754 60063 553757
rect 34237 553752 60063 553754
rect 34237 553696 34242 553752
rect 34298 553696 60002 553752
rect 60058 553696 60063 553752
rect 34237 553694 60063 553696
rect 34237 553691 34303 553694
rect 59997 553691 60063 553694
rect 230197 553754 230263 553757
rect 254761 553754 254827 553757
rect 230197 553752 254827 553754
rect 230197 553696 230202 553752
rect 230258 553696 254766 553752
rect 254822 553696 254827 553752
rect 230197 553694 254827 553696
rect 230197 553691 230263 553694
rect 254761 553691 254827 553694
rect 40718 553556 40724 553620
rect 40788 553618 40794 553620
rect 240041 553618 240107 553621
rect 40788 553616 240107 553618
rect 40788 553560 240046 553616
rect 240102 553560 240107 553616
rect 40788 553558 240107 553560
rect 40788 553556 40794 553558
rect 240041 553555 240107 553558
rect 39798 553420 39804 553484
rect 39868 553482 39874 553484
rect 256693 553482 256759 553485
rect 39868 553480 256759 553482
rect 39868 553424 256698 553480
rect 256754 553424 256759 553480
rect 39868 553422 256759 553424
rect 39868 553420 39874 553422
rect 256693 553419 256759 553422
rect 58341 553346 58407 553349
rect 114461 553346 114527 553349
rect 58341 553344 114527 553346
rect 58341 553288 58346 553344
rect 58402 553288 114466 553344
rect 114522 553288 114527 553344
rect 58341 553286 114527 553288
rect 58341 553283 58407 553286
rect 114461 553283 114527 553286
rect 227345 553346 227411 553349
rect 234613 553346 234679 553349
rect 227345 553344 234679 553346
rect 227345 553288 227350 553344
rect 227406 553288 234618 553344
rect 234674 553288 234679 553344
rect 227345 553286 234679 553288
rect 227345 553283 227411 553286
rect 234613 553283 234679 553286
rect 248505 553346 248571 553349
rect 256509 553346 256575 553349
rect 248505 553344 256575 553346
rect 248505 553288 248510 553344
rect 248566 553288 256514 553344
rect 256570 553288 256575 553344
rect 248505 553286 256575 553288
rect 248505 553283 248571 553286
rect 256509 553283 256575 553286
rect 256693 553346 256759 553349
rect 260189 553346 260255 553349
rect 256693 553344 260255 553346
rect 256693 553288 256698 553344
rect 256754 553288 260194 553344
rect 260250 553288 260255 553344
rect 256693 553286 260255 553288
rect 256693 553283 256759 553286
rect 260189 553283 260255 553286
rect 97809 553210 97875 553213
rect 307201 553210 307267 553213
rect 97809 553208 307267 553210
rect 97809 553152 97814 553208
rect 97870 553152 307206 553208
rect 307262 553152 307267 553208
rect 97809 553150 307267 553152
rect 97809 553147 97875 553150
rect 307201 553147 307267 553150
rect 28441 553074 28507 553077
rect 97901 553074 97967 553077
rect 28441 553072 97967 553074
rect 28441 553016 28446 553072
rect 28502 553016 97906 553072
rect 97962 553016 97967 553072
rect 28441 553014 97967 553016
rect 28441 553011 28507 553014
rect 97901 553011 97967 553014
rect 98913 553074 98979 553077
rect 308213 553074 308279 553077
rect 98913 553072 308279 553074
rect 98913 553016 98918 553072
rect 98974 553016 308218 553072
rect 308274 553016 308279 553072
rect 98913 553014 308279 553016
rect 98913 553011 98979 553014
rect 308213 553011 308279 553014
rect 55765 552938 55831 552941
rect 253197 552938 253263 552941
rect 55765 552936 253263 552938
rect 55765 552880 55770 552936
rect 55826 552880 253202 552936
rect 253258 552880 253263 552936
rect 55765 552878 253263 552880
rect 55765 552875 55831 552878
rect 253197 552875 253263 552878
rect 253565 552938 253631 552941
rect 256693 552938 256759 552941
rect 253565 552936 256759 552938
rect 253565 552880 253570 552936
rect 253626 552880 256698 552936
rect 256754 552880 256759 552936
rect 253565 552878 256759 552880
rect 253565 552875 253631 552878
rect 256693 552875 256759 552878
rect 294873 552938 294939 552941
rect 509693 552938 509759 552941
rect 294873 552936 509759 552938
rect 294873 552880 294878 552936
rect 294934 552880 509698 552936
rect 509754 552880 509759 552936
rect 294873 552878 509759 552880
rect 294873 552875 294939 552878
rect 509693 552875 509759 552878
rect 56041 552802 56107 552805
rect 249701 552802 249767 552805
rect 56041 552800 249767 552802
rect 56041 552744 56046 552800
rect 56102 552744 249706 552800
rect 249762 552744 249767 552800
rect 56041 552742 249767 552744
rect 56041 552739 56107 552742
rect 249701 552739 249767 552742
rect 289537 552802 289603 552805
rect 504633 552802 504699 552805
rect 289537 552800 504699 552802
rect 289537 552744 289542 552800
rect 289598 552744 504638 552800
rect 504694 552744 504699 552800
rect 289537 552742 504699 552744
rect 289537 552739 289603 552742
rect 504633 552739 504699 552742
rect 39205 552666 39271 552669
rect 59169 552666 59235 552669
rect 39205 552664 59235 552666
rect 39205 552608 39210 552664
rect 39266 552608 59174 552664
rect 59230 552608 59235 552664
rect 39205 552606 59235 552608
rect 39205 552603 39271 552606
rect 59169 552603 59235 552606
rect 61561 552666 61627 552669
rect 336917 552666 336983 552669
rect 61561 552664 336983 552666
rect 61561 552608 61566 552664
rect 61622 552608 336922 552664
rect 336978 552608 336983 552664
rect 61561 552606 336983 552608
rect 61561 552603 61627 552606
rect 336917 552603 336983 552606
rect 43897 552530 43963 552533
rect 159541 552530 159607 552533
rect 43897 552528 159607 552530
rect 43897 552472 43902 552528
rect 43958 552472 159546 552528
rect 159602 552472 159607 552528
rect 43897 552470 159607 552472
rect 43897 552467 43963 552470
rect 159541 552467 159607 552470
rect 170029 552530 170095 552533
rect 227253 552530 227319 552533
rect 170029 552528 227319 552530
rect 170029 552472 170034 552528
rect 170090 552472 227258 552528
rect 227314 552472 227319 552528
rect 170029 552470 227319 552472
rect 170029 552467 170095 552470
rect 227253 552467 227319 552470
rect 235349 552530 235415 552533
rect 256233 552530 256299 552533
rect 235349 552528 256299 552530
rect 235349 552472 235354 552528
rect 235410 552472 256238 552528
rect 256294 552472 256299 552528
rect 235349 552470 256299 552472
rect 235349 552467 235415 552470
rect 256233 552467 256299 552470
rect 299749 552530 299815 552533
rect 502333 552530 502399 552533
rect 299749 552528 502399 552530
rect 299749 552472 299754 552528
rect 299810 552472 502338 552528
rect 502394 552472 502399 552528
rect 299749 552470 502399 552472
rect 299749 552467 299815 552470
rect 502333 552467 502399 552470
rect 38101 552394 38167 552397
rect 60825 552394 60891 552397
rect 38101 552392 60891 552394
rect 38101 552336 38106 552392
rect 38162 552336 60830 552392
rect 60886 552336 60891 552392
rect 38101 552334 60891 552336
rect 38101 552331 38167 552334
rect 60825 552331 60891 552334
rect 114093 552394 114159 552397
rect 323393 552394 323459 552397
rect 114093 552392 323459 552394
rect 114093 552336 114098 552392
rect 114154 552336 323398 552392
rect 323454 552336 323459 552392
rect 114093 552334 323459 552336
rect 114093 552331 114159 552334
rect 323393 552331 323459 552334
rect 30046 552196 30052 552260
rect 30116 552258 30122 552260
rect 98637 552258 98703 552261
rect 30116 552256 98703 552258
rect 30116 552200 98642 552256
rect 98698 552200 98703 552256
rect 30116 552198 98703 552200
rect 30116 552196 30122 552198
rect 98637 552195 98703 552198
rect 49417 552122 49483 552125
rect 56501 552122 56567 552125
rect 49417 552120 56567 552122
rect 49417 552064 49422 552120
rect 49478 552064 56506 552120
rect 56562 552064 56567 552120
rect 49417 552062 56567 552064
rect 49417 552059 49483 552062
rect 56501 552059 56567 552062
rect 112069 551986 112135 551989
rect 321369 551986 321435 551989
rect 112069 551984 321435 551986
rect 112069 551928 112074 551984
rect 112130 551928 321374 551984
rect 321430 551928 321435 551984
rect 112069 551926 321435 551928
rect 112069 551923 112135 551926
rect 321369 551923 321435 551926
rect 119153 551850 119219 551853
rect 328453 551850 328519 551853
rect 119153 551848 328519 551850
rect 119153 551792 119158 551848
rect 119214 551792 328458 551848
rect 328514 551792 328519 551848
rect 119153 551790 328519 551792
rect 119153 551787 119219 551790
rect 328453 551787 328519 551790
rect 67541 551714 67607 551717
rect 270769 551714 270835 551717
rect 67541 551712 270835 551714
rect 67541 551656 67546 551712
rect 67602 551656 270774 551712
rect 270830 551656 270835 551712
rect 67541 551654 270835 551656
rect 67541 551651 67607 551654
rect 270769 551651 270835 551654
rect 291142 551652 291148 551716
rect 291212 551714 291218 551716
rect 292297 551714 292363 551717
rect 539542 551714 539548 551716
rect 291212 551712 292363 551714
rect 291212 551656 292302 551712
rect 292358 551656 292363 551712
rect 291212 551654 292363 551656
rect 291212 551652 291218 551654
rect 292297 551651 292363 551654
rect 296670 551654 539548 551714
rect 59670 551516 59676 551580
rect 59740 551578 59746 551580
rect 235993 551578 236059 551581
rect 59740 551576 236059 551578
rect 59740 551520 235998 551576
rect 236054 551520 236059 551576
rect 59740 551518 236059 551520
rect 59740 551516 59746 551518
rect 235993 551515 236059 551518
rect 292062 551516 292068 551580
rect 292132 551578 292138 551580
rect 296670 551578 296730 551654
rect 539542 551652 539548 551654
rect 539612 551652 539618 551716
rect 292132 551518 296730 551578
rect 292132 551516 292138 551518
rect 59169 551442 59235 551445
rect 81433 551442 81499 551445
rect 59169 551440 81499 551442
rect 59169 551384 59174 551440
rect 59230 551384 81438 551440
rect 81494 551384 81499 551440
rect 59169 551382 81499 551384
rect 59169 551379 59235 551382
rect 81433 551379 81499 551382
rect 179454 551380 179460 551444
rect 179524 551442 179530 551444
rect 180057 551442 180123 551445
rect 179524 551440 180123 551442
rect 179524 551384 180062 551440
rect 180118 551384 180123 551440
rect 179524 551382 180123 551384
rect 179524 551380 179530 551382
rect 180057 551379 180123 551382
rect 185485 551442 185551 551445
rect 443821 551442 443887 551445
rect 185485 551440 443887 551442
rect 185485 551384 185490 551440
rect 185546 551384 443826 551440
rect 443882 551384 443887 551440
rect 185485 551382 443887 551384
rect 185485 551379 185551 551382
rect 443821 551379 443887 551382
rect 46565 551306 46631 551309
rect 111793 551306 111859 551309
rect 46565 551304 111859 551306
rect 46565 551248 46570 551304
rect 46626 551248 111798 551304
rect 111854 551248 111859 551304
rect 46565 551246 111859 551248
rect 46565 551243 46631 551246
rect 111793 551243 111859 551246
rect 172237 551306 172303 551309
rect 228265 551306 228331 551309
rect 172237 551304 228331 551306
rect 172237 551248 172242 551304
rect 172298 551248 228270 551304
rect 228326 551248 228331 551304
rect 172237 551246 228331 551248
rect 172237 551243 172303 551246
rect 228265 551243 228331 551246
rect 230381 551306 230447 551309
rect 509601 551306 509667 551309
rect 230381 551304 509667 551306
rect 230381 551248 230386 551304
rect 230442 551248 509606 551304
rect 509662 551248 509667 551304
rect 230381 551246 509667 551248
rect 230381 551243 230447 551246
rect 509601 551243 509667 551246
rect 81709 551170 81775 551173
rect 284937 551170 285003 551173
rect 81709 551168 285003 551170
rect 81709 551112 81714 551168
rect 81770 551112 284942 551168
rect 284998 551112 285003 551168
rect 81709 551110 285003 551112
rect 81709 551107 81775 551110
rect 284937 551107 285003 551110
rect 299105 551170 299171 551173
rect 503529 551170 503595 551173
rect 299105 551168 503595 551170
rect 299105 551112 299110 551168
rect 299166 551112 503534 551168
rect 503590 551112 503595 551168
rect 299105 551110 503595 551112
rect 299105 551107 299171 551110
rect 503529 551107 503595 551110
rect 36997 551034 37063 551037
rect 118693 551034 118759 551037
rect 36997 551032 118759 551034
rect 36997 550976 37002 551032
rect 37058 550976 118698 551032
rect 118754 550976 118759 551032
rect 36997 550974 118759 550976
rect 36997 550971 37063 550974
rect 118693 550971 118759 550974
rect 176469 551034 176535 551037
rect 185485 551034 185551 551037
rect 176469 551032 185551 551034
rect 176469 550976 176474 551032
rect 176530 550976 185490 551032
rect 185546 550976 185551 551032
rect 176469 550974 185551 550976
rect 176469 550971 176535 550974
rect 185485 550971 185551 550974
rect 236453 551034 236519 551037
rect 502057 551034 502123 551037
rect 236453 551032 502123 551034
rect 236453 550976 236458 551032
rect 236514 550976 502062 551032
rect 502118 550976 502123 551032
rect 583520 551020 584960 551260
rect 236453 550974 502123 550976
rect 236453 550971 236519 550974
rect 502057 550971 502123 550974
rect 59118 550836 59124 550900
rect 59188 550898 59194 550900
rect 175825 550898 175891 550901
rect 59188 550896 175891 550898
rect 59188 550840 175830 550896
rect 175886 550840 175891 550896
rect 59188 550838 175891 550840
rect 59188 550836 59194 550838
rect 175825 550835 175891 550838
rect 32438 550700 32444 550764
rect 32508 550762 32514 550764
rect 172421 550762 172487 550765
rect 509233 550764 509299 550765
rect 32508 550760 172487 550762
rect 32508 550704 172426 550760
rect 172482 550704 172487 550760
rect 32508 550702 172487 550704
rect 32508 550700 32514 550702
rect 172421 550699 172487 550702
rect 509182 550700 509188 550764
rect 509252 550762 509299 550764
rect 509252 550760 509344 550762
rect 509294 550704 509344 550760
rect 509252 550702 509344 550704
rect 509252 550700 509299 550702
rect 509233 550699 509299 550700
rect 57789 550626 57855 550629
rect 131113 550626 131179 550629
rect 57789 550624 131179 550626
rect 57789 550568 57794 550624
rect 57850 550568 131118 550624
rect 131174 550568 131179 550624
rect 57789 550566 131179 550568
rect 57789 550563 57855 550566
rect 131113 550563 131179 550566
rect 169477 550626 169543 550629
rect 234337 550626 234403 550629
rect 169477 550624 234403 550626
rect 169477 550568 169482 550624
rect 169538 550568 234342 550624
rect 234398 550568 234403 550624
rect 169477 550566 234403 550568
rect 169477 550563 169543 550566
rect 234337 550563 234403 550566
rect 296478 550564 296484 550628
rect 296548 550626 296554 550628
rect 502374 550626 502380 550628
rect 296548 550566 502380 550626
rect 296548 550564 296554 550566
rect 502374 550564 502380 550566
rect 502444 550564 502450 550628
rect 131297 550490 131363 550493
rect 340597 550490 340663 550493
rect 131297 550488 340663 550490
rect 131297 550432 131302 550488
rect 131358 550432 340602 550488
rect 340658 550432 340663 550488
rect 131297 550430 340663 550432
rect 131297 550427 131363 550430
rect 340597 550427 340663 550430
rect 99925 550354 99991 550357
rect 309225 550354 309291 550357
rect 99925 550352 309291 550354
rect 99925 550296 99930 550352
rect 99986 550296 309230 550352
rect 309286 550296 309291 550352
rect 99925 550294 309291 550296
rect 99925 550291 99991 550294
rect 309225 550291 309291 550294
rect 80697 550218 80763 550221
rect 283925 550218 283991 550221
rect 80697 550216 283991 550218
rect 80697 550160 80702 550216
rect 80758 550160 283930 550216
rect 283986 550160 283991 550216
rect 80697 550158 283991 550160
rect 80697 550155 80763 550158
rect 283925 550155 283991 550158
rect 288341 550218 288407 550221
rect 296529 550220 296595 550221
rect 296478 550218 296484 550220
rect 288341 550216 296362 550218
rect 288341 550160 288346 550216
rect 288402 550160 296362 550216
rect 288341 550158 296362 550160
rect 296438 550158 296484 550218
rect 296548 550216 296595 550220
rect 499021 550218 499087 550221
rect 296590 550160 296595 550216
rect 288341 550155 288407 550158
rect 50521 550082 50587 550085
rect 80053 550082 80119 550085
rect 50521 550080 80119 550082
rect 50521 550024 50526 550080
rect 50582 550024 80058 550080
rect 80114 550024 80119 550080
rect 50521 550022 80119 550024
rect 50521 550019 50587 550022
rect 80053 550019 80119 550022
rect 92841 550082 92907 550085
rect 296069 550082 296135 550085
rect 92841 550080 296135 550082
rect 92841 550024 92846 550080
rect 92902 550024 296074 550080
rect 296130 550024 296135 550080
rect 92841 550022 296135 550024
rect 296302 550082 296362 550158
rect 296478 550156 296484 550158
rect 296548 550156 296595 550160
rect 296529 550155 296595 550156
rect 296670 550216 499087 550218
rect 296670 550160 499026 550216
rect 499082 550160 499087 550216
rect 296670 550158 499087 550160
rect 296670 550082 296730 550158
rect 499021 550155 499087 550158
rect 296302 550022 296730 550082
rect 92841 550019 92907 550022
rect 296069 550019 296135 550022
rect 298870 550020 298876 550084
rect 298940 550082 298946 550084
rect 511022 550082 511028 550084
rect 298940 550022 511028 550082
rect 298940 550020 298946 550022
rect 511022 550020 511028 550022
rect 511092 550020 511098 550084
rect 57237 549946 57303 549949
rect 228357 549946 228423 549949
rect 57237 549944 228423 549946
rect 57237 549888 57242 549944
rect 57298 549888 228362 549944
rect 228418 549888 228423 549944
rect 57237 549886 228423 549888
rect 57237 549883 57303 549886
rect 228357 549883 228423 549886
rect 243261 549946 243327 549949
rect 499757 549946 499823 549949
rect 243261 549944 499823 549946
rect 243261 549888 243266 549944
rect 243322 549888 499762 549944
rect 499818 549888 499823 549944
rect 243261 549886 499823 549888
rect 243261 549883 243327 549886
rect 499757 549883 499823 549886
rect 44633 549810 44699 549813
rect 92473 549810 92539 549813
rect 176561 549812 176627 549813
rect 176510 549810 176516 549812
rect 44633 549808 92539 549810
rect 44633 549752 44638 549808
rect 44694 549752 92478 549808
rect 92534 549752 92539 549808
rect 44633 549750 92539 549752
rect 176470 549750 176516 549810
rect 176580 549808 176627 549812
rect 229277 549810 229343 549813
rect 230197 549810 230263 549813
rect 176622 549752 176627 549808
rect 44633 549747 44699 549750
rect 92473 549747 92539 549750
rect 176510 549748 176516 549750
rect 176580 549748 176627 549752
rect 176561 549747 176627 549748
rect 180750 549808 230263 549810
rect 180750 549752 229282 549808
rect 229338 549752 230202 549808
rect 230258 549752 230263 549808
rect 180750 549750 230263 549752
rect 27245 549674 27311 549677
rect 99373 549674 99439 549677
rect 27245 549672 99439 549674
rect 27245 549616 27250 549672
rect 27306 549616 99378 549672
rect 99434 549616 99439 549672
rect 27245 549614 99439 549616
rect 27245 549611 27311 549614
rect 99373 549611 99439 549614
rect 173709 549674 173775 549677
rect 180750 549674 180810 549750
rect 229277 549747 229343 549750
rect 230197 549747 230263 549750
rect 232313 549810 232379 549813
rect 256141 549810 256207 549813
rect 232313 549808 256207 549810
rect 232313 549752 232318 549808
rect 232374 549752 256146 549808
rect 256202 549752 256207 549808
rect 232313 549750 256207 549752
rect 232313 549747 232379 549750
rect 256141 549747 256207 549750
rect 173709 549672 180810 549674
rect 173709 549616 173714 549672
rect 173770 549616 180810 549672
rect 173709 549614 180810 549616
rect 173709 549611 173775 549614
rect 35617 549538 35683 549541
rect 168373 549538 168439 549541
rect 35617 549536 168439 549538
rect 35617 549480 35622 549536
rect 35678 549480 168378 549536
rect 168434 549480 168439 549536
rect 35617 549478 168439 549480
rect 35617 549475 35683 549478
rect 168373 549475 168439 549478
rect 36854 549340 36860 549404
rect 36924 549402 36930 549404
rect 173801 549402 173867 549405
rect 36924 549400 173867 549402
rect 36924 549344 173806 549400
rect 173862 549344 173867 549400
rect 36924 549342 173867 549344
rect 36924 549340 36930 549342
rect 173801 549339 173867 549342
rect 111057 549266 111123 549269
rect 320357 549266 320423 549269
rect 111057 549264 320423 549266
rect 111057 549208 111062 549264
rect 111118 549208 320362 549264
rect 320418 549208 320423 549264
rect 111057 549206 320423 549208
rect 111057 549203 111123 549206
rect 320357 549203 320423 549206
rect 78673 549130 78739 549133
rect 281901 549130 281967 549133
rect 78673 549128 281967 549130
rect 78673 549072 78678 549128
rect 78734 549072 281906 549128
rect 281962 549072 281967 549128
rect 78673 549070 281967 549072
rect 78673 549067 78739 549070
rect 281901 549067 281967 549070
rect 288566 549068 288572 549132
rect 288636 549130 288642 549132
rect 289721 549130 289787 549133
rect 288636 549128 289787 549130
rect 288636 549072 289726 549128
rect 289782 549072 289787 549128
rect 288636 549070 289787 549072
rect 288636 549068 288642 549070
rect 289721 549067 289787 549070
rect 290958 549068 290964 549132
rect 291028 549130 291034 549132
rect 514150 549130 514156 549132
rect 291028 549070 514156 549130
rect 291028 549068 291034 549070
rect 514150 549068 514156 549070
rect 514220 549068 514226 549132
rect 63493 548994 63559 548997
rect 266721 548994 266787 548997
rect 63493 548992 266787 548994
rect 63493 548936 63498 548992
rect 63554 548936 266726 548992
rect 266782 548936 266787 548992
rect 63493 548934 266787 548936
rect 63493 548931 63559 548934
rect 266721 548931 266787 548934
rect 289486 548932 289492 548996
rect 289556 548994 289562 548996
rect 529054 548994 529060 548996
rect 289556 548934 529060 548994
rect 289556 548932 289562 548934
rect 529054 548932 529060 548934
rect 529124 548932 529130 548996
rect 178677 548858 178743 548861
rect 426617 548858 426683 548861
rect 178677 548856 426683 548858
rect 178677 548800 178682 548856
rect 178738 548800 426622 548856
rect 426678 548800 426683 548856
rect 178677 548798 426683 548800
rect 178677 548795 178743 548798
rect 426617 548795 426683 548798
rect 228081 548722 228147 548725
rect 510889 548722 510955 548725
rect 228081 548720 510955 548722
rect 228081 548664 228086 548720
rect 228142 548664 510894 548720
rect 510950 548664 510955 548720
rect 228081 548662 510955 548664
rect 228081 548659 228147 548662
rect 510889 548659 510955 548662
rect 59721 548586 59787 548589
rect 358813 548586 358879 548589
rect 59721 548584 358879 548586
rect 59721 548528 59726 548584
rect 59782 548528 358818 548584
rect 358874 548528 358879 548584
rect 59721 548526 358879 548528
rect 59721 548523 59787 548526
rect 358813 548523 358879 548526
rect 30230 548388 30236 548452
rect 30300 548450 30306 548452
rect 79317 548450 79383 548453
rect 30300 548448 79383 548450
rect 30300 548392 79322 548448
rect 79378 548392 79383 548448
rect 30300 548390 79383 548392
rect 30300 548388 30306 548390
rect 79317 548387 79383 548390
rect 174813 548450 174879 548453
rect 227713 548450 227779 548453
rect 174813 548448 227779 548450
rect 174813 548392 174818 548448
rect 174874 548392 227718 548448
rect 227774 548392 227779 548448
rect 174813 548390 227779 548392
rect 174813 548387 174879 548390
rect 227713 548387 227779 548390
rect 59077 548314 59143 548317
rect 110413 548314 110479 548317
rect 59077 548312 110479 548314
rect 59077 548256 59082 548312
rect 59138 548256 110418 548312
rect 110474 548256 110479 548312
rect 59077 548254 110479 548256
rect 59077 548251 59143 548254
rect 110413 548251 110479 548254
rect 169937 548314 170003 548317
rect 232313 548314 232379 548317
rect 169937 548312 232379 548314
rect 169937 548256 169942 548312
rect 169998 548256 232318 548312
rect 232374 548256 232379 548312
rect 169937 548254 232379 548256
rect 169937 548251 170003 548254
rect 232313 548251 232379 548254
rect 47761 548178 47827 548181
rect 169753 548178 169819 548181
rect 47761 548176 169819 548178
rect 47761 548120 47766 548176
rect 47822 548120 169758 548176
rect 169814 548120 169819 548176
rect 47761 548118 169819 548120
rect 47761 548115 47827 548118
rect 169753 548115 169819 548118
rect 43161 548042 43227 548045
rect 178033 548042 178099 548045
rect 43161 548040 178099 548042
rect 43161 547984 43166 548040
rect 43222 547984 178038 548040
rect 178094 547984 178099 548040
rect 43161 547982 178099 547984
rect 43161 547979 43227 547982
rect 178033 547979 178099 547982
rect 38377 547906 38443 547909
rect 175181 547906 175247 547909
rect 38377 547904 175247 547906
rect 38377 547848 38382 547904
rect 38438 547848 175186 547904
rect 175242 547848 175247 547904
rect 38377 547846 175247 547848
rect 38377 547843 38443 547846
rect 175181 547843 175247 547846
rect 506473 547906 506539 547909
rect 506606 547906 506612 547908
rect 506473 547904 506612 547906
rect 506473 547848 506478 547904
rect 506534 547848 506612 547904
rect 506473 547846 506612 547848
rect 506473 547843 506539 547846
rect 506606 547844 506612 547846
rect 506676 547844 506682 547908
rect 88793 547770 88859 547773
rect 292021 547770 292087 547773
rect 88793 547768 292087 547770
rect 88793 547712 88798 547768
rect 88854 547712 292026 547768
rect 292082 547712 292087 547768
rect 88793 547710 292087 547712
rect 88793 547707 88859 547710
rect 292021 547707 292087 547710
rect 295057 547770 295123 547773
rect 502517 547770 502583 547773
rect 295057 547768 502583 547770
rect 295057 547712 295062 547768
rect 295118 547712 502522 547768
rect 502578 547712 502583 547768
rect 295057 547710 502583 547712
rect 295057 547707 295123 547710
rect 502517 547707 502583 547710
rect 66529 547634 66595 547637
rect 264237 547634 264303 547637
rect 66529 547632 264303 547634
rect 66529 547576 66534 547632
rect 66590 547576 264242 547632
rect 264298 547576 264303 547632
rect 66529 547574 264303 547576
rect 66529 547571 66595 547574
rect 264237 547571 264303 547574
rect 283966 547572 283972 547636
rect 284036 547634 284042 547636
rect 498694 547634 498700 547636
rect 284036 547574 498700 547634
rect 284036 547572 284042 547574
rect 498694 547572 498700 547574
rect 498764 547572 498770 547636
rect 37038 547436 37044 547500
rect 37108 547498 37114 547500
rect 292246 547498 292252 547500
rect 37108 547438 292252 547498
rect 37108 547436 37114 547438
rect 292246 547436 292252 547438
rect 292316 547436 292322 547500
rect 293166 547436 293172 547500
rect 293236 547498 293242 547500
rect 519302 547498 519308 547500
rect 293236 547438 519308 547498
rect 293236 547436 293242 547438
rect 519302 547436 519308 547438
rect 519372 547436 519378 547500
rect 58249 547362 58315 547365
rect 231761 547362 231827 547365
rect 58249 547360 231827 547362
rect 58249 547304 58254 547360
rect 58310 547304 231766 547360
rect 231822 547304 231827 547360
rect 58249 547302 231827 547304
rect 58249 547299 58315 547302
rect 231761 547299 231827 547302
rect 235165 547362 235231 547365
rect 499665 547362 499731 547365
rect 235165 547360 499731 547362
rect 235165 547304 235170 547360
rect 235226 547304 499670 547360
rect 499726 547304 499731 547360
rect 235165 547302 499731 547304
rect 235165 547299 235231 547302
rect 499665 547299 499731 547302
rect 175038 547164 175044 547228
rect 175108 547226 175114 547228
rect 175181 547226 175247 547229
rect 175108 547224 175247 547226
rect 175108 547168 175186 547224
rect 175242 547168 175247 547224
rect 175108 547166 175247 547168
rect 175108 547164 175114 547166
rect 175181 547163 175247 547166
rect 231117 547226 231183 547229
rect 510981 547226 511047 547229
rect 231117 547224 511047 547226
rect 231117 547168 231122 547224
rect 231178 547168 510986 547224
rect 511042 547168 511047 547224
rect 231117 547166 511047 547168
rect 231117 547163 231183 547166
rect 510981 547163 511047 547166
rect 57421 547090 57487 547093
rect 359825 547090 359891 547093
rect 57421 547088 359891 547090
rect 57421 547032 57426 547088
rect 57482 547032 359830 547088
rect 359886 547032 359891 547088
rect 57421 547030 359891 547032
rect 57421 547027 57487 547030
rect 359825 547027 359891 547030
rect 50429 546954 50495 546957
rect 67541 546954 67607 546957
rect 50429 546952 67607 546954
rect 50429 546896 50434 546952
rect 50490 546896 67546 546952
rect 67602 546896 67607 546952
rect 50429 546894 67607 546896
rect 50429 546891 50495 546894
rect 67541 546891 67607 546894
rect 136173 546954 136239 546957
rect 258625 546954 258691 546957
rect 136173 546952 258691 546954
rect 136173 546896 136178 546952
rect 136234 546896 258630 546952
rect 258686 546896 258691 546952
rect 136173 546894 258691 546896
rect 136173 546891 136239 546894
rect 258625 546891 258691 546894
rect 33869 546818 33935 546821
rect 88977 546818 89043 546821
rect 33869 546816 89043 546818
rect 33869 546760 33874 546816
rect 33930 546760 88982 546816
rect 89038 546760 89043 546816
rect 33869 546758 89043 546760
rect 33869 546755 33935 546758
rect 88977 546755 89043 546758
rect 166809 546818 166875 546821
rect 235349 546818 235415 546821
rect 166809 546816 235415 546818
rect 166809 546760 166814 546816
rect 166870 546760 235354 546816
rect 235410 546760 235415 546816
rect 166809 546758 235415 546760
rect 166809 546755 166875 546758
rect 235349 546755 235415 546758
rect 56041 546682 56107 546685
rect 136541 546682 136607 546685
rect 56041 546680 136607 546682
rect 56041 546624 56046 546680
rect 56102 546624 136546 546680
rect 136602 546624 136607 546680
rect 56041 546622 136607 546624
rect 56041 546619 56107 546622
rect 136541 546619 136607 546622
rect 29862 546484 29868 546548
rect 29932 546546 29938 546548
rect 166165 546546 166231 546549
rect 29932 546544 166231 546546
rect 29932 546488 166170 546544
rect 166226 546488 166231 546544
rect 29932 546486 166231 546488
rect 29932 546484 29938 546486
rect 166165 546483 166231 546486
rect 282862 546484 282868 546548
rect 282932 546546 282938 546548
rect 284201 546546 284267 546549
rect 282932 546544 284267 546546
rect 282932 546488 284206 546544
rect 284262 546488 284267 546544
rect 282932 546486 284267 546488
rect 282932 546484 282938 546486
rect 284201 546483 284267 546486
rect 292614 546484 292620 546548
rect 292684 546546 292690 546548
rect 293861 546546 293927 546549
rect 503713 546548 503779 546549
rect 292684 546544 293927 546546
rect 292684 546488 293866 546544
rect 293922 546488 293927 546544
rect 292684 546486 293927 546488
rect 292684 546484 292690 546486
rect 293861 546483 293927 546486
rect 503662 546484 503668 546548
rect 503732 546546 503779 546548
rect 503732 546544 503824 546546
rect 503774 546488 503824 546544
rect 503732 546486 503824 546488
rect 503732 546484 503779 546486
rect 503713 546483 503779 546484
rect 253933 546410 253999 546413
rect 255078 546410 255084 546412
rect 253933 546408 255084 546410
rect 253933 546352 253938 546408
rect 253994 546352 255084 546408
rect 253933 546350 255084 546352
rect 253933 546347 253999 546350
rect 255078 546348 255084 546350
rect 255148 546348 255154 546412
rect 74625 546274 74691 546277
rect 277853 546274 277919 546277
rect 74625 546272 277919 546274
rect 74625 546216 74630 546272
rect 74686 546216 277858 546272
rect 277914 546216 277919 546272
rect 74625 546214 277919 546216
rect 74625 546211 74691 546214
rect 277853 546211 277919 546214
rect 284886 546212 284892 546276
rect 284956 546274 284962 546276
rect 508262 546274 508268 546276
rect 284956 546214 508268 546274
rect 284956 546212 284962 546214
rect 508262 546212 508268 546214
rect 508332 546212 508338 546276
rect 34094 546076 34100 546140
rect 34164 546138 34170 546140
rect 286542 546138 286548 546140
rect 34164 546078 286548 546138
rect 34164 546076 34170 546078
rect 286542 546076 286548 546078
rect 286612 546076 286618 546140
rect 288198 546076 288204 546140
rect 288268 546138 288274 546140
rect 497406 546138 497412 546140
rect 288268 546078 497412 546138
rect 288268 546076 288274 546078
rect 497406 546076 497412 546078
rect 497476 546076 497482 546140
rect 35525 546002 35591 546005
rect 224125 546002 224191 546005
rect 35525 546000 224191 546002
rect 35525 545944 35530 546000
rect 35586 545944 224130 546000
rect 224186 545944 224191 546000
rect 35525 545942 224191 545944
rect 35525 545939 35591 545942
rect 224125 545939 224191 545942
rect 56133 545866 56199 545869
rect 362861 545866 362927 545869
rect 56133 545864 362927 545866
rect 56133 545808 56138 545864
rect 56194 545808 362866 545864
rect 362922 545808 362927 545864
rect 56133 545806 362927 545808
rect 56133 545803 56199 545806
rect 362861 545803 362927 545806
rect 27470 545668 27476 545732
rect 27540 545730 27546 545732
rect 382222 545730 382228 545732
rect 27540 545670 382228 545730
rect 27540 545668 27546 545670
rect 382222 545668 382228 545670
rect 382292 545668 382298 545732
rect 47669 545594 47735 545597
rect 75821 545594 75887 545597
rect 47669 545592 75887 545594
rect 47669 545536 47674 545592
rect 47730 545536 75826 545592
rect 75882 545536 75887 545592
rect 47669 545534 75887 545536
rect 47669 545531 47735 545534
rect 75821 545531 75887 545534
rect 86769 545594 86835 545597
rect 289997 545594 290063 545597
rect 86769 545592 290063 545594
rect 86769 545536 86774 545592
rect 86830 545536 290002 545592
rect 290058 545536 290063 545592
rect 86769 545534 290063 545536
rect 86769 545531 86835 545534
rect 289997 545531 290063 545534
rect 46381 545458 46447 545461
rect 86861 545458 86927 545461
rect 46381 545456 86927 545458
rect 46381 545400 46386 545456
rect 46442 545400 86866 545456
rect 86922 545400 86927 545456
rect 46381 545398 86927 545400
rect 46381 545395 46447 545398
rect 86861 545395 86927 545398
rect 126237 545458 126303 545461
rect 335537 545458 335603 545461
rect 126237 545456 335603 545458
rect 126237 545400 126242 545456
rect 126298 545400 335542 545456
rect 335598 545400 335603 545456
rect 126237 545398 335603 545400
rect 126237 545395 126303 545398
rect 335537 545395 335603 545398
rect 36905 545322 36971 545325
rect 126881 545322 126947 545325
rect 36905 545320 126947 545322
rect 36905 545264 36910 545320
rect 36966 545264 126886 545320
rect 126942 545264 126947 545320
rect 36905 545262 126947 545264
rect 36905 545259 36971 545262
rect 126881 545259 126947 545262
rect 224033 545322 224099 545325
rect 512085 545322 512151 545325
rect 224033 545320 512151 545322
rect 224033 545264 224038 545320
rect 224094 545264 512090 545320
rect 512146 545264 512151 545320
rect 224033 545262 512151 545264
rect 224033 545259 224099 545262
rect 512085 545259 512151 545262
rect 50337 545186 50403 545189
rect 56501 545186 56567 545189
rect 50337 545184 56567 545186
rect 50337 545128 50342 545184
rect 50398 545128 56506 545184
rect 56562 545128 56567 545184
rect 50337 545126 56567 545128
rect 50337 545123 50403 545126
rect 56501 545123 56567 545126
rect 75637 545050 75703 545053
rect 278865 545050 278931 545053
rect 75637 545048 278931 545050
rect 75637 544992 75642 545048
rect 75698 544992 278870 545048
rect 278926 544992 278931 545048
rect 75637 544990 278931 544992
rect 75637 544987 75703 544990
rect 278865 544987 278931 544990
rect 296294 544988 296300 545052
rect 296364 545050 296370 545052
rect 502558 545050 502564 545052
rect 296364 544990 502564 545050
rect 296364 544988 296370 544990
rect 502558 544988 502564 544990
rect 502628 544988 502634 545052
rect 132309 544914 132375 544917
rect 341609 544914 341675 544917
rect 132309 544912 341675 544914
rect 132309 544856 132314 544912
rect 132370 544856 341614 544912
rect 341670 544856 341675 544912
rect 132309 544854 341675 544856
rect 132309 544851 132375 544854
rect 341609 544851 341675 544854
rect 251357 544778 251423 544781
rect 512269 544778 512335 544781
rect 251357 544776 512335 544778
rect 251357 544720 251362 544776
rect 251418 544720 512274 544776
rect 512330 544720 512335 544776
rect 251357 544718 512335 544720
rect 251357 544715 251423 544718
rect 512269 544715 512335 544718
rect 49325 544642 49391 544645
rect 75821 544642 75887 544645
rect 49325 544640 75887 544642
rect 49325 544584 49330 544640
rect 49386 544584 75826 544640
rect 75882 544584 75887 544640
rect 49325 544582 75887 544584
rect 49325 544579 49391 544582
rect 75821 544579 75887 544582
rect 170673 544642 170739 544645
rect 455965 544642 456031 544645
rect 170673 544640 456031 544642
rect 170673 544584 170678 544640
rect 170734 544584 455970 544640
rect 456026 544584 456031 544640
rect 170673 544582 456031 544584
rect 170673 544579 170739 544582
rect 455965 544579 456031 544582
rect 57697 544506 57763 544509
rect 350717 544506 350783 544509
rect 57697 544504 350783 544506
rect 57697 544448 57702 544504
rect 57758 544448 350722 544504
rect 350778 544448 350783 544504
rect 57697 544446 350783 544448
rect 57697 544443 57763 544446
rect 350717 544443 350783 544446
rect 58985 544370 59051 544373
rect 366909 544370 366975 544373
rect 58985 544368 366975 544370
rect 58985 544312 58990 544368
rect 59046 544312 366914 544368
rect 366970 544312 366975 544368
rect 58985 544310 366975 544312
rect 58985 544307 59051 544310
rect 366909 544307 366975 544310
rect 54661 544234 54727 544237
rect 88241 544234 88307 544237
rect 54661 544232 88307 544234
rect 54661 544176 54666 544232
rect 54722 544176 88246 544232
rect 88302 544176 88307 544232
rect 54661 544174 88307 544176
rect 54661 544171 54727 544174
rect 88241 544171 88307 544174
rect 88425 544234 88491 544237
rect 290825 544234 290891 544237
rect 88425 544232 290891 544234
rect 88425 544176 88430 544232
rect 88486 544176 290830 544232
rect 290886 544176 290891 544232
rect 88425 544174 290891 544176
rect 88425 544171 88491 544174
rect 290825 544171 290891 544174
rect 28349 544098 28415 544101
rect 131113 544098 131179 544101
rect 28349 544096 131179 544098
rect 28349 544040 28354 544096
rect 28410 544040 131118 544096
rect 131174 544040 131179 544096
rect 28349 544038 131179 544040
rect 28349 544035 28415 544038
rect 131113 544035 131179 544038
rect 217961 544098 218027 544101
rect 252461 544098 252527 544101
rect 217961 544096 252527 544098
rect 217961 544040 217966 544096
rect 218022 544040 252466 544096
rect 252522 544040 252527 544096
rect 217961 544038 252527 544040
rect 217961 544035 218027 544038
rect 252461 544035 252527 544038
rect 36813 543962 36879 543965
rect 169753 543962 169819 543965
rect 36813 543960 169819 543962
rect 36813 543904 36818 543960
rect 36874 543904 169758 543960
rect 169814 543904 169819 543960
rect 36813 543902 169819 543904
rect 36813 543899 36879 543902
rect 169753 543899 169819 543902
rect 28758 543764 28764 543828
rect 28828 543826 28834 543828
rect 216673 543826 216739 543829
rect 28828 543824 216739 543826
rect 28828 543768 216678 543824
rect 216734 543768 216739 543824
rect 28828 543766 216739 543768
rect 28828 543764 28834 543766
rect 216673 543763 216739 543766
rect 299197 543826 299263 543829
rect 299197 543824 299490 543826
rect 299197 543768 299202 543824
rect 299258 543768 299490 543824
rect 299197 543766 299490 543768
rect 299197 543763 299263 543766
rect 82721 543690 82787 543693
rect 285949 543690 286015 543693
rect 82721 543688 286015 543690
rect 82721 543632 82726 543688
rect 82782 543632 285954 543688
rect 286010 543632 286015 543688
rect 82721 543630 286015 543632
rect 82721 543627 82787 543630
rect 285949 543627 286015 543630
rect 292481 543690 292547 543693
rect 299197 543690 299263 543693
rect 292481 543688 299263 543690
rect 292481 543632 292486 543688
rect 292542 543632 299202 543688
rect 299258 543632 299263 543688
rect 292481 543630 299263 543632
rect 299430 543690 299490 543766
rect 502609 543690 502675 543693
rect 299430 543688 502675 543690
rect 299430 543632 502614 543688
rect 502670 543632 502675 543688
rect 299430 543630 502675 543632
rect 292481 543627 292547 543630
rect 299197 543627 299263 543630
rect 502609 543627 502675 543630
rect 127249 543554 127315 543557
rect 336549 543554 336615 543557
rect 127249 543552 336615 543554
rect 127249 543496 127254 543552
rect 127310 543496 336554 543552
rect 336610 543496 336615 543552
rect 127249 543494 336615 543496
rect 127249 543491 127315 543494
rect 336549 543491 336615 543494
rect 71589 543418 71655 543421
rect 274817 543418 274883 543421
rect 71589 543416 274883 543418
rect 71589 543360 71594 543416
rect 71650 543360 274822 543416
rect 274878 543360 274883 543416
rect 71589 543358 274883 543360
rect 71589 543355 71655 543358
rect 274817 543355 274883 543358
rect 292982 543356 292988 543420
rect 293052 543418 293058 543420
rect 516174 543418 516180 543420
rect 293052 543358 516180 543418
rect 293052 543356 293058 543358
rect 516174 543356 516180 543358
rect 516244 543356 516250 543420
rect 239213 543282 239279 543285
rect 499849 543282 499915 543285
rect 239213 543280 499915 543282
rect 239213 543224 239218 543280
rect 239274 543224 499854 543280
rect 499910 543224 499915 543280
rect 239213 543222 499915 543224
rect 239213 543219 239279 543222
rect 499849 543219 499915 543222
rect 242249 543146 242315 543149
rect 519445 543146 519511 543149
rect 242249 543144 519511 543146
rect 242249 543088 242254 543144
rect 242310 543088 519450 543144
rect 519506 543088 519511 543144
rect 242249 543086 519511 543088
rect 242249 543083 242315 543086
rect 519445 543083 519511 543086
rect 57145 543010 57211 543013
rect 349705 543010 349771 543013
rect 57145 543008 349771 543010
rect 57145 542952 57150 543008
rect 57206 542952 349710 543008
rect 349766 542952 349771 543008
rect 57145 542950 349771 542952
rect 57145 542947 57211 542950
rect 349705 542947 349771 542950
rect 25497 542874 25563 542877
rect 127617 542874 127683 542877
rect 25497 542872 127683 542874
rect 25497 542816 25502 542872
rect 25558 542816 127622 542872
rect 127678 542816 127683 542872
rect 25497 542814 127683 542816
rect 25497 542811 25563 542814
rect 127617 542811 127683 542814
rect 208853 542874 208919 542877
rect 242801 542874 242867 542877
rect 208853 542872 242867 542874
rect 208853 542816 208858 542872
rect 208914 542816 242806 542872
rect 242862 542816 242867 542872
rect 208853 542814 242867 542816
rect 208853 542811 208919 542814
rect 242801 542811 242867 542814
rect 244365 542874 244431 542877
rect 350533 542874 350599 542877
rect 244365 542872 350599 542874
rect 244365 542816 244370 542872
rect 244426 542816 350538 542872
rect 350594 542816 350599 542872
rect 244365 542814 350599 542816
rect 244365 542811 244431 542814
rect 350533 542811 350599 542814
rect 55673 542738 55739 542741
rect 208393 542738 208459 542741
rect 55673 542736 208459 542738
rect 55673 542680 55678 542736
rect 55734 542680 208398 542736
rect 208454 542680 208459 542736
rect 55673 542678 208459 542680
rect 55673 542675 55739 542678
rect 208393 542675 208459 542678
rect 55949 542602 56015 542605
rect 240041 542602 240107 542605
rect 55949 542600 240107 542602
rect 55949 542544 55954 542600
rect 56010 542544 240046 542600
rect 240102 542544 240107 542600
rect 55949 542542 240107 542544
rect 55949 542539 56015 542542
rect 240041 542539 240107 542542
rect 34145 542466 34211 542469
rect 244273 542466 244339 542469
rect 34145 542464 244339 542466
rect 34145 542408 34150 542464
rect 34206 542408 244278 542464
rect 244334 542408 244339 542464
rect 34145 542406 244339 542408
rect 34145 542403 34211 542406
rect 244273 542403 244339 542406
rect 296662 542404 296668 542468
rect 296732 542466 296738 542468
rect 298001 542466 298067 542469
rect 296732 542464 298067 542466
rect 296732 542408 298006 542464
rect 298062 542408 298067 542464
rect 296732 542406 298067 542408
rect 296732 542404 296738 542406
rect 298001 542403 298067 542406
rect 29126 542268 29132 542332
rect 29196 542330 29202 542332
rect 30097 542330 30163 542333
rect 29196 542328 30163 542330
rect 29196 542272 30102 542328
rect 30158 542272 30163 542328
rect 29196 542270 30163 542272
rect 29196 542268 29202 542270
rect 30097 542267 30163 542270
rect 83733 542330 83799 542333
rect 286961 542330 287027 542333
rect 296294 542330 296300 542332
rect 83733 542328 287027 542330
rect 83733 542272 83738 542328
rect 83794 542272 286966 542328
rect 287022 542272 287027 542328
rect 83733 542270 287027 542272
rect 83733 542267 83799 542270
rect 286961 542267 287027 542270
rect 290782 542270 296300 542330
rect 58382 542132 58388 542196
rect 58452 542194 58458 542196
rect 290782 542194 290842 542270
rect 296294 542268 296300 542270
rect 296364 542268 296370 542332
rect 504541 542330 504607 542333
rect 296670 542328 504607 542330
rect 296670 542272 504546 542328
rect 504602 542272 504607 542328
rect 296670 542270 504607 542272
rect 58452 542134 290842 542194
rect 291009 542194 291075 542197
rect 296670 542194 296730 542270
rect 504541 542267 504607 542270
rect 291009 542192 296730 542194
rect 291009 542136 291014 542192
rect 291070 542136 296730 542192
rect 291009 542134 296730 542136
rect 58452 542132 58458 542134
rect 291009 542131 291075 542134
rect 72601 542058 72667 542061
rect 275829 542058 275895 542061
rect 72601 542056 275895 542058
rect 72601 542000 72606 542056
rect 72662 542000 275834 542056
rect 275890 542000 275895 542056
rect 72601 541998 275895 542000
rect 72601 541995 72667 541998
rect 275829 541995 275895 541998
rect 285254 541996 285260 542060
rect 285324 542058 285330 542060
rect 532734 542058 532740 542060
rect 285324 541998 532740 542058
rect 285324 541996 285330 541998
rect 532734 541996 532740 541998
rect 532804 541996 532810 542060
rect 32622 541860 32628 541924
rect 32692 541922 32698 541924
rect 288566 541922 288572 541924
rect 32692 541862 288572 541922
rect 32692 541860 32698 541862
rect 288566 541860 288572 541862
rect 288636 541860 288642 541924
rect 294454 541860 294460 541924
rect 294524 541922 294530 541924
rect 539726 541922 539732 541924
rect 294524 541862 539732 541922
rect 294524 541860 294530 541862
rect 539726 541860 539732 541862
rect 539796 541860 539802 541924
rect 171542 541724 171548 541788
rect 171612 541786 171618 541788
rect 172421 541786 172487 541789
rect 171612 541784 172487 541786
rect 171612 541728 172426 541784
rect 172482 541728 172487 541784
rect 171612 541726 172487 541728
rect 171612 541724 171618 541726
rect 172421 541723 172487 541726
rect 179229 541786 179295 541789
rect 439773 541786 439839 541789
rect 179229 541784 439839 541786
rect 179229 541728 179234 541784
rect 179290 541728 439778 541784
rect 439834 541728 439839 541784
rect 179229 541726 439839 541728
rect 179229 541723 179295 541726
rect 439773 541723 439839 541726
rect 130285 541650 130351 541653
rect 184197 541650 184263 541653
rect 130285 541648 184263 541650
rect 130285 541592 130290 541648
rect 130346 541592 184202 541648
rect 184258 541592 184263 541648
rect 130285 541590 184263 541592
rect 130285 541587 130351 541590
rect 184197 541587 184263 541590
rect 204805 541650 204871 541653
rect 235993 541650 236059 541653
rect 204805 541648 236059 541650
rect 204805 541592 204810 541648
rect 204866 541592 235998 541648
rect 236054 541592 236059 541648
rect 204805 541590 236059 541592
rect 204805 541587 204871 541590
rect 235993 541587 236059 541590
rect 237189 541650 237255 541653
rect 501137 541650 501203 541653
rect 237189 541648 501203 541650
rect 237189 541592 237194 541648
rect 237250 541592 501142 541648
rect 501198 541592 501203 541648
rect 237189 541590 501203 541592
rect 237189 541587 237255 541590
rect 501137 541587 501203 541590
rect 49233 541514 49299 541517
rect 82813 541514 82879 541517
rect 49233 541512 82879 541514
rect 49233 541456 49238 541512
rect 49294 541456 82818 541512
rect 82874 541456 82879 541512
rect 49233 541454 82879 541456
rect 49233 541451 49299 541454
rect 82813 541451 82879 541454
rect 129273 541514 129339 541517
rect 338573 541514 338639 541517
rect 129273 541512 338639 541514
rect 129273 541456 129278 541512
rect 129334 541456 338578 541512
rect 338634 541456 338639 541512
rect 129273 541454 338639 541456
rect 129273 541451 129339 541454
rect 338573 541451 338639 541454
rect 55765 541378 55831 541381
rect 128353 541378 128419 541381
rect 55765 541376 128419 541378
rect 55765 541320 55770 541376
rect 55826 541320 128358 541376
rect 128414 541320 128419 541376
rect 55765 541318 128419 541320
rect 55765 541315 55831 541318
rect 128353 541315 128419 541318
rect 38193 541242 38259 541245
rect 129733 541242 129799 541245
rect 38193 541240 129799 541242
rect 38193 541184 38198 541240
rect 38254 541184 129738 541240
rect 129794 541184 129799 541240
rect 38193 541182 129799 541184
rect 38193 541179 38259 541182
rect 129733 541179 129799 541182
rect 29678 541044 29684 541108
rect 29748 541106 29754 541108
rect 178033 541106 178099 541109
rect 29748 541104 178099 541106
rect 29748 541048 178038 541104
rect 178094 541048 178099 541104
rect 29748 541046 178099 541048
rect 29748 541044 29754 541046
rect 178033 541043 178099 541046
rect 506473 541106 506539 541109
rect 506790 541106 506796 541108
rect 506473 541104 506796 541106
rect 506473 541048 506478 541104
rect 506534 541048 506796 541104
rect 506473 541046 506796 541048
rect 506473 541043 506539 541046
rect 506790 541044 506796 541046
rect 506860 541044 506866 541108
rect 79685 540970 79751 540973
rect 282913 540970 282979 540973
rect 79685 540968 282979 540970
rect -960 540684 480 540924
rect 79685 540912 79690 540968
rect 79746 540912 282918 540968
rect 282974 540912 282979 540968
rect 79685 540910 282979 540912
rect 79685 540907 79751 540910
rect 282913 540907 282979 540910
rect 295926 540908 295932 540972
rect 295996 540970 296002 540972
rect 502926 540970 502932 540972
rect 295996 540910 502932 540970
rect 295996 540908 296002 540910
rect 502926 540908 502932 540910
rect 502996 540908 503002 540972
rect 107009 540834 107075 540837
rect 316309 540834 316375 540837
rect 107009 540832 316375 540834
rect 107009 540776 107014 540832
rect 107070 540776 316314 540832
rect 316370 540776 316375 540832
rect 107009 540774 316375 540776
rect 107009 540771 107075 540774
rect 316309 540771 316375 540774
rect 73613 540698 73679 540701
rect 276841 540698 276907 540701
rect 73613 540696 276907 540698
rect 73613 540640 73618 540696
rect 73674 540640 276846 540696
rect 276902 540640 276907 540696
rect 73613 540638 276907 540640
rect 73613 540635 73679 540638
rect 276841 540635 276907 540638
rect 298737 540698 298803 540701
rect 510654 540698 510660 540700
rect 298737 540696 510660 540698
rect 298737 540640 298742 540696
rect 298798 540640 510660 540696
rect 298737 540638 510660 540640
rect 298737 540635 298803 540638
rect 510654 540636 510660 540638
rect 510724 540636 510730 540700
rect 170489 540562 170555 540565
rect 175181 540562 175247 540565
rect 170489 540560 175247 540562
rect 170489 540504 170494 540560
rect 170550 540504 175186 540560
rect 175242 540504 175247 540560
rect 170489 540502 175247 540504
rect 170489 540499 170555 540502
rect 175181 540499 175247 540502
rect 175365 540562 175431 540565
rect 428641 540562 428707 540565
rect 175365 540560 428707 540562
rect 175365 540504 175370 540560
rect 175426 540504 428646 540560
rect 428702 540504 428707 540560
rect 175365 540502 428707 540504
rect 175365 540499 175431 540502
rect 428641 540499 428707 540502
rect 58065 540426 58131 540429
rect 247033 540426 247099 540429
rect 58065 540424 247099 540426
rect 58065 540368 58070 540424
rect 58126 540368 247038 540424
rect 247094 540368 247099 540424
rect 58065 540366 247099 540368
rect 58065 540363 58131 540366
rect 247033 540363 247099 540366
rect 218973 540290 219039 540293
rect 244273 540290 244339 540293
rect 218973 540288 244339 540290
rect 218973 540232 218978 540288
rect 219034 540232 244278 540288
rect 244334 540232 244339 540288
rect 218973 540230 244339 540232
rect 218973 540227 219039 540230
rect 244273 540227 244339 540230
rect 247309 540290 247375 540293
rect 512453 540290 512519 540293
rect 247309 540288 512519 540290
rect 247309 540232 247314 540288
rect 247370 540232 512458 540288
rect 512514 540232 512519 540288
rect 247309 540230 512519 540232
rect 247309 540227 247375 540230
rect 512453 540227 512519 540230
rect 91829 540154 91895 540157
rect 295057 540154 295123 540157
rect 91829 540152 295123 540154
rect 91829 540096 91834 540152
rect 91890 540096 295062 540152
rect 295118 540096 295123 540152
rect 91829 540094 295123 540096
rect 91829 540091 91895 540094
rect 295057 540091 295123 540094
rect 50245 540018 50311 540021
rect 91093 540018 91159 540021
rect 50245 540016 91159 540018
rect 50245 539960 50250 540016
rect 50306 539960 91098 540016
rect 91154 539960 91159 540016
rect 50245 539958 91159 539960
rect 50245 539955 50311 539958
rect 91093 539955 91159 539958
rect 245285 540018 245351 540021
rect 507025 540018 507091 540021
rect 245285 540016 507091 540018
rect 245285 539960 245290 540016
rect 245346 539960 507030 540016
rect 507086 539960 507091 540016
rect 245285 539958 507091 539960
rect 245285 539955 245351 539958
rect 507025 539955 507091 539958
rect 32673 539882 32739 539885
rect 107561 539882 107627 539885
rect 32673 539880 107627 539882
rect 32673 539824 32678 539880
rect 32734 539824 107566 539880
rect 107622 539824 107627 539880
rect 32673 539822 107627 539824
rect 32673 539819 32739 539822
rect 107561 539819 107627 539822
rect 36721 539746 36787 539749
rect 169753 539746 169819 539749
rect 521653 539748 521719 539749
rect 521653 539746 521700 539748
rect 36721 539744 169819 539746
rect 36721 539688 36726 539744
rect 36782 539688 169758 539744
rect 169814 539688 169819 539744
rect 36721 539686 169819 539688
rect 521608 539744 521700 539746
rect 521608 539688 521658 539744
rect 521608 539686 521700 539688
rect 36721 539683 36787 539686
rect 169753 539683 169819 539686
rect 521653 539684 521700 539686
rect 521764 539684 521770 539748
rect 521653 539683 521719 539684
rect 33726 539548 33732 539612
rect 33796 539610 33802 539612
rect 218053 539610 218119 539613
rect 33796 539608 218119 539610
rect 33796 539552 218058 539608
rect 218114 539552 218119 539608
rect 33796 539550 218119 539552
rect 33796 539548 33802 539550
rect 218053 539547 218119 539550
rect 222009 539610 222075 539613
rect 225505 539610 225571 539613
rect 222009 539608 225571 539610
rect 222009 539552 222014 539608
rect 222070 539552 225510 539608
rect 225566 539552 225571 539608
rect 222009 539550 225571 539552
rect 222009 539547 222075 539550
rect 225505 539547 225571 539550
rect 521653 539610 521719 539613
rect 521878 539610 521884 539612
rect 521653 539608 521884 539610
rect 521653 539552 521658 539608
rect 521714 539552 521884 539608
rect 521653 539550 521884 539552
rect 521653 539547 521719 539550
rect 521878 539548 521884 539550
rect 521948 539548 521954 539612
rect 57881 539474 57947 539477
rect 104801 539474 104867 539477
rect 57881 539472 104867 539474
rect 57881 539416 57886 539472
rect 57942 539416 104806 539472
rect 104862 539416 104867 539472
rect 57881 539414 104867 539416
rect 57881 539411 57947 539414
rect 104801 539411 104867 539414
rect 350533 539474 350599 539477
rect 500953 539474 501019 539477
rect 350533 539472 501019 539474
rect 350533 539416 350538 539472
rect 350594 539416 500958 539472
rect 501014 539416 501019 539472
rect 350533 539414 501019 539416
rect 350533 539411 350599 539414
rect 500953 539411 501019 539414
rect 85757 539338 85823 539341
rect 288985 539338 289051 539341
rect 85757 539336 289051 539338
rect 85757 539280 85762 539336
rect 85818 539280 288990 539336
rect 289046 539280 289051 539336
rect 85757 539278 289051 539280
rect 85757 539275 85823 539278
rect 288985 539275 289051 539278
rect 290917 539338 290983 539341
rect 522297 539338 522363 539341
rect 290917 539336 522363 539338
rect 290917 539280 290922 539336
rect 290978 539280 522302 539336
rect 522358 539280 522363 539336
rect 290917 539278 522363 539280
rect 290917 539275 290983 539278
rect 522297 539275 522363 539278
rect 61469 539202 61535 539205
rect 253657 539202 253723 539205
rect 61469 539200 253723 539202
rect 61469 539144 61474 539200
rect 61530 539144 253662 539200
rect 253718 539144 253723 539200
rect 61469 539142 253723 539144
rect 61469 539139 61535 539142
rect 253657 539139 253723 539142
rect 282126 539140 282132 539204
rect 282196 539202 282202 539204
rect 514334 539202 514340 539204
rect 282196 539142 514340 539202
rect 282196 539140 282202 539142
rect 514334 539140 514340 539142
rect 514404 539140 514410 539204
rect 103973 539066 104039 539069
rect 226977 539066 227043 539069
rect 103973 539064 227043 539066
rect 103973 539008 103978 539064
rect 104034 539008 226982 539064
rect 227038 539008 227043 539064
rect 103973 539006 227043 539008
rect 103973 539003 104039 539006
rect 226977 539003 227043 539006
rect 253381 539066 253447 539069
rect 508405 539066 508471 539069
rect 253381 539064 508471 539066
rect 253381 539008 253386 539064
rect 253442 539008 508410 539064
rect 508466 539008 508471 539064
rect 253381 539006 508471 539008
rect 253381 539003 253447 539006
rect 508405 539003 508471 539006
rect 59261 538930 59327 538933
rect 352741 538930 352807 538933
rect 59261 538928 352807 538930
rect 59261 538872 59266 538928
rect 59322 538872 352746 538928
rect 352802 538872 352807 538928
rect 59261 538870 352807 538872
rect 59261 538867 59327 538870
rect 352741 538867 352807 538870
rect 49141 538794 49207 538797
rect 60825 538794 60891 538797
rect 49141 538792 60891 538794
rect 49141 538736 49146 538792
rect 49202 538736 60830 538792
rect 60886 538736 60891 538792
rect 49141 538734 60891 538736
rect 49141 538731 49207 538734
rect 60825 538731 60891 538734
rect 225045 538794 225111 538797
rect 522021 538794 522087 538797
rect 225045 538792 522087 538794
rect 225045 538736 225050 538792
rect 225106 538736 522026 538792
rect 522082 538736 522087 538792
rect 225045 538734 522087 538736
rect 225045 538731 225111 538734
rect 522021 538731 522087 538734
rect 35249 538658 35315 538661
rect 86861 538658 86927 538661
rect 35249 538656 86927 538658
rect 35249 538600 35254 538656
rect 35310 538600 86866 538656
rect 86922 538600 86927 538656
rect 35249 538598 86927 538600
rect 35249 538595 35315 538598
rect 86861 538595 86927 538598
rect 135989 538658 136055 538661
rect 254577 538658 254643 538661
rect 135989 538656 254643 538658
rect 135989 538600 135994 538656
rect 136050 538600 254582 538656
rect 254638 538600 254643 538656
rect 135989 538598 254643 538600
rect 135989 538595 136055 538598
rect 254577 538595 254643 538598
rect 295149 538658 295215 538661
rect 502701 538658 502767 538661
rect 295149 538656 502767 538658
rect 295149 538600 295154 538656
rect 295210 538600 502706 538656
rect 502762 538600 502767 538656
rect 295149 538598 502767 538600
rect 295149 538595 295215 538598
rect 502701 538595 502767 538598
rect 26969 538522 27035 538525
rect 100753 538522 100819 538525
rect 26969 538520 100819 538522
rect 26969 538464 26974 538520
rect 27030 538464 100758 538520
rect 100814 538464 100819 538520
rect 26969 538462 100819 538464
rect 26969 538459 27035 538462
rect 100753 538459 100819 538462
rect 101949 538522 102015 538525
rect 311249 538522 311315 538525
rect 101949 538520 311315 538522
rect 101949 538464 101954 538520
rect 102010 538464 311254 538520
rect 311310 538464 311315 538520
rect 101949 538462 311315 538464
rect 101949 538459 102015 538462
rect 311249 538459 311315 538462
rect 54385 538386 54451 538389
rect 136541 538386 136607 538389
rect 54385 538384 136607 538386
rect 54385 538328 54390 538384
rect 54446 538328 136546 538384
rect 136602 538328 136607 538384
rect 54385 538326 136607 538328
rect 54385 538323 54451 538326
rect 136541 538323 136607 538326
rect 44725 538250 44791 538253
rect 222101 538250 222167 538253
rect 44725 538248 222167 538250
rect 44725 538192 44730 538248
rect 44786 538192 222106 538248
rect 222162 538192 222167 538248
rect 44725 538190 222167 538192
rect 44725 538187 44791 538190
rect 222101 538187 222167 538190
rect 58934 538052 58940 538116
rect 59004 538114 59010 538116
rect 109033 538114 109099 538117
rect 59004 538112 109099 538114
rect 59004 538056 109038 538112
rect 109094 538056 109099 538112
rect 59004 538054 109099 538056
rect 59004 538052 59010 538054
rect 109033 538051 109099 538054
rect 110045 537978 110111 537981
rect 319345 537978 319411 537981
rect 110045 537976 319411 537978
rect 110045 537920 110050 537976
rect 110106 537920 319350 537976
rect 319406 537920 319411 537976
rect 110045 537918 319411 537920
rect 110045 537915 110111 537918
rect 319345 537915 319411 537918
rect 68553 537842 68619 537845
rect 270217 537842 270283 537845
rect 68553 537840 270283 537842
rect 68553 537784 68558 537840
rect 68614 537784 270222 537840
rect 270278 537784 270283 537840
rect 68553 537782 270283 537784
rect 68553 537779 68619 537782
rect 270217 537779 270283 537782
rect 283782 537780 283788 537844
rect 283852 537842 283858 537844
rect 534022 537842 534028 537844
rect 283852 537782 534028 537842
rect 283852 537780 283858 537782
rect 534022 537780 534028 537782
rect 534092 537780 534098 537844
rect 580390 537780 580396 537844
rect 580460 537842 580466 537844
rect 583520 537842 584960 537932
rect 580460 537782 584960 537842
rect 580460 537780 580466 537782
rect 31334 537644 31340 537708
rect 31404 537706 31410 537708
rect 286174 537706 286180 537708
rect 31404 537646 286180 537706
rect 31404 537644 31410 537646
rect 286174 537644 286180 537646
rect 286244 537644 286250 537708
rect 290590 537644 290596 537708
rect 290660 537706 290666 537708
rect 520406 537706 520412 537708
rect 290660 537646 520412 537706
rect 290660 537644 290666 537646
rect 520406 537644 520412 537646
rect 520476 537644 520482 537708
rect 583520 537692 584960 537782
rect 166574 537508 166580 537572
rect 166644 537570 166650 537572
rect 166901 537570 166967 537573
rect 166644 537568 166967 537570
rect 166644 537512 166906 537568
rect 166962 537512 166967 537568
rect 166644 537510 166967 537512
rect 166644 537508 166650 537510
rect 166901 537507 166967 537510
rect 252369 537570 252435 537573
rect 512545 537570 512611 537573
rect 252369 537568 512611 537570
rect 252369 537512 252374 537568
rect 252430 537512 512550 537568
rect 512606 537512 512611 537568
rect 252369 537510 512611 537512
rect 252369 537507 252435 537510
rect 512545 537507 512611 537510
rect 35382 537372 35388 537436
rect 35452 537434 35458 537436
rect 379462 537434 379468 537436
rect 35452 537374 379468 537434
rect 35452 537372 35458 537374
rect 379462 537372 379468 537374
rect 379532 537372 379538 537436
rect 84745 537298 84811 537301
rect 287973 537298 288039 537301
rect 84745 537296 288039 537298
rect 84745 537240 84750 537296
rect 84806 537240 287978 537296
rect 288034 537240 288039 537296
rect 84745 537238 288039 537240
rect 84745 537235 84811 537238
rect 287973 537235 288039 537238
rect 49049 537162 49115 537165
rect 85481 537162 85547 537165
rect 49049 537160 85547 537162
rect 49049 537104 49054 537160
rect 49110 537104 85486 537160
rect 85542 537104 85547 537160
rect 49049 537102 85547 537104
rect 49049 537099 49115 537102
rect 85481 537099 85547 537102
rect 116117 537162 116183 537165
rect 325417 537162 325483 537165
rect 116117 537160 325483 537162
rect 116117 537104 116122 537160
rect 116178 537104 325422 537160
rect 325478 537104 325483 537160
rect 116117 537102 325483 537104
rect 116117 537099 116183 537102
rect 325417 537099 325483 537102
rect 35341 537026 35407 537029
rect 117221 537026 117287 537029
rect 35341 537024 117287 537026
rect 35341 536968 35346 537024
rect 35402 536968 117226 537024
rect 117282 536968 117287 537024
rect 35341 536966 117287 536968
rect 35341 536963 35407 536966
rect 117221 536963 117287 536966
rect 40677 536890 40743 536893
rect 252461 536890 252527 536893
rect 40677 536888 252527 536890
rect 40677 536832 40682 536888
rect 40738 536832 252466 536888
rect 252522 536832 252527 536888
rect 40677 536830 252527 536832
rect 40677 536827 40743 536830
rect 252461 536827 252527 536830
rect 59813 536754 59879 536757
rect 299381 536754 299447 536757
rect 59813 536752 299447 536754
rect 59813 536696 59818 536752
rect 59874 536696 299386 536752
rect 299442 536696 299447 536752
rect 59813 536694 299447 536696
rect 59813 536691 59879 536694
rect 299381 536691 299447 536694
rect 416037 536754 416103 536757
rect 436369 536754 436435 536757
rect 416037 536752 436435 536754
rect 416037 536696 416042 536752
rect 416098 536696 436374 536752
rect 436430 536696 436435 536752
rect 416037 536694 436435 536696
rect 416037 536691 416103 536694
rect 436369 536691 436435 536694
rect 169661 536618 169727 536621
rect 231301 536618 231367 536621
rect 169661 536616 231367 536618
rect 169661 536560 169666 536616
rect 169722 536560 231306 536616
rect 231362 536560 231367 536616
rect 169661 536558 231367 536560
rect 169661 536555 169727 536558
rect 231301 536555 231367 536558
rect 233141 536618 233207 536621
rect 241329 536618 241395 536621
rect 233141 536616 241395 536618
rect 233141 536560 233146 536616
rect 233202 536560 241334 536616
rect 241390 536560 241395 536616
rect 233141 536558 241395 536560
rect 233141 536555 233207 536558
rect 241329 536555 241395 536558
rect 298686 536556 298692 536620
rect 298756 536618 298762 536620
rect 518382 536618 518388 536620
rect 298756 536558 518388 536618
rect 298756 536556 298762 536558
rect 518382 536556 518388 536558
rect 518452 536556 518458 536620
rect 90817 536482 90883 536485
rect 294045 536482 294111 536485
rect 90817 536480 294111 536482
rect 90817 536424 90822 536480
rect 90878 536424 294050 536480
rect 294106 536424 294111 536480
rect 90817 536422 294111 536424
rect 90817 536419 90883 536422
rect 294045 536419 294111 536422
rect 299238 536420 299244 536484
rect 299308 536482 299314 536484
rect 526110 536482 526116 536484
rect 299308 536422 526116 536482
rect 299308 536420 299314 536422
rect 526110 536420 526116 536422
rect 526180 536420 526186 536484
rect 76649 536346 76715 536349
rect 279877 536346 279943 536349
rect 76649 536344 279943 536346
rect 76649 536288 76654 536344
rect 76710 536288 279882 536344
rect 279938 536288 279943 536344
rect 76649 536286 279943 536288
rect 76649 536283 76715 536286
rect 279877 536283 279943 536286
rect 291694 536284 291700 536348
rect 291764 536346 291770 536348
rect 519486 536346 519492 536348
rect 291764 536286 519492 536346
rect 291764 536284 291770 536286
rect 519486 536284 519492 536286
rect 519556 536284 519562 536348
rect 57053 536210 57119 536213
rect 175917 536210 175983 536213
rect 57053 536208 175983 536210
rect 57053 536152 57058 536208
rect 57114 536152 175922 536208
rect 175978 536152 175983 536208
rect 57053 536150 175983 536152
rect 57053 536147 57119 536150
rect 175917 536147 175983 536150
rect 241237 536210 241303 536213
rect 504173 536210 504239 536213
rect 241237 536208 504239 536210
rect 241237 536152 241242 536208
rect 241298 536152 504178 536208
rect 504234 536152 504239 536208
rect 241237 536150 504239 536152
rect 241237 536147 241303 536150
rect 504173 536147 504239 536150
rect 176193 536074 176259 536077
rect 444833 536074 444899 536077
rect 176193 536072 444899 536074
rect 176193 536016 176198 536072
rect 176254 536016 444838 536072
rect 444894 536016 444899 536072
rect 176193 536014 444899 536016
rect 176193 536011 176259 536014
rect 444833 536011 444899 536014
rect 465901 536074 465967 536077
rect 517881 536074 517947 536077
rect 465901 536072 517947 536074
rect 465901 536016 465906 536072
rect 465962 536016 517886 536072
rect 517942 536016 517947 536072
rect 465901 536014 517947 536016
rect 465901 536011 465967 536014
rect 517881 536011 517947 536014
rect 48957 535938 49023 535941
rect 89713 535938 89779 535941
rect 48957 535936 89779 535938
rect 48957 535880 48962 535936
rect 49018 535880 89718 535936
rect 89774 535880 89779 535936
rect 48957 535878 89779 535880
rect 48957 535875 49023 535878
rect 89713 535875 89779 535878
rect 109217 535938 109283 535941
rect 318333 535938 318399 535941
rect 109217 535936 318399 535938
rect 109217 535880 109222 535936
rect 109278 535880 318338 535936
rect 318394 535880 318399 535936
rect 109217 535878 318399 535880
rect 109217 535875 109283 535878
rect 318333 535875 318399 535878
rect 58750 535740 58756 535804
rect 58820 535802 58826 535804
rect 117221 535802 117287 535805
rect 326429 535802 326495 535805
rect 58820 535800 117287 535802
rect 58820 535744 117226 535800
rect 117282 535744 117287 535800
rect 58820 535742 117287 535744
rect 58820 535740 58826 535742
rect 117221 535739 117287 535742
rect 122790 535800 326495 535802
rect 122790 535744 326434 535800
rect 326490 535744 326495 535800
rect 122790 535742 326495 535744
rect 32581 535666 32647 535669
rect 109033 535666 109099 535669
rect 32581 535664 109099 535666
rect 32581 535608 32586 535664
rect 32642 535608 109038 535664
rect 109094 535608 109099 535664
rect 32581 535606 109099 535608
rect 32581 535603 32647 535606
rect 109033 535603 109099 535606
rect 117129 535666 117195 535669
rect 122790 535666 122850 535742
rect 326429 535739 326495 535742
rect 117129 535664 122850 535666
rect 117129 535608 117134 535664
rect 117190 535608 122850 535664
rect 117129 535606 122850 535608
rect 117129 535603 117195 535606
rect 39573 535530 39639 535533
rect 168373 535530 168439 535533
rect 39573 535528 168439 535530
rect 39573 535472 39578 535528
rect 39634 535472 168378 535528
rect 168434 535472 168439 535528
rect 39573 535470 168439 535472
rect 39573 535467 39639 535470
rect 168373 535467 168439 535470
rect 535361 535530 535427 535533
rect 535494 535530 535500 535532
rect 535361 535528 535500 535530
rect 535361 535472 535366 535528
rect 535422 535472 535500 535528
rect 535361 535470 535500 535472
rect 535361 535467 535427 535470
rect 535494 535468 535500 535470
rect 535564 535468 535570 535532
rect 108021 535394 108087 535397
rect 317321 535394 317387 535397
rect 108021 535392 317387 535394
rect 108021 535336 108026 535392
rect 108082 535336 317326 535392
rect 317382 535336 317387 535392
rect 108021 535334 317387 535336
rect 108021 535331 108087 535334
rect 317321 535331 317387 535334
rect 100937 535258 101003 535261
rect 310237 535258 310303 535261
rect 100937 535256 310303 535258
rect 100937 535200 100942 535256
rect 100998 535200 310242 535256
rect 310298 535200 310303 535256
rect 100937 535198 310303 535200
rect 100937 535195 101003 535198
rect 310237 535195 310303 535198
rect 62481 535122 62547 535125
rect 265709 535122 265775 535125
rect 62481 535120 265775 535122
rect 62481 535064 62486 535120
rect 62542 535064 265714 535120
rect 265770 535064 265775 535120
rect 62481 535062 265775 535064
rect 62481 535059 62547 535062
rect 265709 535059 265775 535062
rect 295241 535122 295307 535125
rect 521101 535122 521167 535125
rect 295241 535120 521167 535122
rect 295241 535064 295246 535120
rect 295302 535064 521106 535120
rect 521162 535064 521167 535120
rect 295241 535062 521167 535064
rect 295241 535059 295307 535062
rect 521101 535059 521167 535062
rect 38285 534986 38351 534989
rect 255814 534986 255820 534988
rect 38285 534984 255820 534986
rect 38285 534928 38290 534984
rect 38346 534928 255820 534984
rect 38285 534926 255820 534928
rect 38285 534923 38351 534926
rect 255814 534924 255820 534926
rect 255884 534924 255890 534988
rect 285029 534986 285095 534989
rect 515673 534986 515739 534989
rect 285029 534984 515739 534986
rect 285029 534928 285034 534984
rect 285090 534928 515678 534984
rect 515734 534928 515739 534984
rect 285029 534926 515739 534928
rect 285029 534923 285095 534926
rect 515673 534923 515739 534926
rect 57830 534788 57836 534852
rect 57900 534850 57906 534852
rect 108297 534850 108363 534853
rect 57900 534848 108363 534850
rect 57900 534792 108302 534848
rect 108358 534792 108363 534848
rect 57900 534790 108363 534792
rect 57900 534788 57906 534790
rect 108297 534787 108363 534790
rect 250345 534850 250411 534853
rect 512729 534850 512795 534853
rect 250345 534848 512795 534850
rect 250345 534792 250350 534848
rect 250406 534792 512734 534848
rect 512790 534792 512795 534848
rect 250345 534790 512795 534792
rect 250345 534787 250411 534790
rect 512729 534787 512795 534790
rect 170397 534714 170463 534717
rect 464061 534714 464127 534717
rect 170397 534712 464127 534714
rect 170397 534656 170402 534712
rect 170458 534656 464066 534712
rect 464122 534656 464127 534712
rect 170397 534654 464127 534656
rect 170397 534651 170463 534654
rect 464061 534651 464127 534654
rect 89805 534578 89871 534581
rect 293033 534578 293099 534581
rect 89805 534576 293099 534578
rect 89805 534520 89810 534576
rect 89866 534520 293038 534576
rect 293094 534520 293099 534576
rect 89805 534518 293099 534520
rect 89805 534515 89871 534518
rect 293033 534515 293099 534518
rect 299841 534578 299907 534581
rect 502793 534578 502859 534581
rect 299841 534576 502859 534578
rect 299841 534520 299846 534576
rect 299902 534520 502798 534576
rect 502854 534520 502859 534576
rect 299841 534518 502859 534520
rect 299841 534515 299907 534518
rect 502793 534515 502859 534518
rect 58985 534442 59051 534445
rect 100753 534442 100819 534445
rect 58985 534440 100819 534442
rect 58985 534384 58990 534440
rect 59046 534384 100758 534440
rect 100814 534384 100819 534440
rect 58985 534382 100819 534384
rect 58985 534379 59051 534382
rect 100753 534379 100819 534382
rect 46289 534306 46355 534309
rect 169753 534306 169819 534309
rect 46289 534304 169819 534306
rect 46289 534248 46294 534304
rect 46350 534248 169758 534304
rect 169814 534248 169819 534304
rect 46289 534246 169819 534248
rect 46289 534243 46355 534246
rect 169753 534243 169819 534246
rect 27061 534170 27127 534173
rect 251081 534170 251147 534173
rect 27061 534168 251147 534170
rect 27061 534112 27066 534168
rect 27122 534112 251086 534168
rect 251142 534112 251147 534168
rect 27061 534110 251147 534112
rect 27061 534107 27127 534110
rect 251081 534107 251147 534110
rect 499573 534172 499639 534173
rect 499573 534168 499620 534172
rect 499684 534170 499690 534172
rect 499573 534112 499578 534168
rect 499573 534108 499620 534112
rect 499684 534110 499730 534170
rect 499684 534108 499690 534110
rect 499573 534107 499639 534108
rect 115105 534034 115171 534037
rect 324405 534034 324471 534037
rect 115105 534032 324471 534034
rect 115105 533976 115110 534032
rect 115166 533976 324410 534032
rect 324466 533976 324471 534032
rect 115105 533974 324471 533976
rect 115105 533971 115171 533974
rect 324405 533971 324471 533974
rect 478229 534034 478295 534037
rect 535913 534034 535979 534037
rect 478229 534032 535979 534034
rect 478229 533976 478234 534032
rect 478290 533976 535918 534032
rect 535974 533976 535979 534032
rect 478229 533974 535979 533976
rect 478229 533971 478295 533974
rect 535913 533971 535979 533974
rect 105997 533898 106063 533901
rect 315297 533898 315363 533901
rect 105997 533896 315363 533898
rect 105997 533840 106002 533896
rect 106058 533840 315302 533896
rect 315358 533840 315363 533896
rect 105997 533838 315363 533840
rect 105997 533835 106063 533838
rect 315297 533835 315363 533838
rect 471329 533898 471395 533901
rect 533061 533898 533127 533901
rect 471329 533896 533127 533898
rect 471329 533840 471334 533896
rect 471390 533840 533066 533896
rect 533122 533840 533127 533896
rect 471329 533838 533127 533840
rect 471329 533835 471395 533838
rect 533061 533835 533127 533838
rect 34053 533762 34119 533765
rect 259085 533762 259151 533765
rect 34053 533760 259151 533762
rect 34053 533704 34058 533760
rect 34114 533704 259090 533760
rect 259146 533704 259151 533760
rect 34053 533702 259151 533704
rect 34053 533699 34119 533702
rect 259085 533699 259151 533702
rect 287646 533700 287652 533764
rect 287716 533762 287722 533764
rect 498878 533762 498884 533764
rect 287716 533702 498884 533762
rect 287716 533700 287722 533702
rect 498878 533700 498884 533702
rect 498948 533700 498954 533764
rect 500953 533762 501019 533765
rect 518249 533762 518315 533765
rect 500953 533760 518315 533762
rect 500953 533704 500958 533760
rect 501014 533704 518254 533760
rect 518310 533704 518315 533760
rect 500953 533702 518315 533704
rect 500953 533699 501019 533702
rect 518249 533699 518315 533702
rect 44909 533626 44975 533629
rect 292205 533626 292271 533629
rect 44909 533624 292271 533626
rect 44909 533568 44914 533624
rect 44970 533568 292210 533624
rect 292266 533568 292271 533624
rect 44909 533566 292271 533568
rect 44909 533563 44975 533566
rect 292205 533563 292271 533566
rect 465717 533626 465783 533629
rect 536189 533626 536255 533629
rect 465717 533624 536255 533626
rect 465717 533568 465722 533624
rect 465778 533568 536194 533624
rect 536250 533568 536255 533624
rect 465717 533566 536255 533568
rect 465717 533563 465783 533566
rect 536189 533563 536255 533566
rect 175549 533490 175615 533493
rect 429653 533490 429719 533493
rect 175549 533488 429719 533490
rect 175549 533432 175554 533488
rect 175610 533432 429658 533488
rect 429714 533432 429719 533488
rect 175549 533430 429719 533432
rect 175549 533427 175615 533430
rect 429653 533427 429719 533430
rect 463141 533490 463207 533493
rect 534349 533490 534415 533493
rect 463141 533488 534415 533490
rect 463141 533432 463146 533488
rect 463202 533432 534354 533488
rect 534410 533432 534415 533488
rect 463141 533430 534415 533432
rect 463141 533427 463207 533430
rect 534349 533427 534415 533430
rect 51625 533354 51691 533357
rect 106181 533354 106247 533357
rect 51625 533352 106247 533354
rect 51625 533296 51630 533352
rect 51686 533296 106186 533352
rect 106242 533296 106247 533352
rect 51625 533294 106247 533296
rect 51625 533291 51691 533294
rect 106181 533291 106247 533294
rect 223021 533354 223087 533357
rect 504081 533354 504147 533357
rect 223021 533352 504147 533354
rect 223021 533296 223026 533352
rect 223082 533296 504086 533352
rect 504142 533296 504147 533352
rect 223021 533294 504147 533296
rect 223021 533291 223087 533294
rect 504081 533291 504147 533294
rect 65517 533218 65583 533221
rect 224309 533218 224375 533221
rect 65517 533216 224375 533218
rect 65517 533160 65522 533216
rect 65578 533160 224314 533216
rect 224370 533160 224375 533216
rect 65517 533158 224375 533160
rect 65517 533155 65583 533158
rect 224309 533155 224375 533158
rect 485037 533218 485103 533221
rect 533429 533218 533495 533221
rect 485037 533216 533495 533218
rect 485037 533160 485042 533216
rect 485098 533160 533434 533216
rect 533490 533160 533495 533216
rect 485037 533158 533495 533160
rect 485037 533155 485103 533158
rect 533429 533155 533495 533158
rect 36537 533082 36603 533085
rect 115841 533082 115907 533085
rect 36537 533080 115907 533082
rect 36537 533024 36542 533080
rect 36598 533024 115846 533080
rect 115902 533024 115907 533080
rect 36537 533022 115907 533024
rect 36537 533019 36603 533022
rect 115841 533019 115907 533022
rect 475377 533082 475443 533085
rect 485037 533082 485103 533085
rect 475377 533080 485103 533082
rect 475377 533024 475382 533080
rect 475438 533024 485042 533080
rect 485098 533024 485103 533080
rect 475377 533022 485103 533024
rect 475377 533019 475443 533022
rect 485037 533019 485103 533022
rect 31201 532946 31267 532949
rect 175917 532946 175983 532949
rect 31201 532944 175983 532946
rect 31201 532888 31206 532944
rect 31262 532888 175922 532944
rect 175978 532888 175983 532944
rect 31201 532886 175983 532888
rect 31201 532883 31267 532886
rect 175917 532883 175983 532886
rect 40493 532810 40559 532813
rect 223481 532810 223547 532813
rect 40493 532808 223547 532810
rect 40493 532752 40498 532808
rect 40554 532752 223486 532808
rect 223542 532752 223547 532808
rect 40493 532750 223547 532752
rect 40493 532747 40559 532750
rect 223481 532747 223547 532750
rect 509785 532810 509851 532813
rect 514753 532812 514819 532813
rect 518985 532812 519051 532813
rect 510470 532810 510476 532812
rect 509785 532808 510476 532810
rect 509785 532752 509790 532808
rect 509846 532752 510476 532808
rect 509785 532750 510476 532752
rect 509785 532747 509851 532750
rect 510470 532748 510476 532750
rect 510540 532748 510546 532812
rect 514702 532748 514708 532812
rect 514772 532810 514819 532812
rect 514772 532808 514864 532810
rect 514814 532752 514864 532808
rect 514772 532750 514864 532752
rect 514772 532748 514819 532750
rect 518934 532748 518940 532812
rect 519004 532810 519051 532812
rect 519004 532808 519096 532810
rect 519046 532752 519096 532808
rect 519004 532750 519096 532752
rect 519004 532748 519051 532750
rect 514753 532747 514819 532748
rect 518985 532747 519051 532748
rect 177430 532612 177436 532676
rect 177500 532674 177506 532676
rect 177941 532674 178007 532677
rect 177500 532672 178007 532674
rect 177500 532616 177946 532672
rect 178002 532616 178007 532672
rect 177500 532614 178007 532616
rect 177500 532612 177506 532614
rect 177941 532611 178007 532614
rect 215937 532674 216003 532677
rect 512361 532674 512427 532677
rect 215937 532672 512427 532674
rect 215937 532616 215942 532672
rect 215998 532616 512366 532672
rect 512422 532616 512427 532672
rect 215937 532614 512427 532616
rect 215937 532611 216003 532614
rect 512361 532611 512427 532614
rect 59905 532538 59971 532541
rect 356789 532538 356855 532541
rect 59905 532536 356855 532538
rect 59905 532480 59910 532536
rect 59966 532480 356794 532536
rect 356850 532480 356855 532536
rect 59905 532478 356855 532480
rect 59905 532475 59971 532478
rect 356789 532475 356855 532478
rect 436369 532538 436435 532541
rect 440877 532538 440943 532541
rect 436369 532536 440943 532538
rect 436369 532480 436374 532536
rect 436430 532480 440882 532536
rect 440938 532480 440943 532536
rect 436369 532478 440943 532480
rect 436369 532475 436435 532478
rect 440877 532475 440943 532478
rect 56961 532402 57027 532405
rect 375649 532402 375715 532405
rect 56961 532400 375715 532402
rect 56961 532344 56966 532400
rect 57022 532344 375654 532400
rect 375710 532344 375715 532400
rect 56961 532342 375715 532344
rect 56961 532339 57027 532342
rect 375649 532339 375715 532342
rect 57145 532266 57211 532269
rect 378501 532266 378567 532269
rect 57145 532264 378567 532266
rect 57145 532208 57150 532264
rect 57206 532208 378506 532264
rect 378562 532208 378567 532264
rect 57145 532206 378567 532208
rect 57145 532203 57211 532206
rect 378501 532203 378567 532206
rect 57513 532130 57579 532133
rect 378409 532130 378475 532133
rect 57513 532128 378475 532130
rect 57513 532072 57518 532128
rect 57574 532072 378414 532128
rect 378470 532072 378475 532128
rect 57513 532070 378475 532072
rect 57513 532067 57579 532070
rect 378409 532067 378475 532070
rect 37917 531994 37983 531997
rect 386505 531994 386571 531997
rect 37917 531992 386571 531994
rect 37917 531936 37922 531992
rect 37978 531936 386510 531992
rect 386566 531936 386571 531992
rect 37917 531934 386571 531936
rect 37917 531931 37983 531934
rect 386505 531931 386571 531934
rect 52310 531796 52316 531860
rect 52380 531858 52386 531860
rect 296846 531858 296852 531860
rect 52380 531798 296852 531858
rect 52380 531796 52386 531798
rect 296846 531796 296852 531798
rect 296916 531796 296922 531860
rect 57789 531586 57855 531589
rect 59629 531586 59695 531589
rect 57789 531584 59695 531586
rect 57789 531528 57794 531584
rect 57850 531528 59634 531584
rect 59690 531528 59695 531584
rect 57789 531526 59695 531528
rect 57789 531523 57855 531526
rect 59629 531523 59695 531526
rect 57881 531450 57947 531453
rect 215293 531450 215359 531453
rect 57881 531448 215359 531450
rect 57881 531392 57886 531448
rect 57942 531392 215298 531448
rect 215354 531392 215359 531448
rect 57881 531390 215359 531392
rect 57881 531387 57947 531390
rect 215293 531387 215359 531390
rect 499573 531450 499639 531453
rect 499798 531450 499804 531452
rect 499573 531448 499804 531450
rect 499573 531392 499578 531448
rect 499634 531392 499804 531448
rect 499573 531390 499804 531392
rect 499573 531387 499639 531390
rect 499798 531388 499804 531390
rect 499868 531388 499874 531452
rect 521653 531450 521719 531453
rect 525793 531452 525859 531453
rect 522062 531450 522068 531452
rect 521653 531448 522068 531450
rect 521653 531392 521658 531448
rect 521714 531392 522068 531448
rect 521653 531390 522068 531392
rect 521653 531387 521719 531390
rect 522062 531388 522068 531390
rect 522132 531388 522138 531452
rect 525742 531388 525748 531452
rect 525812 531450 525859 531452
rect 529841 531450 529907 531453
rect 529974 531450 529980 531452
rect 525812 531448 525904 531450
rect 525854 531392 525904 531448
rect 525812 531390 525904 531392
rect 529841 531448 529980 531450
rect 529841 531392 529846 531448
rect 529902 531392 529980 531448
rect 529841 531390 529980 531392
rect 525812 531388 525859 531390
rect 525793 531387 525859 531388
rect 529841 531387 529907 531390
rect 529974 531388 529980 531390
rect 530044 531388 530050 531452
rect 137553 531314 137619 531317
rect 175917 531314 175983 531317
rect 137553 531312 175983 531314
rect 137553 531256 137558 531312
rect 137614 531256 175922 531312
rect 175978 531256 175983 531312
rect 137553 531254 175983 531256
rect 137553 531251 137619 531254
rect 175917 531251 175983 531254
rect 179321 531314 179387 531317
rect 436737 531314 436803 531317
rect 179321 531312 436803 531314
rect 179321 531256 179326 531312
rect 179382 531256 436742 531312
rect 436798 531256 436803 531312
rect 179321 531254 436803 531256
rect 179321 531251 179387 531254
rect 436737 531251 436803 531254
rect 163589 531178 163655 531181
rect 178033 531178 178099 531181
rect 163589 531176 178099 531178
rect 163589 531120 163594 531176
rect 163650 531120 178038 531176
rect 178094 531120 178099 531176
rect 163589 531118 178099 531120
rect 163589 531115 163655 531118
rect 178033 531115 178099 531118
rect 179137 531178 179203 531181
rect 437749 531178 437815 531181
rect 179137 531176 437815 531178
rect 179137 531120 179142 531176
rect 179198 531120 437754 531176
rect 437810 531120 437815 531176
rect 179137 531118 437815 531120
rect 179137 531115 179203 531118
rect 437749 531115 437815 531118
rect 137369 531042 137435 531045
rect 164141 531042 164207 531045
rect 137369 531040 164207 531042
rect 137369 530984 137374 531040
rect 137430 530984 164146 531040
rect 164202 530984 164207 531040
rect 137369 530982 164207 530984
rect 137369 530979 137435 530982
rect 164141 530979 164207 530982
rect 178953 531042 179019 531045
rect 438761 531042 438827 531045
rect 178953 531040 438827 531042
rect 178953 530984 178958 531040
rect 179014 530984 438766 531040
rect 438822 530984 438827 531040
rect 178953 530982 438827 530984
rect 178953 530979 179019 530982
rect 438761 530979 438827 530982
rect 166441 530906 166507 530909
rect 173801 530906 173867 530909
rect 166441 530904 173867 530906
rect 166441 530848 166446 530904
rect 166502 530848 173806 530904
rect 173862 530848 173867 530904
rect 166441 530846 173867 530848
rect 166441 530843 166507 530846
rect 173801 530843 173867 530846
rect 176101 530906 176167 530909
rect 440785 530906 440851 530909
rect 176101 530904 440851 530906
rect 176101 530848 176106 530904
rect 176162 530848 440790 530904
rect 440846 530848 440851 530904
rect 176101 530846 440851 530848
rect 176101 530843 176167 530846
rect 440785 530843 440851 530846
rect 482461 530906 482527 530909
rect 516685 530906 516751 530909
rect 482461 530904 516751 530906
rect 482461 530848 482466 530904
rect 482522 530848 516690 530904
rect 516746 530848 516751 530904
rect 482461 530846 516751 530848
rect 482461 530843 482527 530846
rect 516685 530843 516751 530846
rect 33961 530770 34027 530773
rect 310605 530770 310671 530773
rect 33961 530768 310671 530770
rect 33961 530712 33966 530768
rect 34022 530712 310610 530768
rect 310666 530712 310671 530768
rect 33961 530710 310671 530712
rect 33961 530707 34027 530710
rect 310605 530707 310671 530710
rect 461761 530770 461827 530773
rect 526437 530770 526503 530773
rect 461761 530768 526503 530770
rect 461761 530712 461766 530768
rect 461822 530712 526442 530768
rect 526498 530712 526503 530768
rect 461761 530710 526503 530712
rect 461761 530707 461827 530710
rect 526437 530707 526503 530710
rect 41873 530634 41939 530637
rect 153837 530634 153903 530637
rect 41873 530632 153903 530634
rect 41873 530576 41878 530632
rect 41934 530576 153842 530632
rect 153898 530576 153903 530632
rect 41873 530574 153903 530576
rect 41873 530571 41939 530574
rect 153837 530571 153903 530574
rect 162117 530634 162183 530637
rect 459001 530634 459067 530637
rect 162117 530632 459067 530634
rect 162117 530576 162122 530632
rect 162178 530576 459006 530632
rect 459062 530576 459067 530632
rect 162117 530574 459067 530576
rect 162117 530571 162183 530574
rect 459001 530571 459067 530574
rect 467281 530634 467347 530637
rect 533521 530634 533587 530637
rect 467281 530632 533587 530634
rect 467281 530576 467286 530632
rect 467342 530576 533526 530632
rect 533582 530576 533587 530632
rect 467281 530574 533587 530576
rect 467281 530571 467347 530574
rect 533521 530571 533587 530574
rect 61878 530436 61884 530500
rect 61948 530498 61954 530500
rect 137185 530498 137251 530501
rect 61948 530496 137251 530498
rect 61948 530440 137190 530496
rect 137246 530440 137251 530496
rect 61948 530438 137251 530440
rect 61948 530436 61954 530438
rect 137185 530435 137251 530438
rect 173341 530498 173407 530501
rect 256693 530498 256759 530501
rect 173341 530496 256759 530498
rect 173341 530440 173346 530496
rect 173402 530440 256698 530496
rect 256754 530440 256759 530496
rect 173341 530438 256759 530440
rect 173341 530435 173407 530438
rect 256693 530435 256759 530438
rect 257889 530498 257955 530501
rect 507301 530498 507367 530501
rect 257889 530496 507367 530498
rect 257889 530440 257894 530496
rect 257950 530440 507306 530496
rect 507362 530440 507367 530496
rect 257889 530438 507367 530440
rect 257889 530435 257955 530438
rect 507301 530435 507367 530438
rect 50838 530300 50844 530364
rect 50908 530362 50914 530364
rect 135161 530362 135227 530365
rect 50908 530360 135227 530362
rect 50908 530304 135166 530360
rect 135222 530304 135227 530360
rect 50908 530302 135227 530304
rect 50908 530300 50914 530302
rect 135161 530299 135227 530302
rect 43846 530164 43852 530228
rect 43916 530226 43922 530228
rect 166165 530226 166231 530229
rect 43916 530224 166231 530226
rect 43916 530168 166170 530224
rect 166226 530168 166231 530224
rect 43916 530166 166231 530168
rect 43916 530164 43922 530166
rect 166165 530163 166231 530166
rect 40585 530090 40651 530093
rect 178217 530090 178283 530093
rect 40585 530088 178283 530090
rect 40585 530032 40590 530088
rect 40646 530032 178222 530088
rect 178278 530032 178283 530088
rect 40585 530030 178283 530032
rect 40585 530027 40651 530030
rect 178217 530027 178283 530030
rect 36670 529892 36676 529956
rect 36740 529954 36746 529956
rect 178125 529954 178191 529957
rect 36740 529952 178191 529954
rect 36740 529896 178130 529952
rect 178186 529896 178191 529952
rect 36740 529894 178191 529896
rect 36740 529892 36746 529894
rect 178125 529891 178191 529894
rect 53741 529820 53807 529821
rect 53741 529816 53788 529820
rect 53852 529818 53858 529820
rect 58433 529818 58499 529821
rect 299381 529818 299447 529821
rect 53741 529760 53746 529816
rect 53741 529756 53788 529760
rect 53852 529758 53898 529818
rect 58433 529816 299447 529818
rect 58433 529760 58438 529816
rect 58494 529760 299386 529816
rect 299442 529760 299447 529816
rect 58433 529758 299447 529760
rect 53852 529756 53858 529758
rect 53741 529755 53807 529756
rect 58433 529755 58499 529758
rect 299381 529755 299447 529758
rect 95877 529682 95943 529685
rect 306189 529682 306255 529685
rect 95877 529680 306255 529682
rect 95877 529624 95882 529680
rect 95938 529624 306194 529680
rect 306250 529624 306255 529680
rect 95877 529622 306255 529624
rect 95877 529619 95943 529622
rect 306189 529619 306255 529622
rect 93853 529546 93919 529549
rect 95509 529546 95575 529549
rect 93853 529544 95575 529546
rect 93853 529488 93858 529544
rect 93914 529488 95514 529544
rect 95570 529488 95575 529544
rect 93853 529486 95575 529488
rect 93853 529483 93919 529486
rect 95509 529483 95575 529486
rect 286358 529484 286364 529548
rect 286428 529546 286434 529548
rect 497590 529546 497596 529548
rect 286428 529486 497596 529546
rect 286428 529484 286434 529486
rect 497590 529484 497596 529486
rect 497660 529484 497666 529548
rect 61326 529348 61332 529412
rect 61396 529410 61402 529412
rect 96521 529410 96587 529413
rect 61396 529408 96587 529410
rect 61396 529352 96526 529408
rect 96582 529352 96587 529408
rect 61396 529350 96587 529352
rect 61396 529348 61402 529350
rect 96521 529347 96587 529350
rect 299289 529410 299355 529413
rect 525149 529410 525215 529413
rect 299289 529408 525215 529410
rect 299289 529352 299294 529408
rect 299350 529352 525154 529408
rect 525210 529352 525215 529408
rect 299289 529350 525215 529352
rect 299289 529347 299355 529350
rect 525149 529347 525215 529350
rect 58617 529274 58683 529277
rect 347681 529274 347747 529277
rect 58617 529272 347747 529274
rect 58617 529216 58622 529272
rect 58678 529216 347686 529272
rect 347742 529216 347747 529272
rect 58617 529214 347747 529216
rect 58617 529211 58683 529214
rect 347681 529211 347747 529214
rect 500953 529274 501019 529277
rect 501270 529274 501276 529276
rect 500953 529272 501276 529274
rect 500953 529216 500958 529272
rect 501014 529216 501276 529272
rect 500953 529214 501276 529216
rect 500953 529211 501019 529214
rect 501270 529212 501276 529214
rect 501340 529212 501346 529276
rect 58893 529138 58959 529141
rect 363873 529138 363939 529141
rect 58893 529136 363939 529138
rect 58893 529080 58898 529136
rect 58954 529080 363878 529136
rect 363934 529080 363939 529136
rect 58893 529078 363939 529080
rect 58893 529075 58959 529078
rect 363873 529075 363939 529078
rect 450486 529076 450492 529140
rect 450556 529138 450562 529140
rect 514017 529138 514083 529141
rect 450556 529136 514083 529138
rect 450556 529080 514022 529136
rect 514078 529080 514083 529136
rect 450556 529078 514083 529080
rect 450556 529076 450562 529078
rect 514017 529075 514083 529078
rect 51717 529002 51783 529005
rect 95141 529002 95207 529005
rect 305177 529002 305243 529005
rect 51717 529000 95207 529002
rect 51717 528944 51722 529000
rect 51778 528944 95146 529000
rect 95202 528944 95207 529000
rect 51717 528942 95207 528944
rect 51717 528939 51783 528942
rect 95141 528939 95207 528942
rect 95374 529000 305243 529002
rect 95374 528944 305182 529000
rect 305238 528944 305243 529000
rect 95374 528942 305243 528944
rect 94865 528866 94931 528869
rect 95374 528866 95434 528942
rect 305177 528939 305243 528942
rect 94865 528864 95434 528866
rect 94865 528808 94870 528864
rect 94926 528808 95434 528864
rect 94865 528806 95434 528808
rect 95509 528866 95575 528869
rect 302233 528866 302299 528869
rect 95509 528864 302299 528866
rect 95509 528808 95514 528864
rect 95570 528808 302238 528864
rect 302294 528808 302299 528864
rect 95509 528806 302299 528808
rect 94865 528803 94931 528806
rect 95509 528803 95575 528806
rect 302233 528803 302299 528806
rect 44817 528730 44883 528733
rect 95049 528730 95115 528733
rect 44817 528728 95115 528730
rect 44817 528672 44822 528728
rect 44878 528672 95054 528728
rect 95110 528672 95115 528728
rect 44817 528670 95115 528672
rect 44817 528667 44883 528670
rect 95049 528667 95115 528670
rect 42558 528532 42564 528596
rect 42628 528594 42634 528596
rect 285673 528594 285739 528597
rect 42628 528592 285739 528594
rect 42628 528536 285678 528592
rect 285734 528536 285739 528592
rect 42628 528534 285739 528536
rect 42628 528532 42634 528534
rect 285673 528531 285739 528534
rect 500953 528594 501019 528597
rect 501638 528594 501644 528596
rect 500953 528592 501644 528594
rect 500953 528536 500958 528592
rect 501014 528536 501644 528592
rect 500953 528534 501644 528536
rect 500953 528531 501019 528534
rect 501638 528532 501644 528534
rect 501708 528532 501714 528596
rect 122189 528458 122255 528461
rect 331489 528458 331555 528461
rect 122189 528456 331555 528458
rect 122189 528400 122194 528456
rect 122250 528400 331494 528456
rect 331550 528400 331555 528456
rect 122189 528398 331555 528400
rect 122189 528395 122255 528398
rect 331489 528395 331555 528398
rect 440877 528458 440943 528461
rect 444281 528458 444347 528461
rect 440877 528456 444347 528458
rect 440877 528400 440882 528456
rect 440938 528400 444286 528456
rect 444342 528400 444347 528456
rect 440877 528398 444347 528400
rect 440877 528395 440943 528398
rect 444281 528395 444347 528398
rect 123201 528322 123267 528325
rect 332317 528322 332383 528325
rect 123201 528320 332383 528322
rect 123201 528264 123206 528320
rect 123262 528264 332322 528320
rect 332378 528264 332383 528320
rect 123201 528262 332383 528264
rect 123201 528259 123267 528262
rect 332317 528259 332383 528262
rect 487981 528322 488047 528325
rect 531865 528322 531931 528325
rect 487981 528320 531931 528322
rect 487981 528264 487986 528320
rect 488042 528264 531870 528320
rect 531926 528264 531931 528320
rect 487981 528262 531931 528264
rect 487981 528259 488047 528262
rect 531865 528259 531931 528262
rect 25998 528124 26004 528188
rect 26068 528186 26074 528188
rect 125501 528186 125567 528189
rect 26068 528184 125567 528186
rect 26068 528128 125506 528184
rect 125562 528128 125567 528184
rect 26068 528126 125567 528128
rect 26068 528124 26074 528126
rect 125501 528123 125567 528126
rect 468477 528186 468543 528189
rect 527725 528186 527791 528189
rect 468477 528184 527791 528186
rect 468477 528128 468482 528184
rect 468538 528128 527730 528184
rect 527786 528128 527791 528184
rect 468477 528126 527791 528128
rect 468477 528123 468543 528126
rect 527725 528123 527791 528126
rect 80789 528050 80855 528053
rect 120073 528050 120139 528053
rect 80789 528048 120139 528050
rect -960 527914 480 528004
rect 80789 527992 80794 528048
rect 80850 527992 120078 528048
rect 120134 527992 120139 528048
rect 80789 527990 120139 527992
rect 80789 527987 80855 527990
rect 120073 527987 120139 527990
rect 121177 528050 121243 528053
rect 330385 528050 330451 528053
rect 121177 528048 330451 528050
rect 121177 527992 121182 528048
rect 121238 527992 330390 528048
rect 330446 527992 330451 528048
rect 121177 527990 330451 527992
rect 121177 527987 121243 527990
rect 330385 527987 330451 527990
rect 476614 527988 476620 528052
rect 476684 528050 476690 528052
rect 536782 528050 536788 528052
rect 476684 527990 536788 528050
rect 476684 527988 476690 527990
rect 536782 527988 536788 527990
rect 536852 527988 536858 528052
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 120165 527914 120231 527917
rect 329373 527914 329439 527917
rect 120165 527912 329439 527914
rect 120165 527856 120170 527912
rect 120226 527856 329378 527912
rect 329434 527856 329439 527912
rect 120165 527854 329439 527856
rect 120165 527851 120231 527854
rect 329373 527851 329439 527854
rect 467189 527914 467255 527917
rect 531773 527914 531839 527917
rect 467189 527912 531839 527914
rect 467189 527856 467194 527912
rect 467250 527856 531778 527912
rect 531834 527856 531839 527912
rect 467189 527854 531839 527856
rect 467189 527851 467255 527854
rect 531773 527851 531839 527854
rect 102961 527778 103027 527781
rect 312169 527778 312235 527781
rect 102961 527776 312235 527778
rect 102961 527720 102966 527776
rect 103022 527720 312174 527776
rect 312230 527720 312235 527776
rect 102961 527718 312235 527720
rect 102961 527715 103027 527718
rect 312169 527715 312235 527718
rect 467373 527778 467439 527781
rect 534809 527778 534875 527781
rect 467373 527776 534875 527778
rect 467373 527720 467378 527776
rect 467434 527720 534814 527776
rect 534870 527720 534875 527776
rect 467373 527718 534875 527720
rect 467373 527715 467439 527718
rect 534809 527715 534875 527718
rect 43253 527642 43319 527645
rect 121453 527642 121519 527645
rect 43253 527640 121519 527642
rect 43253 527584 43258 527640
rect 43314 527584 121458 527640
rect 121514 527584 121519 527640
rect 43253 527582 121519 527584
rect 43253 527579 43319 527582
rect 121453 527579 121519 527582
rect 125225 527642 125291 527645
rect 334525 527642 334591 527645
rect 125225 527640 334591 527642
rect 125225 527584 125230 527640
rect 125286 527584 334530 527640
rect 334586 527584 334591 527640
rect 125225 527582 334591 527584
rect 125225 527579 125291 527582
rect 334525 527579 334591 527582
rect 44173 527506 44239 527509
rect 125409 527506 125475 527509
rect 44173 527504 125475 527506
rect 44173 527448 44178 527504
rect 44234 527448 125414 527504
rect 125470 527448 125475 527504
rect 44173 527446 125475 527448
rect 44173 527443 44239 527446
rect 125409 527443 125475 527446
rect 39389 527370 39455 527373
rect 124121 527370 124187 527373
rect 39389 527368 124187 527370
rect 39389 527312 39394 527368
rect 39450 527312 124126 527368
rect 124182 527312 124187 527368
rect 39389 527310 124187 527312
rect 39389 527307 39455 527310
rect 124121 527307 124187 527310
rect 124581 527370 124647 527373
rect 333421 527370 333487 527373
rect 124581 527368 333487 527370
rect 124581 527312 124586 527368
rect 124642 527312 333426 527368
rect 333482 527312 333487 527368
rect 124581 527310 333487 527312
rect 124581 527307 124647 527310
rect 333421 527307 333487 527310
rect 49734 527172 49740 527236
rect 49804 527234 49810 527236
rect 50981 527234 51047 527237
rect 55121 527236 55187 527237
rect 55070 527234 55076 527236
rect 49804 527232 51047 527234
rect 49804 527176 50986 527232
rect 51042 527176 51047 527232
rect 49804 527174 51047 527176
rect 55030 527174 55076 527234
rect 55140 527232 55187 527236
rect 55182 527176 55187 527232
rect 49804 527172 49810 527174
rect 50981 527171 51047 527174
rect 55070 527172 55076 527174
rect 55140 527172 55187 527176
rect 55121 527171 55187 527172
rect 59629 527234 59695 527237
rect 120901 527234 120967 527237
rect 511993 527236 512059 527237
rect 59629 527232 120967 527234
rect 59629 527176 59634 527232
rect 59690 527176 120906 527232
rect 120962 527176 120967 527232
rect 59629 527174 120967 527176
rect 59629 527171 59695 527174
rect 120901 527171 120967 527174
rect 511942 527172 511948 527236
rect 512012 527234 512059 527236
rect 514753 527234 514819 527237
rect 514886 527234 514892 527236
rect 512012 527232 512104 527234
rect 512054 527176 512104 527232
rect 512012 527174 512104 527176
rect 514753 527232 514892 527234
rect 514753 527176 514758 527232
rect 514814 527176 514892 527232
rect 514753 527174 514892 527176
rect 512012 527172 512059 527174
rect 511993 527171 512059 527172
rect 514753 527171 514819 527174
rect 514886 527172 514892 527174
rect 514956 527172 514962 527236
rect 517513 527234 517579 527237
rect 518014 527234 518020 527236
rect 517513 527232 518020 527234
rect 517513 527176 517518 527232
rect 517574 527176 518020 527232
rect 517513 527174 518020 527176
rect 517513 527171 517579 527174
rect 518014 527172 518020 527174
rect 518084 527172 518090 527236
rect 523033 527234 523099 527237
rect 523534 527234 523540 527236
rect 523033 527232 523540 527234
rect 523033 527176 523038 527232
rect 523094 527176 523540 527232
rect 523033 527174 523540 527176
rect 523033 527171 523099 527174
rect 523534 527172 523540 527174
rect 523604 527172 523610 527236
rect 113081 527098 113147 527101
rect 322381 527098 322447 527101
rect 113081 527096 322447 527098
rect 113081 527040 113086 527096
rect 113142 527040 322386 527096
rect 322442 527040 322447 527096
rect 113081 527038 322447 527040
rect 113081 527035 113147 527038
rect 322381 527035 322447 527038
rect 479609 527098 479675 527101
rect 531957 527098 532023 527101
rect 479609 527096 532023 527098
rect 479609 527040 479614 527096
rect 479670 527040 531962 527096
rect 532018 527040 532023 527096
rect 479609 527038 532023 527040
rect 479609 527035 479675 527038
rect 531957 527035 532023 527038
rect 32489 526962 32555 526965
rect 106181 526962 106247 526965
rect 32489 526960 106247 526962
rect 32489 526904 32494 526960
rect 32550 526904 106186 526960
rect 106242 526904 106247 526960
rect 32489 526902 106247 526904
rect 32489 526899 32555 526902
rect 106181 526899 106247 526902
rect 214925 526962 214991 526965
rect 237465 526962 237531 526965
rect 214925 526960 237531 526962
rect 214925 526904 214930 526960
rect 214986 526904 237470 526960
rect 237526 526904 237531 526960
rect 214925 526902 237531 526904
rect 214925 526899 214991 526902
rect 237465 526899 237531 526902
rect 238201 526962 238267 526965
rect 288341 526962 288407 526965
rect 512310 526962 512316 526964
rect 238201 526960 288407 526962
rect 238201 526904 238206 526960
rect 238262 526904 288346 526960
rect 288402 526904 288407 526960
rect 238201 526902 288407 526904
rect 238201 526899 238267 526902
rect 288341 526899 288407 526902
rect 291334 526902 512316 526962
rect 44950 526764 44956 526828
rect 45020 526826 45026 526828
rect 291142 526826 291148 526828
rect 45020 526766 291148 526826
rect 45020 526764 45026 526766
rect 291142 526764 291148 526766
rect 291212 526764 291218 526828
rect 51533 526690 51599 526693
rect 62021 526690 62087 526693
rect 51533 526688 62087 526690
rect 51533 526632 51538 526688
rect 51594 526632 62026 526688
rect 62082 526632 62087 526688
rect 51533 526630 62087 526632
rect 51533 526627 51599 526630
rect 62021 526627 62087 526630
rect 234153 526690 234219 526693
rect 256693 526690 256759 526693
rect 234153 526688 256759 526690
rect 234153 526632 234158 526688
rect 234214 526632 256698 526688
rect 256754 526632 256759 526688
rect 234153 526630 256759 526632
rect 234153 526627 234219 526630
rect 256693 526627 256759 526630
rect 288014 526628 288020 526692
rect 288084 526690 288090 526692
rect 291334 526690 291394 526902
rect 512310 526900 512316 526902
rect 512380 526900 512386 526964
rect 296110 526764 296116 526828
rect 296180 526826 296186 526828
rect 502742 526826 502748 526828
rect 296180 526766 502748 526826
rect 296180 526764 296186 526766
rect 502742 526764 502748 526766
rect 502812 526764 502818 526828
rect 288084 526630 291394 526690
rect 288084 526628 288090 526630
rect 35157 526554 35223 526557
rect 111793 526554 111859 526557
rect 35157 526552 111859 526554
rect 35157 526496 35162 526552
rect 35218 526496 111798 526552
rect 111854 526496 111859 526552
rect 35157 526494 111859 526496
rect 35157 526491 35223 526494
rect 111793 526491 111859 526494
rect 178861 526554 178927 526557
rect 441705 526554 441771 526557
rect 178861 526552 441771 526554
rect 178861 526496 178866 526552
rect 178922 526496 441710 526552
rect 441766 526496 441771 526552
rect 178861 526494 441771 526496
rect 178861 526491 178927 526494
rect 441705 526491 441771 526494
rect 444281 526554 444347 526557
rect 501454 526554 501460 526556
rect 444281 526552 501460 526554
rect 444281 526496 444286 526552
rect 444342 526496 501460 526552
rect 444281 526494 501460 526496
rect 444281 526491 444347 526494
rect 501454 526492 501460 526494
rect 501524 526492 501530 526556
rect 518249 526554 518315 526557
rect 544561 526554 544627 526557
rect 518249 526552 544627 526554
rect 518249 526496 518254 526552
rect 518310 526496 544566 526552
rect 544622 526496 544627 526552
rect 518249 526494 544627 526496
rect 518249 526491 518315 526494
rect 544561 526491 544627 526494
rect 57053 526418 57119 526421
rect 178033 526418 178099 526421
rect 57053 526416 178099 526418
rect 57053 526360 57058 526416
rect 57114 526360 178038 526416
rect 178094 526360 178099 526416
rect 57053 526358 178099 526360
rect 57053 526355 57119 526358
rect 178033 526355 178099 526358
rect 249333 526418 249399 526421
rect 519537 526418 519603 526421
rect 249333 526416 519603 526418
rect 249333 526360 249338 526416
rect 249394 526360 519542 526416
rect 519598 526360 519603 526416
rect 249333 526358 519603 526360
rect 249333 526355 249399 526358
rect 519537 526355 519603 526358
rect 104985 526282 105051 526285
rect 298001 526282 298067 526285
rect 104985 526280 298067 526282
rect 104985 526224 104990 526280
rect 105046 526224 298006 526280
rect 298062 526224 298067 526280
rect 104985 526222 298067 526224
rect 104985 526219 105051 526222
rect 298001 526219 298067 526222
rect 61745 526146 61811 526149
rect 214557 526146 214623 526149
rect 61745 526144 214623 526146
rect 61745 526088 61750 526144
rect 61806 526088 214562 526144
rect 214618 526088 214623 526144
rect 61745 526086 214623 526088
rect 61745 526083 61811 526086
rect 214557 526083 214623 526086
rect 257102 526084 257108 526148
rect 257172 526146 257178 526148
rect 514518 526146 514524 526148
rect 257172 526086 514524 526146
rect 257172 526084 257178 526086
rect 514518 526084 514524 526086
rect 514588 526084 514594 526148
rect 35198 525948 35204 526012
rect 35268 526010 35274 526012
rect 233877 526010 233943 526013
rect 35268 526008 233943 526010
rect 35268 525952 233882 526008
rect 233938 525952 233943 526008
rect 35268 525950 233943 525952
rect 35268 525948 35274 525950
rect 233877 525947 233943 525950
rect 41086 525812 41092 525876
rect 41156 525874 41162 525876
rect 249701 525874 249767 525877
rect 41156 525872 249767 525874
rect 41156 525816 249706 525872
rect 249762 525816 249767 525872
rect 41156 525814 249767 525816
rect 41156 525812 41162 525814
rect 249701 525811 249767 525814
rect 514201 525874 514267 525877
rect 514334 525874 514340 525876
rect 514201 525872 514340 525874
rect 514201 525816 514206 525872
rect 514262 525816 514340 525872
rect 514201 525814 514340 525816
rect 514201 525811 514267 525814
rect 514334 525812 514340 525814
rect 514404 525812 514410 525876
rect 177614 525676 177620 525740
rect 177684 525738 177690 525740
rect 177941 525738 178007 525741
rect 177684 525736 178007 525738
rect 177684 525680 177946 525736
rect 178002 525680 178007 525736
rect 177684 525678 178007 525680
rect 177684 525676 177690 525678
rect 177941 525675 178007 525678
rect 487797 525738 487863 525741
rect 523677 525738 523743 525741
rect 487797 525736 523743 525738
rect 487797 525680 487802 525736
rect 487858 525680 523682 525736
rect 523738 525680 523743 525736
rect 487797 525678 523743 525680
rect 487797 525675 487863 525678
rect 523677 525675 523743 525678
rect 69565 525602 69631 525605
rect 272701 525602 272767 525605
rect 69565 525600 272767 525602
rect 69565 525544 69570 525600
rect 69626 525544 272706 525600
rect 272762 525544 272767 525600
rect 69565 525542 272767 525544
rect 69565 525539 69631 525542
rect 272701 525539 272767 525542
rect 280654 525540 280660 525604
rect 280724 525602 280730 525604
rect 499430 525602 499436 525604
rect 280724 525542 499436 525602
rect 280724 525540 280730 525542
rect 499430 525540 499436 525542
rect 499500 525540 499506 525604
rect 44766 525404 44772 525468
rect 44836 525466 44842 525468
rect 289118 525466 289124 525468
rect 44836 525406 289124 525466
rect 44836 525404 44842 525406
rect 289118 525404 289124 525406
rect 289188 525404 289194 525468
rect 296621 525466 296687 525469
rect 503069 525466 503135 525469
rect 296621 525464 503135 525466
rect 296621 525408 296626 525464
rect 296682 525408 503074 525464
rect 503130 525408 503135 525464
rect 296621 525406 503135 525408
rect 296621 525403 296687 525406
rect 503069 525403 503135 525406
rect 70577 525330 70643 525333
rect 273805 525330 273871 525333
rect 70577 525328 273871 525330
rect 70577 525272 70582 525328
rect 70638 525272 273810 525328
rect 273866 525272 273871 525328
rect 70577 525270 273871 525272
rect 70577 525267 70643 525270
rect 273805 525267 273871 525270
rect 285070 525268 285076 525332
rect 285140 525330 285146 525332
rect 530158 525330 530164 525332
rect 285140 525270 530164 525330
rect 285140 525268 285146 525270
rect 530158 525268 530164 525270
rect 530228 525268 530234 525332
rect 31109 525194 31175 525197
rect 44173 525194 44239 525197
rect 31109 525192 44239 525194
rect 31109 525136 31114 525192
rect 31170 525136 44178 525192
rect 44234 525136 44239 525192
rect 31109 525134 44239 525136
rect 31109 525131 31175 525134
rect 44173 525131 44239 525134
rect 46422 525132 46428 525196
rect 46492 525194 46498 525196
rect 282862 525194 282868 525196
rect 46492 525134 282868 525194
rect 46492 525132 46498 525134
rect 282862 525132 282868 525134
rect 282932 525132 282938 525196
rect 285438 525132 285444 525196
rect 285508 525194 285514 525196
rect 535678 525194 535684 525196
rect 285508 525134 535684 525194
rect 285508 525132 285514 525134
rect 535678 525132 535684 525134
rect 535748 525132 535754 525196
rect 41270 524996 41276 525060
rect 41340 525058 41346 525060
rect 69013 525058 69079 525061
rect 41340 525056 69079 525058
rect 41340 525000 69018 525056
rect 69074 525000 69079 525056
rect 41340 524998 69079 525000
rect 41340 524996 41346 524998
rect 69013 524995 69079 524998
rect 248321 525058 248387 525061
rect 507117 525058 507183 525061
rect 248321 525056 507183 525058
rect 248321 525000 248326 525056
rect 248382 525000 507122 525056
rect 507178 525000 507183 525056
rect 248321 524998 507183 525000
rect 248321 524995 248387 524998
rect 507117 524995 507183 524998
rect 36486 524860 36492 524924
rect 36556 524922 36562 524924
rect 70393 524922 70459 524925
rect 36556 524920 70459 524922
rect 36556 524864 70398 524920
rect 70454 524864 70459 524920
rect 36556 524862 70459 524864
rect 36556 524860 36562 524862
rect 70393 524859 70459 524862
rect 118141 524922 118207 524925
rect 225321 524922 225387 524925
rect 258073 524922 258139 524925
rect 118141 524920 122850 524922
rect 118141 524864 118146 524920
rect 118202 524864 122850 524920
rect 118141 524862 122850 524864
rect 118141 524859 118207 524862
rect 42374 524724 42380 524788
rect 42444 524786 42450 524788
rect 117957 524786 118023 524789
rect 42444 524784 118023 524786
rect 42444 524728 117962 524784
rect 118018 524728 118023 524784
rect 42444 524726 118023 524728
rect 122790 524786 122850 524862
rect 225321 524920 258139 524922
rect 225321 524864 225326 524920
rect 225382 524864 258078 524920
rect 258134 524864 258139 524920
rect 225321 524862 258139 524864
rect 225321 524859 225387 524862
rect 258073 524859 258139 524862
rect 327349 524786 327415 524789
rect 122790 524784 327415 524786
rect 122790 524728 327354 524784
rect 327410 524728 327415 524784
rect 122790 524726 327415 524728
rect 42444 524724 42450 524726
rect 117957 524723 118023 524726
rect 327349 524723 327415 524726
rect 35433 524650 35499 524653
rect 224953 524650 225019 524653
rect 35433 524648 225019 524650
rect 35433 524592 35438 524648
rect 35494 524592 224958 524648
rect 225014 524592 225019 524648
rect 35433 524590 225019 524592
rect 35433 524587 35499 524590
rect 224953 524587 225019 524590
rect 39430 524452 39436 524516
rect 39500 524514 39506 524516
rect 247033 524514 247099 524517
rect 39500 524512 247099 524514
rect 39500 524456 247038 524512
rect 247094 524456 247099 524512
rect 39500 524454 247099 524456
rect 39500 524452 39506 524454
rect 247033 524451 247099 524454
rect 511993 524514 512059 524517
rect 512494 524514 512500 524516
rect 511993 524512 512500 524514
rect 511993 524456 511998 524512
rect 512054 524456 512500 524512
rect 511993 524454 512500 524456
rect 511993 524451 512059 524454
rect 512494 524452 512500 524454
rect 512564 524452 512570 524516
rect 548374 524452 548380 524516
rect 548444 524514 548450 524516
rect 583520 524514 584960 524604
rect 548444 524454 584960 524514
rect 548444 524452 548450 524454
rect 54702 524316 54708 524380
rect 54772 524378 54778 524380
rect 296478 524378 296484 524380
rect 54772 524318 296484 524378
rect 54772 524316 54778 524318
rect 296478 524316 296484 524318
rect 296548 524316 296554 524380
rect 480294 524316 480300 524380
rect 480364 524378 480370 524380
rect 481541 524378 481607 524381
rect 480364 524376 481607 524378
rect 480364 524320 481546 524376
rect 481602 524320 481607 524376
rect 583520 524364 584960 524454
rect 480364 524318 481607 524320
rect 480364 524316 480370 524318
rect 481541 524315 481607 524318
rect 68277 524242 68343 524245
rect 267733 524242 267799 524245
rect 68277 524240 267799 524242
rect 68277 524184 68282 524240
rect 68338 524184 267738 524240
rect 267794 524184 267799 524240
rect 68277 524182 267799 524184
rect 68277 524179 68343 524182
rect 267733 524179 267799 524182
rect 281022 524180 281028 524244
rect 281092 524242 281098 524244
rect 527398 524242 527404 524244
rect 281092 524182 527404 524242
rect 281092 524180 281098 524182
rect 527398 524180 527404 524182
rect 527468 524180 527474 524244
rect 37406 524044 37412 524108
rect 37476 524106 37482 524108
rect 288934 524106 288940 524108
rect 37476 524046 288940 524106
rect 37476 524044 37482 524046
rect 288934 524044 288940 524046
rect 289004 524044 289010 524108
rect 291101 524106 291167 524109
rect 532049 524106 532115 524109
rect 291101 524104 532115 524106
rect 291101 524048 291106 524104
rect 291162 524048 532054 524104
rect 532110 524048 532115 524104
rect 291101 524046 532115 524048
rect 291101 524043 291167 524046
rect 532049 524043 532115 524046
rect 77661 523970 77727 523973
rect 280705 523970 280771 523973
rect 77661 523968 280771 523970
rect 77661 523912 77666 523968
rect 77722 523912 280710 523968
rect 280766 523912 280771 523968
rect 77661 523910 280771 523912
rect 77661 523907 77727 523910
rect 280705 523907 280771 523910
rect 283598 523908 283604 523972
rect 283668 523970 283674 523972
rect 536966 523970 536972 523972
rect 283668 523910 536972 523970
rect 283668 523908 283674 523910
rect 536966 523908 536972 523910
rect 537036 523908 537042 523972
rect 44582 523772 44588 523836
rect 44652 523834 44658 523836
rect 241329 523834 241395 523837
rect 44652 523832 241395 523834
rect 44652 523776 241334 523832
rect 241390 523776 241395 523832
rect 44652 523774 241395 523776
rect 44652 523772 44658 523774
rect 241329 523771 241395 523774
rect 38009 523698 38075 523701
rect 380985 523698 381051 523701
rect 38009 523696 381051 523698
rect 38009 523640 38014 523696
rect 38070 523640 380990 523696
rect 381046 523640 381051 523696
rect 38009 523638 381051 523640
rect 38009 523635 38075 523638
rect 380985 523635 381051 523638
rect 461577 523698 461643 523701
rect 523769 523698 523835 523701
rect 461577 523696 523835 523698
rect 461577 523640 461582 523696
rect 461638 523640 523774 523696
rect 523830 523640 523835 523696
rect 461577 523638 523835 523640
rect 461577 523635 461643 523638
rect 523769 523635 523835 523638
rect 46606 523500 46612 523564
rect 46676 523562 46682 523564
rect 288382 523562 288388 523564
rect 46676 523502 288388 523562
rect 46676 523500 46682 523502
rect 288382 523500 288388 523502
rect 288452 523500 288458 523564
rect 469857 523562 469923 523565
rect 519721 523562 519787 523565
rect 469857 523560 519787 523562
rect 469857 523504 469862 523560
rect 469918 523504 519726 523560
rect 519782 523504 519787 523560
rect 469857 523502 519787 523504
rect 469857 523499 469923 523502
rect 519721 523499 519787 523502
rect 32397 523426 32463 523429
rect 68921 523426 68987 523429
rect 32397 523424 68987 523426
rect 32397 523368 32402 523424
rect 32458 523368 68926 523424
rect 68982 523368 68987 523424
rect 32397 523366 68987 523368
rect 32397 523363 32463 523366
rect 68921 523363 68987 523366
rect 177798 523364 177804 523428
rect 177868 523426 177874 523428
rect 177941 523426 178007 523429
rect 177868 523424 178007 523426
rect 177868 523368 177946 523424
rect 178002 523368 178007 523424
rect 177868 523366 178007 523368
rect 177868 523364 177874 523366
rect 177941 523363 178007 523366
rect 299933 523426 299999 523429
rect 503253 523426 503319 523429
rect 299933 523424 503319 523426
rect 299933 523368 299938 523424
rect 299994 523368 503258 523424
rect 503314 523368 503319 523424
rect 299933 523366 503319 523368
rect 299933 523363 299999 523366
rect 503253 523363 503319 523366
rect 39246 523228 39252 523292
rect 39316 523290 39322 523292
rect 78581 523290 78647 523293
rect 39316 523288 78647 523290
rect 39316 523232 78586 523288
rect 78642 523232 78647 523288
rect 39316 523230 78647 523232
rect 39316 523228 39322 523230
rect 78581 523227 78647 523230
rect 240225 523290 240291 523293
rect 501505 523290 501571 523293
rect 240225 523288 501571 523290
rect 240225 523232 240230 523288
rect 240286 523232 501510 523288
rect 501566 523232 501571 523288
rect 240225 523230 501571 523232
rect 240225 523227 240291 523230
rect 501505 523227 501571 523230
rect 50153 523154 50219 523157
rect 53833 523154 53899 523157
rect 57697 523156 57763 523157
rect 57646 523154 57652 523156
rect 50153 523152 53899 523154
rect 50153 523096 50158 523152
rect 50214 523096 53838 523152
rect 53894 523096 53899 523152
rect 50153 523094 53899 523096
rect 57606 523094 57652 523154
rect 57716 523152 57763 523156
rect 313365 523154 313431 523157
rect 57758 523096 57763 523152
rect 50153 523091 50219 523094
rect 53833 523091 53899 523094
rect 57646 523092 57652 523094
rect 57716 523092 57763 523096
rect 57697 523091 57763 523092
rect 313046 523152 313431 523154
rect 313046 523096 313370 523152
rect 313426 523096 313431 523152
rect 313046 523094 313431 523096
rect 59997 523018 60063 523021
rect 224125 523018 224191 523021
rect 59997 523016 224191 523018
rect 59997 522960 60002 523016
rect 60058 522960 224130 523016
rect 224186 522960 224191 523016
rect 59997 522958 224191 522960
rect 59997 522955 60063 522958
rect 224125 522955 224191 522958
rect 226977 523018 227043 523021
rect 313046 523018 313106 523094
rect 313365 523091 313431 523094
rect 503713 523154 503779 523157
rect 503846 523154 503852 523156
rect 503713 523152 503852 523154
rect 503713 523096 503718 523152
rect 503774 523096 503852 523152
rect 503713 523094 503852 523096
rect 503713 523091 503779 523094
rect 503846 523092 503852 523094
rect 503916 523092 503922 523156
rect 517830 523092 517836 523156
rect 517900 523154 517906 523156
rect 518065 523154 518131 523157
rect 517900 523152 518131 523154
rect 517900 523096 518070 523152
rect 518126 523096 518131 523152
rect 517900 523094 518131 523096
rect 517900 523092 517906 523094
rect 518065 523091 518131 523094
rect 525793 523154 525859 523157
rect 525926 523154 525932 523156
rect 525793 523152 525932 523154
rect 525793 523096 525798 523152
rect 525854 523096 525932 523152
rect 525793 523094 525932 523096
rect 525793 523091 525859 523094
rect 525926 523092 525932 523094
rect 525996 523092 526002 523156
rect 226977 523016 313106 523018
rect 226977 522960 226982 523016
rect 227038 522960 313106 523016
rect 226977 522958 313106 522960
rect 313273 523018 313339 523021
rect 380893 523018 380959 523021
rect 313273 523016 380959 523018
rect 313273 522960 313278 523016
rect 313334 522960 380898 523016
rect 380954 522960 380959 523016
rect 313273 522958 380959 522960
rect 226977 522955 227043 522958
rect 313273 522955 313339 522958
rect 380893 522955 380959 522958
rect 483606 522956 483612 523020
rect 483676 523018 483682 523020
rect 519118 523018 519124 523020
rect 483676 522958 519124 523018
rect 483676 522956 483682 522958
rect 519118 522956 519124 522958
rect 519188 522956 519194 523020
rect 179045 522882 179111 522885
rect 257521 522882 257587 522885
rect 179045 522880 257587 522882
rect 179045 522824 179050 522880
rect 179106 522824 257526 522880
rect 257582 522824 257587 522880
rect 179045 522822 257587 522824
rect 179045 522819 179111 522822
rect 257521 522819 257587 522822
rect 264237 522882 264303 522885
rect 269665 522882 269731 522885
rect 264237 522880 269731 522882
rect 264237 522824 264242 522880
rect 264298 522824 269670 522880
rect 269726 522824 269731 522880
rect 264237 522822 269731 522824
rect 264237 522819 264303 522822
rect 269665 522819 269731 522822
rect 270217 522882 270283 522885
rect 271597 522882 271663 522885
rect 270217 522880 271663 522882
rect 270217 522824 270222 522880
rect 270278 522824 271602 522880
rect 271658 522824 271663 522880
rect 270217 522822 271663 522824
rect 270217 522819 270283 522822
rect 271597 522819 271663 522822
rect 271965 522882 272031 522885
rect 377949 522882 378015 522885
rect 271965 522880 378015 522882
rect 271965 522824 271970 522880
rect 272026 522824 377954 522880
rect 378010 522824 378015 522880
rect 271965 522822 378015 522824
rect 271965 522819 272031 522822
rect 377949 522819 378015 522822
rect 482134 522820 482140 522884
rect 482204 522882 482210 522884
rect 520222 522882 520228 522884
rect 482204 522822 520228 522882
rect 482204 522820 482210 522822
rect 520222 522820 520228 522822
rect 520292 522820 520298 522884
rect 37222 522684 37228 522748
rect 37292 522746 37298 522748
rect 253197 522746 253263 522749
rect 37292 522744 253263 522746
rect 37292 522688 253202 522744
rect 253258 522688 253263 522744
rect 37292 522686 253263 522688
rect 37292 522684 37298 522686
rect 253197 522683 253263 522686
rect 256693 522746 256759 522749
rect 376661 522746 376727 522749
rect 256693 522744 376727 522746
rect 256693 522688 256698 522744
rect 256754 522688 376666 522744
rect 376722 522688 376727 522744
rect 256693 522686 376727 522688
rect 256693 522683 256759 522686
rect 376661 522683 376727 522686
rect 478086 522684 478092 522748
rect 478156 522746 478162 522748
rect 520825 522746 520891 522749
rect 478156 522744 520891 522746
rect 478156 522688 520830 522744
rect 520886 522688 520891 522744
rect 478156 522686 520891 522688
rect 478156 522684 478162 522686
rect 520825 522683 520891 522686
rect 46105 522610 46171 522613
rect 178033 522610 178099 522613
rect 46105 522608 178099 522610
rect 46105 522552 46110 522608
rect 46166 522552 178038 522608
rect 178094 522552 178099 522608
rect 46105 522550 178099 522552
rect 46105 522547 46171 522550
rect 178033 522547 178099 522550
rect 228357 522610 228423 522613
rect 361849 522610 361915 522613
rect 228357 522608 361915 522610
rect 228357 522552 228362 522608
rect 228418 522552 361854 522608
rect 361910 522552 361915 522608
rect 228357 522550 361915 522552
rect 228357 522547 228423 522550
rect 361849 522547 361915 522550
rect 479374 522548 479380 522612
rect 479444 522610 479450 522612
rect 525190 522610 525196 522612
rect 479444 522550 525196 522610
rect 479444 522548 479450 522550
rect 525190 522548 525196 522550
rect 525260 522548 525266 522612
rect 184197 522474 184263 522477
rect 339493 522474 339559 522477
rect 184197 522472 339559 522474
rect 184197 522416 184202 522472
rect 184258 522416 339498 522472
rect 339554 522416 339559 522472
rect 184197 522414 339559 522416
rect 184197 522411 184263 522414
rect 339493 522411 339559 522414
rect 393957 522474 394023 522477
rect 420453 522474 420519 522477
rect 393957 522472 420519 522474
rect 393957 522416 393962 522472
rect 394018 522416 420458 522472
rect 420514 522416 420519 522472
rect 393957 522414 420519 522416
rect 393957 522411 394023 522414
rect 420453 522411 420519 522414
rect 475561 522474 475627 522477
rect 523585 522474 523651 522477
rect 475561 522472 523651 522474
rect 475561 522416 475566 522472
rect 475622 522416 523590 522472
rect 523646 522416 523651 522472
rect 475561 522414 523651 522416
rect 475561 522411 475627 522414
rect 523585 522411 523651 522414
rect 39614 522276 39620 522340
rect 39684 522338 39690 522340
rect 292614 522338 292620 522340
rect 39684 522278 292620 522338
rect 39684 522276 39690 522278
rect 292614 522276 292620 522278
rect 292684 522276 292690 522340
rect 295977 522338 296043 522341
rect 296897 522338 296963 522341
rect 295977 522336 296963 522338
rect 295977 522280 295982 522336
rect 296038 522280 296902 522336
rect 296958 522280 296963 522336
rect 295977 522278 296963 522280
rect 295977 522275 296043 522278
rect 296897 522275 296963 522278
rect 302233 522338 302299 522341
rect 304073 522338 304139 522341
rect 302233 522336 304139 522338
rect 302233 522280 302238 522336
rect 302294 522280 304078 522336
rect 304134 522280 304139 522336
rect 302233 522278 304139 522280
rect 302233 522275 302299 522278
rect 304073 522275 304139 522278
rect 314009 522338 314075 522341
rect 431677 522338 431743 522341
rect 314009 522336 431743 522338
rect 314009 522280 314014 522336
rect 314070 522280 431682 522336
rect 431738 522280 431743 522336
rect 314009 522278 431743 522280
rect 314009 522275 314075 522278
rect 431677 522275 431743 522278
rect 475745 522338 475811 522341
rect 524781 522338 524847 522341
rect 475745 522336 524847 522338
rect 475745 522280 475750 522336
rect 475806 522280 524786 522336
rect 524842 522280 524847 522336
rect 475745 522278 524847 522280
rect 475745 522275 475811 522278
rect 524781 522275 524847 522278
rect 224309 522202 224375 522205
rect 268745 522202 268811 522205
rect 224309 522200 268811 522202
rect 224309 522144 224314 522200
rect 224370 522144 268750 522200
rect 268806 522144 268811 522200
rect 224309 522142 268811 522144
rect 224309 522139 224375 522142
rect 268745 522139 268811 522142
rect 269021 522202 269087 522205
rect 271965 522202 272031 522205
rect 269021 522200 272031 522202
rect 269021 522144 269026 522200
rect 269082 522144 271970 522200
rect 272026 522144 272031 522200
rect 269021 522142 272031 522144
rect 269021 522139 269087 522142
rect 271965 522139 272031 522142
rect 296161 522202 296227 522205
rect 303061 522202 303127 522205
rect 296161 522200 303127 522202
rect 296161 522144 296166 522200
rect 296222 522144 303066 522200
rect 303122 522144 303127 522200
rect 296161 522142 303127 522144
rect 296161 522139 296227 522142
rect 303061 522139 303127 522142
rect 303613 522202 303679 522205
rect 378777 522202 378843 522205
rect 303613 522200 378843 522202
rect 303613 522144 303618 522200
rect 303674 522144 378782 522200
rect 378838 522144 378843 522200
rect 303613 522142 378843 522144
rect 303613 522139 303679 522142
rect 378777 522139 378843 522142
rect 490557 522202 490623 522205
rect 501965 522202 502031 522205
rect 490557 522200 502031 522202
rect 490557 522144 490562 522200
rect 490618 522144 501970 522200
rect 502026 522144 502031 522200
rect 490557 522142 502031 522144
rect 490557 522139 490623 522142
rect 501965 522139 502031 522142
rect 47577 522066 47643 522069
rect 226333 522066 226399 522069
rect 47577 522064 226399 522066
rect 47577 522008 47582 522064
rect 47638 522008 226338 522064
rect 226394 522008 226399 522064
rect 47577 522006 226399 522008
rect 47577 522003 47643 522006
rect 226333 522003 226399 522006
rect 253657 522066 253723 522069
rect 264605 522066 264671 522069
rect 253657 522064 264671 522066
rect 253657 522008 253662 522064
rect 253718 522008 264610 522064
rect 264666 522008 264671 522064
rect 253657 522006 264671 522008
rect 253657 522003 253723 522006
rect 264605 522003 264671 522006
rect 298001 522066 298067 522069
rect 314285 522066 314351 522069
rect 298001 522064 314351 522066
rect 298001 522008 298006 522064
rect 298062 522008 314290 522064
rect 314346 522008 314351 522064
rect 298001 522006 314351 522008
rect 298001 522003 298067 522006
rect 314285 522003 314351 522006
rect 43478 521868 43484 521932
rect 43548 521930 43554 521932
rect 43805 521930 43871 521933
rect 43548 521928 43871 521930
rect 43548 521872 43810 521928
rect 43866 521872 43871 521928
rect 43548 521870 43871 521872
rect 43548 521868 43554 521870
rect 43805 521867 43871 521870
rect 47853 521930 47919 521933
rect 227713 521930 227779 521933
rect 47853 521928 227779 521930
rect 47853 521872 47858 521928
rect 47914 521872 227718 521928
rect 227774 521872 227779 521928
rect 47853 521870 227779 521872
rect 47853 521867 47919 521870
rect 227713 521867 227779 521870
rect 500033 521930 500099 521933
rect 500718 521930 500724 521932
rect 500033 521928 500724 521930
rect 500033 521872 500038 521928
rect 500094 521872 500724 521928
rect 500033 521870 500724 521872
rect 500033 521867 500099 521870
rect 500718 521868 500724 521870
rect 500788 521868 500794 521932
rect 43662 521732 43668 521796
rect 43732 521794 43738 521796
rect 44081 521794 44147 521797
rect 43732 521792 44147 521794
rect 43732 521736 44086 521792
rect 44142 521736 44147 521792
rect 43732 521734 44147 521736
rect 43732 521732 43738 521734
rect 44081 521731 44147 521734
rect 48865 521794 48931 521797
rect 184841 521794 184907 521797
rect 48865 521792 184907 521794
rect 48865 521736 48870 521792
rect 48926 521736 184846 521792
rect 184902 521736 184907 521792
rect 48865 521734 184907 521736
rect 48865 521731 48931 521734
rect 184841 521731 184907 521734
rect 499246 521732 499252 521796
rect 499316 521794 499322 521796
rect 500861 521794 500927 521797
rect 499316 521792 500927 521794
rect 499316 521736 500866 521792
rect 500922 521736 500927 521792
rect 499316 521734 500927 521736
rect 499316 521732 499322 521734
rect 500861 521731 500927 521734
rect 517513 521794 517579 521797
rect 518198 521794 518204 521796
rect 517513 521792 518204 521794
rect 517513 521736 517518 521792
rect 517574 521736 518204 521792
rect 517513 521734 518204 521736
rect 517513 521731 517579 521734
rect 518198 521732 518204 521734
rect 518268 521732 518274 521796
rect 167637 521658 167703 521661
rect 301129 521658 301195 521661
rect 167637 521656 301195 521658
rect 167637 521600 167642 521656
rect 167698 521600 301134 521656
rect 301190 521600 301195 521656
rect 167637 521598 301195 521600
rect 167637 521595 167703 521598
rect 301129 521595 301195 521598
rect 468569 521658 468635 521661
rect 498101 521658 498167 521661
rect 468569 521656 498167 521658
rect 468569 521600 468574 521656
rect 468630 521600 498106 521656
rect 498162 521600 498167 521656
rect 468569 521598 498167 521600
rect 468569 521595 468635 521598
rect 498101 521595 498167 521598
rect 498694 521596 498700 521660
rect 498764 521658 498770 521660
rect 500534 521658 500540 521660
rect 498764 521598 500540 521658
rect 498764 521596 498770 521598
rect 500534 521596 500540 521598
rect 500604 521596 500610 521660
rect 530526 521596 530532 521660
rect 530596 521658 530602 521660
rect 531221 521658 531287 521661
rect 530596 521656 531287 521658
rect 530596 521600 531226 521656
rect 531282 521600 531287 521656
rect 530596 521598 531287 521600
rect 530596 521596 530602 521598
rect 531221 521595 531287 521598
rect 166441 521522 166507 521525
rect 300025 521522 300091 521525
rect 166441 521520 300091 521522
rect 166441 521464 166446 521520
rect 166502 521464 300030 521520
rect 300086 521464 300091 521520
rect 166441 521462 300091 521464
rect 166441 521459 166507 521462
rect 300025 521459 300091 521462
rect 461669 521522 461735 521525
rect 518341 521522 518407 521525
rect 461669 521520 518407 521522
rect 461669 521464 461674 521520
rect 461730 521464 518346 521520
rect 518402 521464 518407 521520
rect 461669 521462 518407 521464
rect 461669 521459 461735 521462
rect 518341 521459 518407 521462
rect 167821 521386 167887 521389
rect 299013 521386 299079 521389
rect 167821 521384 299079 521386
rect 167821 521328 167826 521384
rect 167882 521328 299018 521384
rect 299074 521328 299079 521384
rect 167821 521326 299079 521328
rect 167821 521323 167887 521326
rect 299013 521323 299079 521326
rect 299790 521324 299796 521388
rect 299860 521386 299866 521388
rect 503110 521386 503116 521388
rect 299860 521326 503116 521386
rect 299860 521324 299866 521326
rect 503110 521324 503116 521326
rect 503180 521324 503186 521388
rect 39297 521250 39363 521253
rect 222101 521250 222167 521253
rect 39297 521248 222167 521250
rect 39297 521192 39302 521248
rect 39358 521192 222106 521248
rect 222162 521192 222167 521248
rect 39297 521190 222167 521192
rect 39297 521187 39363 521190
rect 222101 521187 222167 521190
rect 287830 521188 287836 521252
rect 287900 521250 287906 521252
rect 505318 521250 505324 521252
rect 287900 521190 505324 521250
rect 287900 521188 287906 521190
rect 505318 521188 505324 521190
rect 505388 521188 505394 521252
rect 517053 521250 517119 521253
rect 527214 521250 527220 521252
rect 517053 521248 527220 521250
rect 517053 521192 517058 521248
rect 517114 521192 527220 521248
rect 517053 521190 527220 521192
rect 517053 521187 517119 521190
rect 527214 521188 527220 521190
rect 527284 521188 527290 521252
rect 47485 521114 47551 521117
rect 166993 521114 167059 521117
rect 47485 521112 167059 521114
rect 47485 521056 47490 521112
rect 47546 521056 166998 521112
rect 167054 521056 167059 521112
rect 47485 521054 167059 521056
rect 47485 521051 47551 521054
rect 166993 521051 167059 521054
rect 220997 521114 221063 521117
rect 291837 521114 291903 521117
rect 220997 521112 291903 521114
rect 220997 521056 221002 521112
rect 221058 521056 291842 521112
rect 291898 521056 291903 521112
rect 220997 521054 291903 521056
rect 220997 521051 221063 521054
rect 291837 521051 291903 521054
rect 500125 521114 500191 521117
rect 508078 521114 508084 521116
rect 500125 521112 508084 521114
rect 500125 521056 500130 521112
rect 500186 521056 508084 521112
rect 500125 521054 508084 521056
rect 500125 521051 500191 521054
rect 508078 521052 508084 521054
rect 508148 521052 508154 521116
rect 57830 520916 57836 520980
rect 57900 520978 57906 520980
rect 254526 520978 254532 520980
rect 57900 520918 254532 520978
rect 57900 520916 57906 520918
rect 254526 520916 254532 520918
rect 254596 520916 254602 520980
rect 283414 520916 283420 520980
rect 283484 520978 283490 520980
rect 531446 520978 531452 520980
rect 283484 520918 531452 520978
rect 283484 520916 283490 520918
rect 531446 520916 531452 520918
rect 531516 520916 531522 520980
rect 46197 520842 46263 520845
rect 167085 520842 167151 520845
rect 46197 520840 167151 520842
rect 46197 520784 46202 520840
rect 46258 520784 167090 520840
rect 167146 520784 167151 520840
rect 46197 520782 167151 520784
rect 46197 520779 46263 520782
rect 167085 520779 167151 520782
rect 169017 520842 169083 520845
rect 302049 520842 302115 520845
rect 169017 520840 302115 520842
rect 169017 520784 169022 520840
rect 169078 520784 302054 520840
rect 302110 520784 302115 520840
rect 169017 520782 302115 520784
rect 169017 520779 169083 520782
rect 302049 520779 302115 520782
rect 497590 520780 497596 520844
rect 497660 520842 497666 520844
rect 508446 520842 508452 520844
rect 497660 520782 508452 520842
rect 497660 520780 497666 520782
rect 508446 520780 508452 520782
rect 508516 520780 508522 520844
rect 41965 520706 42031 520709
rect 166257 520706 166323 520709
rect 41965 520704 166323 520706
rect 41965 520648 41970 520704
rect 42026 520648 166262 520704
rect 166318 520648 166323 520704
rect 41965 520646 166323 520648
rect 41965 520643 42031 520646
rect 166257 520643 166323 520646
rect 219985 520706 220051 520709
rect 288341 520706 288407 520709
rect 219985 520704 288407 520706
rect 219985 520648 219990 520704
rect 220046 520648 288346 520704
rect 288402 520648 288407 520704
rect 219985 520646 288407 520648
rect 219985 520643 220051 520646
rect 288341 520643 288407 520646
rect 499430 520644 499436 520708
rect 499500 520706 499506 520708
rect 500350 520706 500356 520708
rect 499500 520646 500356 520706
rect 499500 520644 499506 520646
rect 500350 520644 500356 520646
rect 500420 520644 500426 520708
rect 40902 520508 40908 520572
rect 40972 520570 40978 520572
rect 168373 520570 168439 520573
rect 40972 520568 168439 520570
rect 40972 520512 168378 520568
rect 168434 520512 168439 520568
rect 40972 520510 168439 520512
rect 40972 520508 40978 520510
rect 168373 520507 168439 520510
rect 489545 520570 489611 520573
rect 498101 520570 498167 520573
rect 489545 520568 498167 520570
rect 489545 520512 489550 520568
rect 489606 520512 498106 520568
rect 498162 520512 498167 520568
rect 489545 520510 498167 520512
rect 489545 520507 489611 520510
rect 498101 520507 498167 520510
rect 499430 520508 499436 520572
rect 499500 520570 499506 520572
rect 500309 520570 500375 520573
rect 499500 520568 500375 520570
rect 499500 520512 500314 520568
rect 500370 520512 500375 520568
rect 499500 520510 500375 520512
rect 499500 520508 499506 520510
rect 500309 520507 500375 520510
rect 504633 520570 504699 520573
rect 511625 520570 511691 520573
rect 504633 520568 511691 520570
rect 504633 520512 504638 520568
rect 504694 520512 511630 520568
rect 511686 520512 511691 520568
rect 504633 520510 511691 520512
rect 504633 520507 504699 520510
rect 511625 520507 511691 520510
rect 46473 520434 46539 520437
rect 220721 520434 220787 520437
rect 46473 520432 220787 520434
rect 46473 520376 46478 520432
rect 46534 520376 220726 520432
rect 220782 520376 220787 520432
rect 46473 520374 220787 520376
rect 46473 520371 46539 520374
rect 220721 520371 220787 520374
rect 291878 520372 291884 520436
rect 291948 520434 291954 520436
rect 538438 520434 538444 520436
rect 291948 520374 538444 520434
rect 291948 520372 291954 520374
rect 538438 520372 538444 520374
rect 538508 520372 538514 520436
rect 50286 520236 50292 520300
rect 50356 520298 50362 520300
rect 50981 520298 51047 520301
rect 50356 520296 51047 520298
rect 50356 520240 50986 520296
rect 51042 520240 51047 520296
rect 50356 520238 51047 520240
rect 50356 520236 50362 520238
rect 50981 520235 51047 520238
rect 51206 520236 51212 520300
rect 51276 520298 51282 520300
rect 51533 520298 51599 520301
rect 51276 520296 51599 520298
rect 51276 520240 51538 520296
rect 51594 520240 51599 520296
rect 51276 520238 51599 520240
rect 51276 520236 51282 520238
rect 51533 520235 51599 520238
rect 52126 520236 52132 520300
rect 52196 520298 52202 520300
rect 52361 520298 52427 520301
rect 61837 520300 61903 520301
rect 52196 520296 52427 520298
rect 52196 520240 52366 520296
rect 52422 520240 52427 520296
rect 52196 520238 52427 520240
rect 52196 520236 52202 520238
rect 52361 520235 52427 520238
rect 59670 520236 59676 520300
rect 59740 520298 59746 520300
rect 61326 520298 61332 520300
rect 59740 520238 61332 520298
rect 59740 520236 59746 520238
rect 61326 520236 61332 520238
rect 61396 520236 61402 520300
rect 61837 520298 61884 520300
rect 61792 520296 61884 520298
rect 61792 520240 61842 520296
rect 61792 520238 61884 520240
rect 61837 520236 61884 520238
rect 61948 520236 61954 520300
rect 497406 520236 497412 520300
rect 497476 520298 497482 520300
rect 499982 520298 499988 520300
rect 497476 520238 499988 520298
rect 497476 520236 497482 520238
rect 499982 520236 499988 520238
rect 500052 520236 500058 520300
rect 502241 520298 502307 520301
rect 500174 520296 502307 520298
rect 500174 520240 502246 520296
rect 502302 520240 502307 520296
rect 500174 520238 502307 520240
rect 61837 520235 61903 520236
rect 55029 520162 55095 520165
rect 62113 520162 62179 520165
rect 55029 520160 62179 520162
rect 55029 520104 55034 520160
rect 55090 520104 62118 520160
rect 62174 520104 62179 520160
rect 55029 520102 62179 520104
rect 55029 520099 55095 520102
rect 62113 520099 62179 520102
rect 497365 520162 497431 520165
rect 499430 520162 499436 520164
rect 497365 520160 499436 520162
rect 497365 520104 497370 520160
rect 497426 520104 499436 520160
rect 497365 520102 499436 520104
rect 497365 520099 497431 520102
rect 499430 520100 499436 520102
rect 499500 520100 499506 520164
rect 499573 520162 499639 520165
rect 500174 520162 500234 520238
rect 502241 520235 502307 520238
rect 502926 520236 502932 520300
rect 502996 520298 503002 520300
rect 503161 520298 503227 520301
rect 502996 520296 503227 520298
rect 502996 520240 503166 520296
rect 503222 520240 503227 520296
rect 502996 520238 503227 520240
rect 502996 520236 503002 520238
rect 503161 520235 503227 520238
rect 514753 520298 514819 520301
rect 515070 520298 515076 520300
rect 514753 520296 515076 520298
rect 514753 520240 514758 520296
rect 514814 520240 515076 520296
rect 514753 520238 515076 520240
rect 514753 520235 514819 520238
rect 515070 520236 515076 520238
rect 515140 520236 515146 520300
rect 499573 520160 500234 520162
rect 499573 520104 499578 520160
rect 499634 520104 500234 520160
rect 499573 520102 500234 520104
rect 500309 520162 500375 520165
rect 500309 520160 505110 520162
rect 500309 520104 500314 520160
rect 500370 520104 505110 520160
rect 500309 520102 505110 520104
rect 499573 520099 499639 520102
rect 500309 520099 500375 520102
rect 55438 519964 55444 520028
rect 55508 520026 55514 520028
rect 59721 520026 59787 520029
rect 55508 520024 59787 520026
rect 55508 519968 59726 520024
rect 59782 519968 59787 520024
rect 55508 519966 59787 519968
rect 55508 519964 55514 519966
rect 59721 519963 59787 519966
rect 500401 520026 500467 520029
rect 501086 520026 501092 520028
rect 500401 520024 501092 520026
rect 500401 519968 500406 520024
rect 500462 519968 501092 520024
rect 500401 519966 501092 519968
rect 500401 519963 500467 519966
rect 501086 519964 501092 519966
rect 501156 519964 501162 520028
rect 505050 520026 505110 520102
rect 529238 520026 529244 520028
rect 505050 519966 529244 520026
rect 529238 519964 529244 519966
rect 529308 519964 529314 520028
rect 59813 519890 59879 519893
rect 60641 519890 60707 519893
rect 59813 519888 60707 519890
rect 59813 519832 59818 519888
rect 59874 519832 60646 519888
rect 60702 519832 60707 519888
rect 59813 519830 60707 519832
rect 59813 519827 59879 519830
rect 60641 519827 60707 519830
rect 500861 519890 500927 519893
rect 514109 519890 514175 519893
rect 500861 519888 514175 519890
rect 500861 519832 500866 519888
rect 500922 519832 514114 519888
rect 514170 519832 514175 519888
rect 500861 519830 514175 519832
rect 500861 519827 500927 519830
rect 514109 519827 514175 519830
rect 500534 519692 500540 519756
rect 500604 519754 500610 519756
rect 506013 519754 506079 519757
rect 507158 519754 507164 519756
rect 500604 519694 505110 519754
rect 500604 519692 500610 519694
rect 50654 519556 50660 519620
rect 50724 519618 50730 519620
rect 60641 519618 60707 519621
rect 50724 519616 60707 519618
rect 50724 519560 60646 519616
rect 60702 519560 60707 519616
rect 50724 519558 60707 519560
rect 50724 519556 50730 519558
rect 60641 519555 60707 519558
rect 499573 519618 499639 519621
rect 500718 519618 500724 519620
rect 499573 519616 500724 519618
rect 499573 519560 499578 519616
rect 499634 519560 500724 519616
rect 499573 519558 500724 519560
rect 499573 519555 499639 519558
rect 500718 519556 500724 519558
rect 500788 519556 500794 519620
rect 503713 519618 503779 519621
rect 504030 519618 504036 519620
rect 503713 519616 504036 519618
rect 503713 519560 503718 519616
rect 503774 519560 504036 519616
rect 503713 519558 504036 519560
rect 503713 519555 503779 519558
rect 504030 519556 504036 519558
rect 504100 519556 504106 519620
rect 505050 519618 505110 519694
rect 506013 519752 507164 519754
rect 506013 519696 506018 519752
rect 506074 519696 507164 519752
rect 506013 519694 507164 519696
rect 506013 519691 506079 519694
rect 507158 519692 507164 519694
rect 507228 519692 507234 519756
rect 507945 519754 508011 519757
rect 510705 519754 510771 519757
rect 507945 519752 510771 519754
rect 507945 519696 507950 519752
rect 508006 519696 510710 519752
rect 510766 519696 510771 519752
rect 507945 519694 510771 519696
rect 507945 519691 508011 519694
rect 510705 519691 510771 519694
rect 511533 519754 511599 519757
rect 526294 519754 526300 519756
rect 511533 519752 526300 519754
rect 511533 519696 511538 519752
rect 511594 519696 526300 519752
rect 511533 519694 526300 519696
rect 511533 519691 511599 519694
rect 526294 519692 526300 519694
rect 526364 519692 526370 519756
rect 516358 519618 516364 519620
rect 505050 519558 516364 519618
rect 516358 519556 516364 519558
rect 516428 519556 516434 519620
rect 46013 519482 46079 519485
rect 59261 519482 59327 519485
rect 46013 519480 59327 519482
rect 46013 519424 46018 519480
rect 46074 519424 59266 519480
rect 59322 519424 59327 519480
rect 46013 519422 59327 519424
rect 46013 519419 46079 519422
rect 59261 519419 59327 519422
rect 500350 519420 500356 519484
rect 500420 519482 500426 519484
rect 522246 519482 522252 519484
rect 500420 519422 522252 519482
rect 500420 519420 500426 519422
rect 522246 519420 522252 519422
rect 522316 519420 522322 519484
rect 51574 519284 51580 519348
rect 51644 519346 51650 519348
rect 52361 519346 52427 519349
rect 60641 519346 60707 519349
rect 51644 519344 52427 519346
rect 51644 519288 52366 519344
rect 52422 519288 52427 519344
rect 51644 519286 52427 519288
rect 51644 519284 51650 519286
rect 52361 519283 52427 519286
rect 55170 519344 60707 519346
rect 55170 519288 60646 519344
rect 60702 519288 60707 519344
rect 55170 519286 60707 519288
rect 47393 519210 47459 519213
rect 55170 519210 55230 519286
rect 60641 519283 60707 519286
rect 500861 519346 500927 519349
rect 510613 519346 510679 519349
rect 511206 519346 511212 519348
rect 500861 519344 510354 519346
rect 500861 519288 500866 519344
rect 500922 519288 510354 519344
rect 500861 519286 510354 519288
rect 500861 519283 500927 519286
rect 47393 519208 55230 519210
rect 47393 519152 47398 519208
rect 47454 519152 55230 519208
rect 47393 519150 55230 519152
rect 501873 519210 501939 519213
rect 509417 519210 509483 519213
rect 501873 519208 509483 519210
rect 501873 519152 501878 519208
rect 501934 519152 509422 519208
rect 509478 519152 509483 519208
rect 501873 519150 509483 519152
rect 47393 519147 47459 519150
rect 501873 519147 501939 519150
rect 509417 519147 509483 519150
rect 502149 519074 502215 519077
rect 507945 519074 508011 519077
rect 502149 519072 508011 519074
rect 502149 519016 502154 519072
rect 502210 519016 507950 519072
rect 508006 519016 508011 519072
rect 502149 519014 508011 519016
rect 510294 519074 510354 519286
rect 510613 519344 511212 519346
rect 510613 519288 510618 519344
rect 510674 519288 511212 519344
rect 510613 519286 511212 519288
rect 510613 519283 510679 519286
rect 511206 519284 511212 519286
rect 511276 519284 511282 519348
rect 512637 519074 512703 519077
rect 510294 519072 512703 519074
rect 510294 519016 512642 519072
rect 512698 519016 512703 519072
rect 510294 519014 512703 519016
rect 502149 519011 502215 519014
rect 507945 519011 508011 519014
rect 512637 519011 512703 519014
rect 44030 518740 44036 518804
rect 44100 518802 44106 518804
rect 44100 518742 60076 518802
rect 44100 518740 44106 518742
rect 59813 518258 59879 518261
rect 59813 518256 60076 518258
rect 59813 518200 59818 518256
rect 59874 518200 60076 518256
rect 59813 518198 60076 518200
rect 59813 518195 59879 518198
rect 60089 517986 60155 517989
rect 60046 517984 60155 517986
rect 60046 517928 60094 517984
rect 60150 517928 60155 517984
rect 60046 517923 60155 517928
rect 60046 517684 60106 517923
rect 57329 517170 57395 517173
rect 57329 517168 60076 517170
rect 57329 517112 57334 517168
rect 57390 517112 60076 517168
rect 57329 517110 60076 517112
rect 57329 517107 57395 517110
rect 46565 516626 46631 516629
rect 46565 516624 60076 516626
rect 46565 516568 46570 516624
rect 46626 516568 60076 516624
rect 46565 516566 60076 516568
rect 46565 516563 46631 516566
rect 57605 516082 57671 516085
rect 57605 516080 60076 516082
rect 57605 516024 57610 516080
rect 57666 516024 60076 516080
rect 57605 516022 60076 516024
rect 57605 516019 57671 516022
rect 57421 515538 57487 515541
rect 57421 515536 60076 515538
rect 57421 515480 57426 515536
rect 57482 515480 60076 515536
rect 57421 515478 60076 515480
rect 57421 515475 57487 515478
rect 31150 514994 31156 514996
rect -960 514858 480 514948
rect 26190 514934 31156 514994
rect 26190 514858 26250 514934
rect 31150 514932 31156 514934
rect 31220 514932 31226 514996
rect 57789 514994 57855 514997
rect 57789 514992 60076 514994
rect 57789 514936 57794 514992
rect 57850 514936 60076 514992
rect 57789 514934 60076 514936
rect 57789 514931 57855 514934
rect -960 514798 26250 514858
rect -960 514708 480 514798
rect 30414 514796 30420 514860
rect 30484 514858 30490 514860
rect 31385 514858 31451 514861
rect 30484 514856 31451 514858
rect 30484 514800 31390 514856
rect 31446 514800 31451 514856
rect 30484 514798 31451 514800
rect 30484 514796 30490 514798
rect 31385 514795 31451 514798
rect 514661 514724 514727 514725
rect 514661 514722 514708 514724
rect 514616 514720 514708 514722
rect 514616 514664 514666 514720
rect 514616 514662 514708 514664
rect 514661 514660 514708 514662
rect 514772 514660 514778 514724
rect 514661 514659 514727 514660
rect 55990 514388 55996 514452
rect 56060 514450 56066 514452
rect 56060 514390 60076 514450
rect 56060 514388 56066 514390
rect 55622 513980 55628 514044
rect 55692 514042 55698 514044
rect 56501 514042 56567 514045
rect 55692 514040 56567 514042
rect 55692 513984 56506 514040
rect 56562 513984 56567 514040
rect 55692 513982 56567 513984
rect 55692 513980 55698 513982
rect 56501 513979 56567 513982
rect 57881 513906 57947 513909
rect 57881 513904 60076 513906
rect 57881 513848 57886 513904
rect 57942 513848 60076 513904
rect 57881 513846 60076 513848
rect 57881 513843 57947 513846
rect 509969 513498 510035 513501
rect 510838 513498 510844 513500
rect 509969 513496 510844 513498
rect 509969 513440 509974 513496
rect 510030 513440 510844 513496
rect 509969 513438 510844 513440
rect 509969 513435 510035 513438
rect 510838 513436 510844 513438
rect 510908 513436 510914 513500
rect 53782 513300 53788 513364
rect 53852 513362 53858 513364
rect 54569 513362 54635 513365
rect 53852 513360 54635 513362
rect 53852 513304 54574 513360
rect 54630 513304 54635 513360
rect 53852 513302 54635 513304
rect 53852 513300 53858 513302
rect 54569 513299 54635 513302
rect 57237 513362 57303 513365
rect 57237 513360 60076 513362
rect 57237 513304 57242 513360
rect 57298 513304 60076 513360
rect 57237 513302 60076 513304
rect 57237 513299 57303 513302
rect 57053 512818 57119 512821
rect 57053 512816 60076 512818
rect 57053 512760 57058 512816
rect 57114 512760 60076 512816
rect 57053 512758 60076 512760
rect 57053 512755 57119 512758
rect 57513 512274 57579 512277
rect 57513 512272 60076 512274
rect 57513 512216 57518 512272
rect 57574 512216 60076 512272
rect 57513 512214 60076 512216
rect 57513 512211 57579 512214
rect 502241 512002 502307 512005
rect 504030 512002 504036 512004
rect 502241 512000 504036 512002
rect 502241 511944 502246 512000
rect 502302 511944 504036 512000
rect 502241 511942 504036 511944
rect 502241 511939 502307 511942
rect 504030 511940 504036 511942
rect 504100 511940 504106 512004
rect 500585 511866 500651 511869
rect 504030 511866 504036 511868
rect 500585 511864 504036 511866
rect 500585 511808 500590 511864
rect 500646 511808 504036 511864
rect 500585 511806 504036 511808
rect 500585 511803 500651 511806
rect 504030 511804 504036 511806
rect 504100 511804 504106 511868
rect 56961 511730 57027 511733
rect 56961 511728 60076 511730
rect 56961 511672 56966 511728
rect 57022 511672 60076 511728
rect 56961 511670 60076 511672
rect 56961 511667 57027 511670
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 57145 511186 57211 511189
rect 57145 511184 60076 511186
rect 57145 511128 57150 511184
rect 57206 511128 60076 511184
rect 583520 511172 584960 511262
rect 57145 511126 60076 511128
rect 57145 511123 57211 511126
rect 50654 510580 50660 510644
rect 50724 510642 50730 510644
rect 57513 510642 57579 510645
rect 50724 510640 57579 510642
rect 50724 510584 57518 510640
rect 57574 510584 57579 510640
rect 50724 510582 57579 510584
rect 50724 510580 50730 510582
rect 57513 510579 57579 510582
rect 57646 510580 57652 510644
rect 57716 510642 57722 510644
rect 57716 510582 60076 510642
rect 57716 510580 57722 510582
rect 44633 510098 44699 510101
rect 44633 510096 60076 510098
rect 44633 510040 44638 510096
rect 44694 510040 60076 510096
rect 44633 510038 60076 510040
rect 44633 510035 44699 510038
rect 43846 509492 43852 509556
rect 43916 509554 43922 509556
rect 43916 509494 60076 509554
rect 43916 509492 43922 509494
rect 41873 509010 41939 509013
rect 41873 509008 60076 509010
rect 41873 508952 41878 509008
rect 41934 508952 60076 509008
rect 41873 508950 60076 508952
rect 41873 508947 41939 508950
rect 47393 508602 47459 508605
rect 57646 508602 57652 508604
rect 47393 508600 57652 508602
rect 47393 508544 47398 508600
rect 47454 508544 57652 508600
rect 47393 508542 57652 508544
rect 47393 508539 47459 508542
rect 57646 508540 57652 508542
rect 57716 508540 57722 508604
rect 46105 508466 46171 508469
rect 46105 508464 60076 508466
rect 46105 508408 46110 508464
rect 46166 508408 60076 508464
rect 46105 508406 60076 508408
rect 46105 508403 46171 508406
rect 39205 507922 39271 507925
rect 39205 507920 60076 507922
rect 39205 507864 39210 507920
rect 39266 507864 60076 507920
rect 39205 507862 60076 507864
rect 39205 507859 39271 507862
rect 41270 507316 41276 507380
rect 41340 507378 41346 507380
rect 41340 507318 60076 507378
rect 41340 507316 41346 507318
rect 48865 506834 48931 506837
rect 48865 506832 60076 506834
rect 48865 506776 48870 506832
rect 48926 506776 60076 506832
rect 48865 506774 60076 506776
rect 48865 506771 48931 506774
rect 40769 506562 40835 506565
rect 41270 506562 41276 506564
rect 40769 506560 41276 506562
rect 40769 506504 40774 506560
rect 40830 506504 41276 506560
rect 40769 506502 41276 506504
rect 40769 506499 40835 506502
rect 41270 506500 41276 506502
rect 41340 506500 41346 506564
rect 47393 506562 47459 506565
rect 49734 506562 49740 506564
rect 47393 506560 49740 506562
rect 47393 506504 47398 506560
rect 47454 506504 49740 506560
rect 47393 506502 49740 506504
rect 47393 506499 47459 506502
rect 49734 506500 49740 506502
rect 49804 506500 49810 506564
rect 38101 506290 38167 506293
rect 38101 506288 60076 506290
rect 38101 506232 38106 506288
rect 38162 506232 60076 506288
rect 38101 506230 60076 506232
rect 38101 506227 38167 506230
rect 47853 505882 47919 505885
rect 57605 505882 57671 505885
rect 47853 505880 57671 505882
rect 47853 505824 47858 505880
rect 47914 505824 57610 505880
rect 57666 505824 57671 505880
rect 47853 505822 57671 505824
rect 47853 505819 47919 505822
rect 57605 505819 57671 505822
rect 57646 505684 57652 505748
rect 57716 505746 57722 505748
rect 57716 505686 60076 505746
rect 57716 505684 57722 505686
rect 57462 505276 57468 505340
rect 57532 505338 57538 505340
rect 60181 505338 60247 505341
rect 514661 505340 514727 505341
rect 514661 505338 514708 505340
rect 57532 505336 60247 505338
rect 57532 505280 60186 505336
rect 60242 505280 60247 505336
rect 57532 505278 60247 505280
rect 514616 505336 514708 505338
rect 514616 505280 514666 505336
rect 514616 505278 514708 505280
rect 57532 505276 57538 505278
rect 60181 505275 60247 505278
rect 514661 505276 514708 505278
rect 514772 505276 514778 505340
rect 514661 505275 514727 505276
rect 35566 505140 35572 505204
rect 35636 505202 35642 505204
rect 35636 505142 60076 505202
rect 35636 505140 35642 505142
rect 33869 504658 33935 504661
rect 33869 504656 60076 504658
rect 33869 504600 33874 504656
rect 33930 504600 60076 504656
rect 33869 504598 60076 504600
rect 33869 504595 33935 504598
rect 37917 504114 37983 504117
rect 37917 504112 60076 504114
rect 37917 504056 37922 504112
rect 37978 504056 60076 504112
rect 37917 504054 60076 504056
rect 37917 504051 37983 504054
rect 31109 503706 31175 503709
rect 37917 503706 37983 503709
rect 31109 503704 37983 503706
rect 31109 503648 31114 503704
rect 31170 503648 37922 503704
rect 37978 503648 37983 503704
rect 31109 503646 37983 503648
rect 31109 503643 31175 503646
rect 37917 503643 37983 503646
rect 51022 503644 51028 503708
rect 51092 503706 51098 503708
rect 53097 503706 53163 503709
rect 51092 503704 53163 503706
rect 51092 503648 53102 503704
rect 53158 503648 53163 503704
rect 51092 503646 53163 503648
rect 51092 503644 51098 503646
rect 53097 503643 53163 503646
rect 55438 503644 55444 503708
rect 55508 503706 55514 503708
rect 57421 503706 57487 503709
rect 55508 503704 57487 503706
rect 55508 503648 57426 503704
rect 57482 503648 57487 503704
rect 55508 503646 57487 503648
rect 55508 503644 55514 503646
rect 57421 503643 57487 503646
rect 54518 503508 54524 503572
rect 54588 503570 54594 503572
rect 54588 503510 60076 503570
rect 54588 503508 54594 503510
rect 58566 502964 58572 503028
rect 58636 503026 58642 503028
rect 58636 502966 60076 503026
rect 58636 502964 58642 502966
rect 40718 502420 40724 502484
rect 40788 502482 40794 502484
rect 40788 502422 60076 502482
rect 40788 502420 40794 502422
rect 38878 502284 38884 502348
rect 38948 502346 38954 502348
rect 39665 502346 39731 502349
rect 38948 502344 39731 502346
rect 38948 502288 39670 502344
rect 39726 502288 39731 502344
rect 38948 502286 39731 502288
rect 38948 502284 38954 502286
rect 39665 502283 39731 502286
rect -960 501802 480 501892
rect 36670 501876 36676 501940
rect 36740 501938 36746 501940
rect 36740 501878 60076 501938
rect 36740 501876 36746 501878
rect 22686 501802 22692 501804
rect -960 501742 22692 501802
rect -960 501652 480 501742
rect 22686 501740 22692 501742
rect 22756 501740 22762 501804
rect 39798 501332 39804 501396
rect 39868 501394 39874 501396
rect 39868 501334 60076 501394
rect 39868 501332 39874 501334
rect 44725 500850 44791 500853
rect 44725 500848 60076 500850
rect 44725 500792 44730 500848
rect 44786 500792 60076 500848
rect 44725 500790 60076 500792
rect 44725 500787 44791 500790
rect 55622 500652 55628 500716
rect 55692 500714 55698 500716
rect 57329 500714 57395 500717
rect 55692 500712 57395 500714
rect 55692 500656 57334 500712
rect 57390 500656 57395 500712
rect 55692 500654 57395 500656
rect 55692 500652 55698 500654
rect 57329 500651 57395 500654
rect 59997 500578 60063 500581
rect 59997 500576 60106 500578
rect 59997 500520 60002 500576
rect 60058 500520 60106 500576
rect 59997 500515 60106 500520
rect 60046 500276 60106 500515
rect 52126 499836 52132 499900
rect 52196 499898 52202 499900
rect 55857 499898 55923 499901
rect 52196 499896 55923 499898
rect 52196 499840 55862 499896
rect 55918 499840 55923 499896
rect 52196 499838 55923 499840
rect 52196 499836 52202 499838
rect 55857 499835 55923 499838
rect 47485 499762 47551 499765
rect 47485 499760 60076 499762
rect 47485 499704 47490 499760
rect 47546 499704 60076 499760
rect 47485 499702 60076 499704
rect 47485 499699 47551 499702
rect 57462 499156 57468 499220
rect 57532 499218 57538 499220
rect 57532 499158 60076 499218
rect 57532 499156 57538 499158
rect 46197 498946 46263 498949
rect 57646 498946 57652 498948
rect 46197 498944 57652 498946
rect 46197 498888 46202 498944
rect 46258 498888 57652 498944
rect 46197 498886 57652 498888
rect 46197 498883 46263 498886
rect 57646 498884 57652 498886
rect 57716 498884 57722 498948
rect 43253 498810 43319 498813
rect 57513 498810 57579 498813
rect 43253 498808 57579 498810
rect 43253 498752 43258 498808
rect 43314 498752 57518 498808
rect 57574 498752 57579 498808
rect 43253 498750 57579 498752
rect 43253 498747 43319 498750
rect 57513 498747 57579 498750
rect 32397 498674 32463 498677
rect 32397 498672 60076 498674
rect 32397 498616 32402 498672
rect 32458 498616 60076 498672
rect 32397 498614 60076 498616
rect 32397 498611 32463 498614
rect 42149 498130 42215 498133
rect 42374 498130 42380 498132
rect 42149 498128 42380 498130
rect 42149 498072 42154 498128
rect 42210 498072 42380 498128
rect 42149 498070 42380 498072
rect 42149 498067 42215 498070
rect 42374 498068 42380 498070
rect 42444 498068 42450 498132
rect 57513 498130 57579 498133
rect 57513 498128 60076 498130
rect 57513 498072 57518 498128
rect 57574 498072 60076 498128
rect 57513 498070 60076 498072
rect 57513 498067 57579 498070
rect 583520 497844 584960 498084
rect 36486 497524 36492 497588
rect 36556 497586 36562 497588
rect 36556 497526 60076 497586
rect 36556 497524 36562 497526
rect 55990 497116 55996 497180
rect 56060 497178 56066 497180
rect 60273 497178 60339 497181
rect 56060 497176 60339 497178
rect 56060 497120 60278 497176
rect 60334 497120 60339 497176
rect 56060 497118 60339 497120
rect 56060 497116 56066 497118
rect 60273 497115 60339 497118
rect 42742 496980 42748 497044
rect 42812 497042 42818 497044
rect 42812 496982 60076 497042
rect 42812 496980 42818 496982
rect 43253 496770 43319 496773
rect 43478 496770 43484 496772
rect 43253 496768 43484 496770
rect 43253 496712 43258 496768
rect 43314 496712 43484 496768
rect 43253 496710 43484 496712
rect 43253 496707 43319 496710
rect 43478 496708 43484 496710
rect 43548 496708 43554 496772
rect 57646 496436 57652 496500
rect 57716 496498 57722 496500
rect 57716 496438 60076 496498
rect 57716 496436 57722 496438
rect 47577 496362 47643 496365
rect 57513 496362 57579 496365
rect 47577 496360 57579 496362
rect 47577 496304 47582 496360
rect 47638 496304 57518 496360
rect 57574 496304 57579 496360
rect 47577 496302 57579 496304
rect 47577 496299 47643 496302
rect 57513 496299 57579 496302
rect 46473 496226 46539 496229
rect 57697 496226 57763 496229
rect 46473 496224 57763 496226
rect 46473 496168 46478 496224
rect 46534 496168 57702 496224
rect 57758 496168 57763 496224
rect 46473 496166 57763 496168
rect 46473 496163 46539 496166
rect 57697 496163 57763 496166
rect 43161 496090 43227 496093
rect 57053 496090 57119 496093
rect 43161 496088 57119 496090
rect 43161 496032 43166 496088
rect 43222 496032 57058 496088
rect 57114 496032 57119 496088
rect 43161 496030 57119 496032
rect 43161 496027 43227 496030
rect 57053 496027 57119 496030
rect 32438 495892 32444 495956
rect 32508 495954 32514 495956
rect 32508 495894 60076 495954
rect 32508 495892 32514 495894
rect 35198 495348 35204 495412
rect 35268 495410 35274 495412
rect 35268 495350 60076 495410
rect 35268 495348 35274 495350
rect 40902 494804 40908 494868
rect 40972 494866 40978 494868
rect 40972 494806 60076 494866
rect 40972 494804 40978 494806
rect 39062 494668 39068 494732
rect 39132 494730 39138 494732
rect 39757 494730 39823 494733
rect 39132 494728 39823 494730
rect 39132 494672 39762 494728
rect 39818 494672 39823 494728
rect 39132 494670 39823 494672
rect 39132 494668 39138 494670
rect 39757 494667 39823 494670
rect 46422 494668 46428 494732
rect 46492 494730 46498 494732
rect 57278 494730 57284 494732
rect 46492 494670 57284 494730
rect 46492 494668 46498 494670
rect 57278 494668 57284 494670
rect 57348 494668 57354 494732
rect 39246 494260 39252 494324
rect 39316 494322 39322 494324
rect 39316 494262 60076 494322
rect 39316 494260 39322 494262
rect 44398 493988 44404 494052
rect 44468 494050 44474 494052
rect 45001 494050 45067 494053
rect 44468 494048 45067 494050
rect 44468 493992 45006 494048
rect 45062 493992 45067 494048
rect 44468 493990 45067 493992
rect 44468 493988 44474 493990
rect 45001 493987 45067 493990
rect 59670 493716 59676 493780
rect 59740 493778 59746 493780
rect 59740 493718 60076 493778
rect 59740 493716 59746 493718
rect 43437 493370 43503 493373
rect 57145 493370 57211 493373
rect 43437 493368 57211 493370
rect 43437 493312 43442 493368
rect 43498 493312 57150 493368
rect 57206 493312 57211 493368
rect 43437 493310 57211 493312
rect 43437 493307 43503 493310
rect 57145 493307 57211 493310
rect 44582 493172 44588 493236
rect 44652 493234 44658 493236
rect 44652 493174 60076 493234
rect 44652 493172 44658 493174
rect 57513 492690 57579 492693
rect 57513 492688 60076 492690
rect 57513 492632 57518 492688
rect 57574 492632 60076 492688
rect 57513 492630 60076 492632
rect 57513 492627 57579 492630
rect 35750 492084 35756 492148
rect 35820 492146 35826 492148
rect 35820 492086 60076 492146
rect 35820 492084 35826 492086
rect 37917 491874 37983 491877
rect 46054 491874 46060 491876
rect 37917 491872 46060 491874
rect 37917 491816 37922 491872
rect 37978 491816 46060 491872
rect 37917 491814 46060 491816
rect 37917 491811 37983 491814
rect 46054 491812 46060 491814
rect 46124 491812 46130 491876
rect 42558 491540 42564 491604
rect 42628 491602 42634 491604
rect 42628 491542 60076 491602
rect 42628 491540 42634 491542
rect 39246 491132 39252 491196
rect 39316 491194 39322 491196
rect 39849 491194 39915 491197
rect 39316 491192 39915 491194
rect 39316 491136 39854 491192
rect 39910 491136 39915 491192
rect 39316 491134 39915 491136
rect 39316 491132 39322 491134
rect 39849 491131 39915 491134
rect 57145 491194 57211 491197
rect 58801 491194 58867 491197
rect 57145 491192 58867 491194
rect 57145 491136 57150 491192
rect 57206 491136 58806 491192
rect 58862 491136 58867 491192
rect 57145 491134 58867 491136
rect 57145 491131 57211 491134
rect 58801 491131 58867 491134
rect 57697 491058 57763 491061
rect 57697 491056 60076 491058
rect 57697 491000 57702 491056
rect 57758 491000 60076 491056
rect 57697 490998 60076 491000
rect 57697 490995 57763 490998
rect 39430 490452 39436 490516
rect 39500 490514 39506 490516
rect 39500 490454 60076 490514
rect 39500 490452 39506 490454
rect 57053 489970 57119 489973
rect 57053 489968 60076 489970
rect 57053 489912 57058 489968
rect 57114 489912 60076 489968
rect 57053 489910 60076 489912
rect 57053 489907 57119 489910
rect 35382 489364 35388 489428
rect 35452 489426 35458 489428
rect 35452 489366 60076 489426
rect 35452 489364 35458 489366
rect 38009 488882 38075 488885
rect 38009 488880 60076 488882
rect -960 488596 480 488836
rect 38009 488824 38014 488880
rect 38070 488824 60076 488880
rect 38009 488822 60076 488824
rect 38009 488819 38075 488822
rect 30966 488276 30972 488340
rect 31036 488338 31042 488340
rect 31036 488278 60076 488338
rect 31036 488276 31042 488278
rect 499430 488276 499436 488340
rect 499500 488338 499506 488340
rect 500585 488338 500651 488341
rect 499500 488336 500651 488338
rect 499500 488280 500590 488336
rect 500646 488280 500651 488336
rect 499500 488278 500651 488280
rect 499500 488276 499506 488278
rect 500585 488275 500651 488278
rect 55806 487732 55812 487796
rect 55876 487794 55882 487796
rect 55876 487734 60076 487794
rect 55876 487732 55882 487734
rect 503621 487522 503687 487525
rect 499836 487520 503687 487522
rect 499836 487464 503626 487520
rect 503682 487464 503687 487520
rect 499836 487462 503687 487464
rect 503621 487459 503687 487462
rect 27470 487188 27476 487252
rect 27540 487250 27546 487252
rect 500217 487250 500283 487253
rect 27540 487190 60076 487250
rect 499836 487248 500283 487250
rect 499836 487192 500222 487248
rect 500278 487192 500283 487248
rect 499836 487190 500283 487192
rect 27540 487188 27546 487190
rect 500217 487187 500283 487190
rect 525149 486978 525215 486981
rect 499836 486976 525215 486978
rect 499836 486920 525154 486976
rect 525210 486920 525215 486976
rect 499836 486918 525215 486920
rect 525149 486915 525215 486918
rect 57605 486706 57671 486709
rect 532049 486706 532115 486709
rect 57605 486704 60076 486706
rect 57605 486648 57610 486704
rect 57666 486648 60076 486704
rect 57605 486646 60076 486648
rect 499836 486704 532115 486706
rect 499836 486648 532054 486704
rect 532110 486648 532115 486704
rect 499836 486646 532115 486648
rect 57605 486643 57671 486646
rect 532049 486643 532115 486646
rect 503069 486434 503135 486437
rect 499836 486432 503135 486434
rect 499836 486376 503074 486432
rect 503130 486376 503135 486432
rect 499836 486374 503135 486376
rect 503069 486371 503135 486374
rect 29678 486100 29684 486164
rect 29748 486162 29754 486164
rect 512637 486162 512703 486165
rect 29748 486102 60076 486162
rect 499836 486160 512703 486162
rect 499836 486104 512642 486160
rect 512698 486104 512703 486160
rect 499836 486102 512703 486104
rect 29748 486100 29754 486102
rect 512637 486099 512703 486102
rect 503161 485890 503227 485893
rect 499836 485888 503227 485890
rect 499836 485832 503166 485888
rect 503222 485832 503227 485888
rect 499836 485830 503227 485832
rect 503161 485827 503227 485830
rect 29862 485556 29868 485620
rect 29932 485618 29938 485620
rect 514201 485618 514267 485621
rect 29932 485558 60076 485618
rect 499836 485616 514267 485618
rect 499836 485560 514206 485616
rect 514262 485560 514267 485616
rect 499836 485558 514267 485560
rect 29932 485556 29938 485558
rect 514201 485555 514267 485558
rect 511349 485346 511415 485349
rect 499836 485344 511415 485346
rect 499836 485288 511354 485344
rect 511410 485288 511415 485344
rect 499836 485286 511415 485288
rect 511349 485283 511415 485286
rect 30046 485012 30052 485076
rect 30116 485074 30122 485076
rect 521101 485074 521167 485077
rect 30116 485014 60076 485074
rect 499836 485072 521167 485074
rect 499836 485016 521106 485072
rect 521162 485016 521167 485072
rect 499836 485014 521167 485016
rect 30116 485012 30122 485014
rect 521101 485011 521167 485014
rect 522246 484802 522252 484804
rect 499836 484742 522252 484802
rect 522246 484740 522252 484742
rect 522316 484740 522322 484804
rect 580574 484604 580580 484668
rect 580644 484666 580650 484668
rect 583520 484666 584960 484756
rect 580644 484606 584960 484666
rect 580644 484604 580650 484606
rect 33726 484468 33732 484532
rect 33796 484530 33802 484532
rect 502701 484530 502767 484533
rect 33796 484470 60076 484530
rect 499836 484528 502767 484530
rect 499836 484472 502706 484528
rect 502762 484472 502767 484528
rect 583520 484516 584960 484606
rect 499836 484470 502767 484472
rect 33796 484468 33802 484470
rect 502701 484467 502767 484470
rect 503621 484394 503687 484397
rect 505921 484394 505987 484397
rect 503621 484392 505987 484394
rect 503621 484336 503626 484392
rect 503682 484336 505926 484392
rect 505982 484336 505987 484392
rect 503621 484334 505987 484336
rect 503621 484331 503687 484334
rect 505921 484331 505987 484334
rect 508262 484258 508268 484260
rect 499836 484198 508268 484258
rect 508262 484196 508268 484198
rect 508332 484196 508338 484260
rect 36854 483924 36860 483988
rect 36924 483986 36930 483988
rect 501597 483986 501663 483989
rect 36924 483926 60076 483986
rect 499836 483984 501663 483986
rect 499836 483928 501602 483984
rect 501658 483928 501663 483984
rect 499836 483926 501663 483928
rect 36924 483924 36930 483926
rect 501597 483923 501663 483926
rect 502701 483986 502767 483989
rect 507158 483986 507164 483988
rect 502701 483984 507164 483986
rect 502701 483928 502706 483984
rect 502762 483928 507164 483984
rect 502701 483926 507164 483928
rect 502701 483923 502767 483926
rect 507158 483924 507164 483926
rect 507228 483924 507234 483988
rect 502609 483714 502675 483717
rect 499836 483712 502675 483714
rect 499836 483656 502614 483712
rect 502670 483656 502675 483712
rect 499836 483654 502675 483656
rect 502609 483651 502675 483654
rect 37222 483380 37228 483444
rect 37292 483442 37298 483444
rect 502517 483442 502583 483445
rect 37292 483382 60076 483442
rect 499836 483440 502583 483442
rect 499836 483384 502522 483440
rect 502578 483384 502583 483440
rect 499836 483382 502583 483384
rect 37292 483380 37298 483382
rect 502517 483379 502583 483382
rect 504541 483170 504607 483173
rect 499836 483168 504607 483170
rect 499836 483112 504546 483168
rect 504602 483112 504607 483168
rect 499836 483110 504607 483112
rect 504541 483107 504607 483110
rect 50613 483034 50679 483037
rect 50613 483032 50906 483034
rect 50613 482976 50618 483032
rect 50674 482976 50906 483032
rect 50613 482974 50906 482976
rect 50613 482971 50679 482974
rect 50286 482836 50292 482900
rect 50356 482898 50362 482900
rect 50613 482898 50679 482901
rect 50356 482896 50679 482898
rect 50356 482840 50618 482896
rect 50674 482840 50679 482896
rect 50356 482838 50679 482840
rect 50846 482898 50906 482974
rect 500217 482900 500283 482901
rect 50846 482838 60076 482898
rect 499836 482838 500050 482898
rect 50356 482836 50362 482838
rect 50613 482835 50679 482838
rect 499990 482762 500050 482838
rect 500166 482836 500172 482900
rect 500236 482898 500283 482900
rect 502793 482898 502859 482901
rect 500236 482896 500328 482898
rect 500278 482840 500328 482896
rect 500236 482838 500328 482840
rect 500542 482896 502859 482898
rect 500542 482840 502798 482896
rect 502854 482840 502859 482896
rect 500542 482838 502859 482840
rect 500236 482836 500283 482838
rect 500217 482835 500283 482836
rect 500542 482762 500602 482838
rect 502793 482835 502859 482838
rect 499990 482702 500602 482762
rect 502885 482626 502951 482629
rect 499836 482624 502951 482626
rect 499836 482568 502890 482624
rect 502946 482568 502951 482624
rect 499836 482566 502951 482568
rect 502885 482563 502951 482566
rect 51809 482354 51875 482357
rect 500493 482354 500559 482357
rect 51809 482352 60076 482354
rect 51809 482296 51814 482352
rect 51870 482296 60076 482352
rect 51809 482294 60076 482296
rect 499836 482352 500559 482354
rect 499836 482296 500498 482352
rect 500554 482296 500559 482352
rect 499836 482294 500559 482296
rect 51809 482291 51875 482294
rect 500493 482291 500559 482294
rect 500534 482156 500540 482220
rect 500604 482218 500610 482220
rect 512494 482218 512500 482220
rect 500604 482158 512500 482218
rect 500604 482156 500610 482158
rect 512494 482156 512500 482158
rect 512564 482156 512570 482220
rect 502333 482082 502399 482085
rect 499836 482080 502399 482082
rect 499836 482024 502338 482080
rect 502394 482024 502399 482080
rect 499836 482022 502399 482024
rect 502333 482019 502399 482022
rect 54753 481810 54819 481813
rect 503345 481810 503411 481813
rect 54753 481808 60076 481810
rect 54753 481752 54758 481808
rect 54814 481752 60076 481808
rect 54753 481750 60076 481752
rect 499836 481808 503411 481810
rect 499836 481752 503350 481808
rect 503406 481752 503411 481808
rect 499836 481750 503411 481752
rect 54753 481747 54819 481750
rect 503345 481747 503411 481750
rect 529238 481538 529244 481540
rect 499836 481478 529244 481538
rect 529238 481476 529244 481478
rect 529308 481476 529314 481540
rect 501454 481340 501460 481404
rect 501524 481402 501530 481404
rect 502333 481402 502399 481405
rect 501524 481400 502399 481402
rect 501524 481344 502338 481400
rect 502394 481344 502399 481400
rect 501524 481342 502399 481344
rect 501524 481340 501530 481342
rect 502333 481339 502399 481342
rect 503110 481340 503116 481404
rect 503180 481402 503186 481404
rect 503529 481402 503595 481405
rect 503180 481400 503595 481402
rect 503180 481344 503534 481400
rect 503590 481344 503595 481400
rect 503180 481342 503595 481344
rect 503180 481340 503186 481342
rect 503529 481339 503595 481342
rect 511349 481402 511415 481405
rect 512126 481402 512132 481404
rect 511349 481400 512132 481402
rect 511349 481344 511354 481400
rect 511410 481344 512132 481400
rect 511349 481342 512132 481344
rect 511349 481339 511415 481342
rect 512126 481340 512132 481342
rect 512196 481340 512202 481404
rect 25681 481266 25747 481269
rect 518382 481266 518388 481268
rect 25681 481264 60076 481266
rect 25681 481208 25686 481264
rect 25742 481208 60076 481264
rect 25681 481206 60076 481208
rect 499836 481206 518388 481266
rect 25681 481203 25747 481206
rect 518382 481204 518388 481206
rect 518452 481204 518458 481268
rect 503253 480994 503319 480997
rect 499836 480992 503319 480994
rect 499836 480936 503258 480992
rect 503314 480936 503319 480992
rect 499836 480934 503319 480936
rect 503253 480931 503319 480934
rect 512637 480858 512703 480861
rect 526294 480858 526300 480860
rect 512637 480856 526300 480858
rect 512637 480800 512642 480856
rect 512698 480800 526300 480856
rect 512637 480798 526300 480800
rect 512637 480795 512703 480798
rect 526294 480796 526300 480798
rect 526364 480796 526370 480860
rect 31293 480722 31359 480725
rect 534257 480722 534323 480725
rect 31293 480720 60076 480722
rect 31293 480664 31298 480720
rect 31354 480664 60076 480720
rect 31293 480662 60076 480664
rect 499836 480720 534323 480722
rect 499836 480664 534262 480720
rect 534318 480664 534323 480720
rect 499836 480662 534323 480664
rect 31293 480659 31359 480662
rect 534257 480659 534323 480662
rect 502558 480450 502564 480452
rect 499836 480390 502564 480450
rect 502558 480388 502564 480390
rect 502628 480388 502634 480452
rect 505829 480314 505895 480317
rect 511206 480314 511212 480316
rect 505829 480312 511212 480314
rect 505829 480256 505834 480312
rect 505890 480256 511212 480312
rect 505829 480254 511212 480256
rect 505829 480251 505895 480254
rect 511206 480252 511212 480254
rect 511276 480252 511282 480316
rect 35709 480178 35775 480181
rect 502374 480178 502380 480180
rect 35709 480176 60076 480178
rect 35709 480120 35714 480176
rect 35770 480120 60076 480176
rect 35709 480118 60076 480120
rect 499836 480118 502380 480178
rect 35709 480115 35775 480118
rect 502374 480116 502380 480118
rect 502444 480116 502450 480180
rect 501413 479906 501479 479909
rect 499836 479904 501479 479906
rect 499836 479848 501418 479904
rect 501474 479848 501479 479904
rect 499836 479846 501479 479848
rect 501413 479843 501479 479846
rect 56225 479634 56291 479637
rect 504449 479634 504515 479637
rect 56225 479632 60076 479634
rect 56225 479576 56230 479632
rect 56286 479576 60076 479632
rect 56225 479574 60076 479576
rect 499836 479632 504515 479634
rect 499836 479576 504454 479632
rect 504510 479576 504515 479632
rect 499836 479574 504515 479576
rect 56225 479571 56291 479574
rect 504449 479571 504515 479574
rect 502742 479362 502748 479364
rect 499836 479302 502748 479362
rect 502742 479300 502748 479302
rect 502812 479300 502818 479364
rect 42517 479090 42583 479093
rect 502926 479090 502932 479092
rect 42517 479088 60076 479090
rect 42517 479032 42522 479088
rect 42578 479032 60076 479088
rect 42517 479030 60076 479032
rect 499836 479030 502932 479090
rect 42517 479027 42583 479030
rect 502926 479028 502932 479030
rect 502996 479028 503002 479092
rect 55990 478892 55996 478956
rect 56060 478954 56066 478956
rect 56225 478954 56291 478957
rect 56060 478952 56291 478954
rect 56060 478896 56230 478952
rect 56286 478896 56291 478952
rect 56060 478894 56291 478896
rect 56060 478892 56066 478894
rect 56225 478891 56291 478894
rect 505134 478818 505140 478820
rect 499836 478758 505140 478818
rect 505134 478756 505140 478758
rect 505204 478756 505210 478820
rect 53557 478546 53623 478549
rect 519486 478546 519492 478548
rect 53557 478544 60076 478546
rect 53557 478488 53562 478544
rect 53618 478488 60076 478544
rect 53557 478486 60076 478488
rect 499836 478486 519492 478546
rect 53557 478483 53623 478486
rect 519486 478484 519492 478486
rect 519556 478484 519562 478548
rect 516358 478274 516364 478276
rect 499836 478214 516364 478274
rect 516358 478212 516364 478214
rect 516428 478212 516434 478276
rect 54845 478002 54911 478005
rect 511022 478002 511028 478004
rect 54845 478000 60076 478002
rect 54845 477944 54850 478000
rect 54906 477944 60076 478000
rect 54845 477942 60076 477944
rect 499836 477942 511028 478002
rect 54845 477939 54911 477942
rect 511022 477940 511028 477942
rect 511092 477940 511098 478004
rect 527398 477730 527404 477732
rect 499836 477670 527404 477730
rect 527398 477668 527404 477670
rect 527468 477668 527474 477732
rect 38469 477458 38535 477461
rect 532734 477458 532740 477460
rect 38469 477456 60076 477458
rect 38469 477400 38474 477456
rect 38530 477400 60076 477456
rect 38469 477398 60076 477400
rect 499836 477398 532740 477458
rect 38469 477395 38535 477398
rect 532734 477396 532740 477398
rect 532804 477396 532810 477460
rect 509693 477186 509759 477189
rect 499836 477184 509759 477186
rect 499836 477128 509698 477184
rect 509754 477128 509759 477184
rect 499836 477126 509759 477128
rect 509693 477123 509759 477126
rect 52085 476914 52151 476917
rect 534022 476914 534028 476916
rect 52085 476912 60076 476914
rect 52085 476856 52090 476912
rect 52146 476856 60076 476912
rect 52085 476854 60076 476856
rect 499836 476854 534028 476914
rect 52085 476851 52151 476854
rect 534022 476852 534028 476854
rect 534092 476852 534098 476916
rect 539726 476642 539732 476644
rect 499836 476582 539732 476642
rect 539726 476580 539732 476582
rect 539796 476580 539802 476644
rect 51901 476370 51967 476373
rect 525374 476370 525380 476372
rect 51901 476368 60076 476370
rect 51901 476312 51906 476368
rect 51962 476312 60076 476368
rect 51901 476310 60076 476312
rect 499836 476310 525380 476370
rect 51901 476307 51967 476310
rect 525374 476308 525380 476310
rect 525444 476308 525450 476372
rect 51574 476172 51580 476236
rect 51644 476234 51650 476236
rect 52361 476234 52427 476237
rect 51644 476232 52427 476234
rect 51644 476176 52366 476232
rect 52422 476176 52427 476232
rect 51644 476174 52427 476176
rect 51644 476172 51650 476174
rect 52361 476171 52427 476174
rect 540421 476234 540487 476237
rect 544561 476234 544627 476237
rect 540421 476232 544627 476234
rect 540421 476176 540426 476232
rect 540482 476176 544566 476232
rect 544622 476176 544627 476232
rect 540421 476174 544627 476176
rect 540421 476171 540487 476174
rect 544561 476171 544627 476174
rect 514109 476098 514175 476101
rect 499836 476096 514175 476098
rect 499836 476040 514114 476096
rect 514170 476040 514175 476096
rect 499836 476038 514175 476040
rect 514109 476035 514175 476038
rect 25865 475826 25931 475829
rect 505318 475826 505324 475828
rect 25865 475824 60076 475826
rect -960 475690 480 475780
rect 25865 475768 25870 475824
rect 25926 475768 60076 475824
rect 25865 475766 60076 475768
rect 499836 475766 505324 475826
rect 25865 475763 25931 475766
rect 505318 475764 505324 475766
rect 505388 475764 505394 475828
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 44817 475554 44883 475557
rect 51901 475554 51967 475557
rect 522297 475554 522363 475557
rect 44817 475552 51967 475554
rect 44817 475496 44822 475552
rect 44878 475496 51906 475552
rect 51962 475496 51967 475552
rect 44817 475494 51967 475496
rect 499836 475552 522363 475554
rect 499836 475496 522302 475552
rect 522358 475496 522363 475552
rect 499836 475494 522363 475496
rect 44817 475491 44883 475494
rect 51901 475491 51967 475494
rect 522297 475491 522363 475494
rect 46054 475356 46060 475420
rect 46124 475418 46130 475420
rect 54334 475418 54340 475420
rect 46124 475358 54340 475418
rect 46124 475356 46130 475358
rect 54334 475356 54340 475358
rect 54404 475356 54410 475420
rect 53373 475282 53439 475285
rect 500350 475282 500356 475284
rect 53373 475280 60076 475282
rect 53373 475224 53378 475280
rect 53434 475224 60076 475280
rect 53373 475222 60076 475224
rect 499836 475222 500356 475282
rect 53373 475219 53439 475222
rect 500350 475220 500356 475222
rect 500420 475220 500426 475284
rect 508446 475010 508452 475012
rect 499836 474950 508452 475010
rect 508446 474948 508452 474950
rect 508516 474948 508522 475012
rect 52177 474738 52243 474741
rect 530158 474738 530164 474740
rect 52177 474736 60076 474738
rect 52177 474680 52182 474736
rect 52238 474680 60076 474736
rect 52177 474678 60076 474680
rect 499836 474678 530164 474738
rect 52177 474675 52243 474678
rect 530158 474676 530164 474678
rect 530228 474676 530234 474740
rect 500217 474602 500283 474605
rect 500350 474602 500356 474604
rect 500217 474600 500356 474602
rect 500217 474544 500222 474600
rect 500278 474544 500356 474600
rect 500217 474542 500356 474544
rect 500217 474539 500283 474542
rect 500350 474540 500356 474542
rect 500420 474540 500426 474604
rect 500493 474602 500559 474605
rect 501689 474602 501755 474605
rect 500493 474600 501755 474602
rect 500493 474544 500498 474600
rect 500554 474544 501694 474600
rect 501750 474544 501755 474600
rect 500493 474542 501755 474544
rect 500493 474539 500559 474542
rect 501689 474539 501755 474542
rect 531446 474466 531452 474468
rect 499836 474406 531452 474466
rect 531446 474404 531452 474406
rect 531516 474404 531522 474468
rect 52269 474194 52335 474197
rect 536966 474194 536972 474196
rect 52269 474192 60076 474194
rect 52269 474136 52274 474192
rect 52330 474136 60076 474192
rect 52269 474134 60076 474136
rect 499836 474134 536972 474194
rect 52269 474131 52335 474134
rect 536966 474132 536972 474134
rect 537036 474132 537042 474196
rect 514150 473922 514156 473924
rect 499836 473862 514156 473922
rect 514150 473860 514156 473862
rect 514220 473860 514226 473924
rect 56409 473650 56475 473653
rect 529054 473650 529060 473652
rect 56409 473648 60076 473650
rect 56409 473592 56414 473648
rect 56470 473592 60076 473648
rect 56409 473590 60076 473592
rect 499836 473590 529060 473650
rect 56409 473587 56475 473590
rect 529054 473588 529060 473590
rect 529124 473588 529130 473652
rect 519302 473378 519308 473380
rect 499836 473318 519308 473378
rect 519302 473316 519308 473318
rect 519372 473316 519378 473380
rect 538622 473180 538628 473244
rect 538692 473242 538698 473244
rect 539501 473242 539567 473245
rect 538692 473240 539567 473242
rect 538692 473184 539506 473240
rect 539562 473184 539567 473240
rect 538692 473182 539567 473184
rect 538692 473180 538698 473182
rect 539501 473179 539567 473182
rect 41229 473106 41295 473109
rect 520406 473106 520412 473108
rect 41229 473104 60076 473106
rect 41229 473048 41234 473104
rect 41290 473048 60076 473104
rect 41229 473046 60076 473048
rect 499836 473046 520412 473106
rect 41229 473043 41295 473046
rect 520406 473044 520412 473046
rect 520476 473044 520482 473108
rect 512310 472834 512316 472836
rect 499836 472774 512316 472834
rect 512310 472772 512316 472774
rect 512380 472772 512386 472836
rect 44909 472698 44975 472701
rect 52177 472698 52243 472701
rect 44909 472696 52243 472698
rect 44909 472640 44914 472696
rect 44970 472640 52182 472696
rect 52238 472640 52243 472696
rect 44909 472638 52243 472640
rect 44909 472635 44975 472638
rect 52177 472635 52243 472638
rect 51993 472562 52059 472565
rect 539542 472562 539548 472564
rect 51993 472560 60076 472562
rect 51993 472504 51998 472560
rect 52054 472504 60076 472560
rect 51993 472502 60076 472504
rect 499836 472502 539548 472562
rect 51993 472499 52059 472502
rect 539542 472500 539548 472502
rect 539612 472500 539618 472564
rect 507301 472290 507367 472293
rect 499836 472288 507367 472290
rect 499836 472232 507306 472288
rect 507362 472232 507367 472288
rect 499836 472230 507367 472232
rect 507301 472227 507367 472230
rect 43989 472018 44055 472021
rect 538438 472018 538444 472020
rect 43989 472016 60076 472018
rect 43989 471960 43994 472016
rect 44050 471960 60076 472016
rect 43989 471958 60076 471960
rect 499836 471958 538444 472018
rect 43989 471955 44055 471958
rect 538438 471956 538444 471958
rect 538508 471956 538514 472020
rect 535678 471746 535684 471748
rect 499836 471686 535684 471746
rect 535678 471684 535684 471686
rect 535748 471684 535754 471748
rect 26049 471474 26115 471477
rect 515397 471474 515463 471477
rect 26049 471472 60076 471474
rect 26049 471416 26054 471472
rect 26110 471416 60076 471472
rect 26049 471414 60076 471416
rect 499836 471472 515463 471474
rect 499836 471416 515402 471472
rect 515458 471416 515463 471472
rect 499836 471414 515463 471416
rect 26049 471411 26115 471414
rect 515397 471411 515463 471414
rect 547086 471412 547092 471476
rect 547156 471474 547162 471476
rect 583520 471474 584960 471564
rect 547156 471414 584960 471474
rect 547156 471412 547162 471414
rect 583520 471324 584960 471414
rect 515489 471202 515555 471205
rect 499836 471200 515555 471202
rect 499836 471144 515494 471200
rect 515550 471144 515555 471200
rect 499836 471142 515555 471144
rect 515489 471139 515555 471142
rect 54109 470930 54175 470933
rect 514518 470930 514524 470932
rect 54109 470928 60076 470930
rect 54109 470872 54114 470928
rect 54170 470872 60076 470928
rect 54109 470870 60076 470872
rect 499836 470870 514524 470930
rect 54109 470867 54175 470870
rect 514518 470868 514524 470870
rect 514588 470868 514594 470932
rect 515254 470658 515260 470660
rect 499836 470598 515260 470658
rect 515254 470596 515260 470598
rect 515324 470596 515330 470660
rect 53005 470386 53071 470389
rect 526110 470386 526116 470388
rect 53005 470384 60076 470386
rect 53005 470328 53010 470384
rect 53066 470328 60076 470384
rect 53005 470326 60076 470328
rect 499836 470326 526116 470386
rect 53005 470323 53071 470326
rect 526110 470324 526116 470326
rect 526180 470324 526186 470388
rect 523166 470114 523172 470116
rect 499836 470054 523172 470114
rect 523166 470052 523172 470054
rect 523236 470052 523242 470116
rect 42701 469842 42767 469845
rect 516174 469842 516180 469844
rect 42701 469840 60076 469842
rect 42701 469784 42706 469840
rect 42762 469784 60076 469840
rect 42701 469782 60076 469784
rect 499836 469782 516180 469842
rect 42701 469779 42767 469782
rect 516174 469780 516180 469782
rect 516244 469780 516250 469844
rect 518341 469570 518407 469573
rect 499836 469568 518407 469570
rect 499836 469512 518346 469568
rect 518402 469512 518407 469568
rect 499836 469510 518407 469512
rect 518341 469507 518407 469510
rect 32857 469298 32923 469301
rect 502885 469298 502951 469301
rect 32857 469296 60076 469298
rect 32857 469240 32862 469296
rect 32918 469240 60076 469296
rect 32857 469238 60076 469240
rect 499836 469296 502951 469298
rect 499836 469240 502890 469296
rect 502946 469240 502951 469296
rect 499836 469238 502951 469240
rect 32857 469235 32923 469238
rect 502885 469235 502951 469238
rect 531957 469026 532023 469029
rect 499836 469024 532023 469026
rect 499836 468968 531962 469024
rect 532018 468968 532023 469024
rect 499836 468966 532023 468968
rect 531957 468963 532023 468966
rect 56317 468754 56383 468757
rect 533429 468754 533495 468757
rect 56317 468752 60076 468754
rect 56317 468696 56322 468752
rect 56378 468696 60076 468752
rect 56317 468694 60076 468696
rect 499836 468752 533495 468754
rect 499836 468696 533434 468752
rect 533490 468696 533495 468752
rect 499836 468694 533495 468696
rect 56317 468691 56383 468694
rect 533429 468691 533495 468694
rect 502885 468482 502951 468485
rect 499836 468480 502951 468482
rect 499836 468424 502890 468480
rect 502946 468424 502951 468480
rect 499836 468422 502951 468424
rect 502885 468419 502951 468422
rect 534993 468482 535059 468485
rect 540421 468482 540487 468485
rect 534993 468480 540487 468482
rect 534993 468424 534998 468480
rect 535054 468424 540426 468480
rect 540482 468424 540487 468480
rect 534993 468422 540487 468424
rect 534993 468419 535059 468422
rect 540421 468419 540487 468422
rect 30005 468210 30071 468213
rect 502793 468210 502859 468213
rect 30005 468208 60076 468210
rect 30005 468152 30010 468208
rect 30066 468152 60076 468208
rect 30005 468150 60076 468152
rect 499836 468208 502859 468210
rect 499836 468152 502798 468208
rect 502854 468152 502859 468208
rect 499836 468150 502859 468152
rect 30005 468147 30071 468150
rect 502793 468147 502859 468150
rect 523769 468074 523835 468077
rect 509190 468072 523835 468074
rect 509190 468016 523774 468072
rect 523830 468016 523835 468072
rect 509190 468014 523835 468016
rect 509190 467938 509250 468014
rect 523769 468011 523835 468014
rect 499836 467878 509250 467938
rect 523534 467876 523540 467940
rect 523604 467938 523610 467940
rect 523953 467938 524019 467941
rect 523604 467936 524019 467938
rect 523604 467880 523958 467936
rect 524014 467880 524019 467936
rect 523604 467878 524019 467880
rect 523604 467876 523610 467878
rect 523953 467875 524019 467878
rect 28533 467666 28599 467669
rect 526437 467666 526503 467669
rect 28533 467664 60076 467666
rect 28533 467608 28538 467664
rect 28594 467608 60076 467664
rect 28533 467606 60076 467608
rect 499836 467664 526503 467666
rect 499836 467608 526442 467664
rect 526498 467608 526503 467664
rect 499836 467606 526503 467608
rect 28533 467603 28599 467606
rect 526437 467603 526503 467606
rect 502885 467394 502951 467397
rect 499836 467392 502951 467394
rect 499836 467336 502890 467392
rect 502946 467336 502951 467392
rect 499836 467334 502951 467336
rect 502885 467331 502951 467334
rect 34329 467122 34395 467125
rect 533521 467122 533587 467125
rect 34329 467120 60076 467122
rect 34329 467064 34334 467120
rect 34390 467064 60076 467120
rect 34329 467062 60076 467064
rect 499836 467120 533587 467122
rect 499836 467064 533526 467120
rect 533582 467064 533587 467120
rect 499836 467062 533587 467064
rect 34329 467059 34395 467062
rect 533521 467059 533587 467062
rect 502701 466850 502767 466853
rect 499836 466848 502767 466850
rect 499836 466792 502706 466848
rect 502762 466792 502767 466848
rect 499836 466790 502767 466792
rect 502701 466787 502767 466790
rect 55581 466578 55647 466581
rect 502793 466578 502859 466581
rect 55581 466576 60076 466578
rect 55581 466520 55586 466576
rect 55642 466520 60076 466576
rect 55581 466518 60076 466520
rect 499836 466576 502859 466578
rect 499836 466520 502798 466576
rect 502854 466520 502859 466576
rect 499836 466518 502859 466520
rect 55581 466515 55647 466518
rect 502793 466515 502859 466518
rect 502885 466306 502951 466309
rect 499836 466304 502951 466306
rect 499836 466248 502890 466304
rect 502946 466248 502951 466304
rect 499836 466246 502951 466248
rect 502885 466243 502951 466246
rect 54937 466034 55003 466037
rect 502701 466034 502767 466037
rect 54937 466032 60076 466034
rect 54937 465976 54942 466032
rect 54998 465976 60076 466032
rect 54937 465974 60076 465976
rect 499836 466032 502767 466034
rect 499836 465976 502706 466032
rect 502762 465976 502767 466032
rect 499836 465974 502767 465976
rect 54937 465971 55003 465974
rect 502701 465971 502767 465974
rect 502793 465762 502859 465765
rect 499836 465760 502859 465762
rect 499836 465704 502798 465760
rect 502854 465704 502859 465760
rect 499836 465702 502859 465704
rect 502793 465699 502859 465702
rect 51441 465490 51507 465493
rect 502609 465490 502675 465493
rect 51441 465488 60076 465490
rect 51441 465432 51446 465488
rect 51502 465432 60076 465488
rect 51441 465430 60076 465432
rect 499836 465488 502675 465490
rect 499836 465432 502614 465488
rect 502670 465432 502675 465488
rect 499836 465430 502675 465432
rect 51441 465427 51507 465430
rect 502609 465427 502675 465430
rect 534809 465218 534875 465221
rect 499836 465216 534875 465218
rect 499836 465160 534814 465216
rect 534870 465160 534875 465216
rect 499836 465158 534875 465160
rect 534809 465155 534875 465158
rect 32949 464946 33015 464949
rect 531865 464946 531931 464949
rect 32949 464944 60076 464946
rect 32949 464888 32954 464944
rect 33010 464888 60076 464944
rect 32949 464886 60076 464888
rect 499836 464944 531931 464946
rect 499836 464888 531870 464944
rect 531926 464888 531931 464944
rect 499836 464886 531931 464888
rect 32949 464883 33015 464886
rect 531865 464883 531931 464886
rect 531773 464674 531839 464677
rect 499836 464672 531839 464674
rect 499836 464616 531778 464672
rect 531834 464616 531839 464672
rect 499836 464614 531839 464616
rect 531773 464611 531839 464614
rect 50705 464402 50771 464405
rect 519721 464402 519787 464405
rect 50705 464400 60076 464402
rect 50705 464344 50710 464400
rect 50766 464344 60076 464400
rect 50705 464342 60076 464344
rect 499836 464400 519787 464402
rect 499836 464344 519726 464400
rect 519782 464344 519787 464400
rect 499836 464342 519787 464344
rect 50705 464339 50771 464342
rect 519721 464339 519787 464342
rect 502885 464130 502951 464133
rect 499836 464128 502951 464130
rect 499836 464072 502890 464128
rect 502946 464072 502951 464128
rect 499836 464070 502951 464072
rect 502885 464067 502951 464070
rect 52913 463858 52979 463861
rect 527725 463858 527791 463861
rect 52913 463856 60076 463858
rect 52913 463800 52918 463856
rect 52974 463800 60076 463856
rect 52913 463798 60076 463800
rect 499836 463856 527791 463858
rect 499836 463800 527730 463856
rect 527786 463800 527791 463856
rect 499836 463798 527791 463800
rect 52913 463795 52979 463798
rect 527725 463795 527791 463798
rect 523677 463586 523743 463589
rect 499836 463584 523743 463586
rect 499836 463528 523682 463584
rect 523738 463528 523743 463584
rect 499836 463526 523743 463528
rect 523677 463523 523743 463526
rect 50061 463314 50127 463317
rect 502701 463314 502767 463317
rect 50061 463312 60076 463314
rect 50061 463256 50066 463312
rect 50122 463256 60076 463312
rect 50061 463254 60076 463256
rect 499836 463312 502767 463314
rect 499836 463256 502706 463312
rect 502762 463256 502767 463312
rect 499836 463254 502767 463256
rect 50061 463251 50127 463254
rect 502701 463251 502767 463254
rect 502885 463042 502951 463045
rect 499836 463040 502951 463042
rect 499836 462984 502890 463040
rect 502946 462984 502951 463040
rect 499836 462982 502951 462984
rect 502885 462979 502951 462982
rect 37181 462770 37247 462773
rect 502793 462770 502859 462773
rect 37181 462768 60076 462770
rect -960 462634 480 462724
rect 37181 462712 37186 462768
rect 37242 462712 60076 462768
rect 37181 462710 60076 462712
rect 499836 462768 502859 462770
rect 499836 462712 502798 462768
rect 502854 462712 502859 462768
rect 499836 462710 502859 462712
rect 37181 462707 37247 462710
rect 502793 462707 502859 462710
rect 3366 462634 3372 462636
rect -960 462574 3372 462634
rect -960 462484 480 462574
rect 3366 462572 3372 462574
rect 3436 462572 3442 462636
rect 502609 462498 502675 462501
rect 499836 462496 502675 462498
rect 499836 462440 502614 462496
rect 502670 462440 502675 462496
rect 499836 462438 502675 462440
rect 502609 462435 502675 462438
rect 50889 462226 50955 462229
rect 502885 462226 502951 462229
rect 50889 462224 60076 462226
rect 50889 462168 50894 462224
rect 50950 462168 60076 462224
rect 50889 462166 60076 462168
rect 499836 462224 502951 462226
rect 499836 462168 502890 462224
rect 502946 462168 502951 462224
rect 499836 462166 502951 462168
rect 50889 462163 50955 462166
rect 502885 462163 502951 462166
rect 502517 461954 502583 461957
rect 499836 461952 502583 461954
rect 499836 461896 502522 461952
rect 502578 461896 502583 461952
rect 499836 461894 502583 461896
rect 502517 461891 502583 461894
rect 41321 461682 41387 461685
rect 502885 461682 502951 461685
rect 41321 461680 60076 461682
rect 41321 461624 41326 461680
rect 41382 461624 60076 461680
rect 41321 461622 60076 461624
rect 499836 461680 502951 461682
rect 499836 461624 502890 461680
rect 502946 461624 502951 461680
rect 499836 461622 502951 461624
rect 41321 461619 41387 461622
rect 502885 461619 502951 461622
rect 502609 461410 502675 461413
rect 499836 461408 502675 461410
rect 499836 461352 502614 461408
rect 502670 461352 502675 461408
rect 499836 461350 502675 461352
rect 502609 461347 502675 461350
rect 28717 461138 28783 461141
rect 502793 461138 502859 461141
rect 28717 461136 60076 461138
rect 28717 461080 28722 461136
rect 28778 461080 60076 461136
rect 28717 461078 60076 461080
rect 499836 461136 502859 461138
rect 499836 461080 502798 461136
rect 502854 461080 502859 461136
rect 499836 461078 502859 461080
rect 28717 461075 28783 461078
rect 502793 461075 502859 461078
rect 533061 460866 533127 460869
rect 499836 460864 533127 460866
rect 499836 460808 533066 460864
rect 533122 460808 533127 460864
rect 499836 460806 533127 460808
rect 533061 460803 533127 460806
rect 28809 460594 28875 460597
rect 502793 460594 502859 460597
rect 28809 460592 60076 460594
rect 28809 460536 28814 460592
rect 28870 460536 60076 460592
rect 28809 460534 60076 460536
rect 499836 460592 502859 460594
rect 499836 460536 502798 460592
rect 502854 460536 502859 460592
rect 499836 460534 502859 460536
rect 28809 460531 28875 460534
rect 502793 460531 502859 460534
rect 502885 460322 502951 460325
rect 499836 460320 502951 460322
rect 499836 460264 502890 460320
rect 502946 460264 502951 460320
rect 499836 460262 502951 460264
rect 502885 460259 502951 460262
rect 536373 460186 536439 460189
rect 544377 460186 544443 460189
rect 536373 460184 544443 460186
rect 536373 460128 536378 460184
rect 536434 460128 544382 460184
rect 544438 460128 544443 460184
rect 536373 460126 544443 460128
rect 536373 460123 536439 460126
rect 544377 460123 544443 460126
rect 54293 460050 54359 460053
rect 536189 460050 536255 460053
rect 54293 460048 60076 460050
rect 54293 459992 54298 460048
rect 54354 459992 60076 460048
rect 54293 459990 60076 459992
rect 499836 460048 536255 460050
rect 499836 459992 536194 460048
rect 536250 459992 536255 460048
rect 499836 459990 536255 459992
rect 54293 459987 54359 459990
rect 536189 459987 536255 459990
rect 534349 459778 534415 459781
rect 499836 459776 534415 459778
rect 499836 459720 534354 459776
rect 534410 459720 534415 459776
rect 499836 459718 534415 459720
rect 534349 459715 534415 459718
rect 49601 459506 49667 459509
rect 535913 459506 535979 459509
rect 49601 459504 60076 459506
rect 49601 459448 49606 459504
rect 49662 459448 60076 459504
rect 49601 459446 60076 459448
rect 499836 459504 535979 459506
rect 499836 459448 535918 459504
rect 535974 459448 535979 459504
rect 499836 459446 535979 459448
rect 49601 459443 49667 459446
rect 535913 459443 535979 459446
rect 502885 459234 502951 459237
rect 499836 459232 502951 459234
rect 499836 459176 502890 459232
rect 502946 459176 502951 459232
rect 499836 459174 502951 459176
rect 502885 459171 502951 459174
rect 48037 458962 48103 458965
rect 502609 458962 502675 458965
rect 48037 458960 60076 458962
rect 48037 458904 48042 458960
rect 48098 458904 60076 458960
rect 48037 458902 60076 458904
rect 499836 458960 502675 458962
rect 499836 458904 502614 458960
rect 502670 458904 502675 458960
rect 499836 458902 502675 458904
rect 48037 458899 48103 458902
rect 502609 458899 502675 458902
rect 502793 458690 502859 458693
rect 499836 458688 502859 458690
rect 499836 458632 502798 458688
rect 502854 458632 502859 458688
rect 499836 458630 502859 458632
rect 502793 458627 502859 458630
rect 46790 458356 46796 458420
rect 46860 458418 46866 458420
rect 502701 458418 502767 458421
rect 46860 458358 60076 458418
rect 499836 458416 502767 458418
rect 499836 458360 502706 458416
rect 502762 458360 502767 458416
rect 499836 458358 502767 458360
rect 46860 458356 46866 458358
rect 502701 458355 502767 458358
rect 502885 458146 502951 458149
rect 499836 458144 502951 458146
rect 499836 458088 502890 458144
rect 502946 458088 502951 458144
rect 499836 458086 502951 458088
rect 502885 458083 502951 458086
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 48630 457812 48636 457876
rect 48700 457874 48706 457876
rect 502793 457874 502859 457877
rect 48700 457814 60076 457874
rect 499836 457872 502859 457874
rect 499836 457816 502798 457872
rect 502854 457816 502859 457872
rect 499836 457814 502859 457816
rect 48700 457812 48706 457814
rect 502793 457811 502859 457814
rect 514017 457602 514083 457605
rect 499836 457600 514083 457602
rect 499836 457544 514022 457600
rect 514078 457544 514083 457600
rect 499836 457542 514083 457544
rect 514017 457539 514083 457542
rect 48221 457330 48287 457333
rect 502701 457330 502767 457333
rect 48221 457328 60076 457330
rect 48221 457272 48226 457328
rect 48282 457272 60076 457328
rect 48221 457270 60076 457272
rect 499836 457328 502767 457330
rect 499836 457272 502706 457328
rect 502762 457272 502767 457328
rect 499836 457270 502767 457272
rect 48221 457267 48287 457270
rect 502701 457267 502767 457270
rect 502609 457058 502675 457061
rect 499836 457056 502675 457058
rect 499836 457000 502614 457056
rect 502670 457000 502675 457056
rect 499836 456998 502675 457000
rect 502609 456995 502675 456998
rect 48129 456786 48195 456789
rect 502885 456786 502951 456789
rect 48129 456784 60076 456786
rect 48129 456728 48134 456784
rect 48190 456728 60076 456784
rect 48129 456726 60076 456728
rect 499836 456784 502951 456786
rect 499836 456728 502890 456784
rect 502946 456728 502951 456784
rect 499836 456726 502951 456728
rect 48129 456723 48195 456726
rect 502885 456723 502951 456726
rect 502885 456514 502951 456517
rect 499836 456512 502951 456514
rect 499836 456456 502890 456512
rect 502946 456456 502951 456512
rect 499836 456454 502951 456456
rect 502885 456451 502951 456454
rect 54886 456180 54892 456244
rect 54956 456242 54962 456244
rect 516685 456242 516751 456245
rect 54956 456182 60076 456242
rect 499836 456240 516751 456242
rect 499836 456184 516690 456240
rect 516746 456184 516751 456240
rect 499836 456182 516751 456184
rect 54956 456180 54962 456182
rect 516685 456179 516751 456182
rect 502793 455970 502859 455973
rect 499836 455968 502859 455970
rect 499836 455912 502798 455968
rect 502854 455912 502859 455968
rect 499836 455910 502859 455912
rect 502793 455907 502859 455910
rect 47894 455636 47900 455700
rect 47964 455698 47970 455700
rect 502609 455698 502675 455701
rect 47964 455638 60076 455698
rect 499836 455696 502675 455698
rect 499836 455640 502614 455696
rect 502670 455640 502675 455696
rect 499836 455638 502675 455640
rect 47964 455636 47970 455638
rect 502609 455635 502675 455638
rect 502793 455426 502859 455429
rect 499836 455424 502859 455426
rect 499836 455368 502798 455424
rect 502854 455368 502859 455424
rect 499836 455366 502859 455368
rect 502793 455363 502859 455366
rect 47710 455092 47716 455156
rect 47780 455154 47786 455156
rect 502885 455154 502951 455157
rect 47780 455094 60076 455154
rect 499836 455152 502951 455154
rect 499836 455096 502890 455152
rect 502946 455096 502951 455152
rect 499836 455094 502951 455096
rect 47780 455092 47786 455094
rect 502885 455091 502951 455094
rect 502701 454882 502767 454885
rect 499836 454880 502767 454882
rect 499836 454824 502706 454880
rect 502762 454824 502767 454880
rect 499836 454822 502767 454824
rect 502701 454819 502767 454822
rect 48446 454548 48452 454612
rect 48516 454610 48522 454612
rect 501270 454610 501276 454612
rect 48516 454550 60076 454610
rect 499836 454550 501276 454610
rect 48516 454548 48522 454550
rect 501270 454548 501276 454550
rect 501340 454548 501346 454612
rect 502609 454338 502675 454341
rect 499836 454336 502675 454338
rect 499836 454280 502614 454336
rect 502670 454280 502675 454336
rect 499836 454278 502675 454280
rect 502609 454275 502675 454278
rect 33910 454004 33916 454068
rect 33980 454066 33986 454068
rect 502517 454066 502583 454069
rect 33980 454006 60076 454066
rect 499836 454064 502583 454066
rect 499836 454008 502522 454064
rect 502578 454008 502583 454064
rect 499836 454006 502583 454008
rect 33980 454004 33986 454006
rect 502517 454003 502583 454006
rect 502885 453794 502951 453797
rect 499836 453792 502951 453794
rect 499836 453736 502890 453792
rect 502946 453736 502951 453792
rect 499836 453734 502951 453736
rect 502885 453731 502951 453734
rect 58750 453460 58756 453524
rect 58820 453522 58826 453524
rect 536782 453522 536788 453524
rect 58820 453462 60076 453522
rect 499836 453462 536788 453522
rect 58820 453460 58826 453462
rect 536782 453460 536788 453462
rect 536852 453460 536858 453524
rect 502793 453250 502859 453253
rect 499836 453248 502859 453250
rect 499836 453192 502798 453248
rect 502854 453192 502859 453248
rect 499836 453190 502859 453192
rect 502793 453187 502859 453190
rect 54334 452916 54340 452980
rect 54404 452978 54410 452980
rect 503989 452978 504055 452981
rect 54404 452918 60076 452978
rect 499836 452976 504055 452978
rect 499836 452920 503994 452976
rect 504050 452920 504055 452976
rect 499836 452918 504055 452920
rect 54404 452916 54410 452918
rect 503989 452915 504055 452918
rect 502701 452706 502767 452709
rect 499836 452704 502767 452706
rect 499836 452648 502706 452704
rect 502762 452648 502767 452704
rect 499836 452646 502767 452648
rect 502701 452643 502767 452646
rect 25998 452372 26004 452436
rect 26068 452434 26074 452436
rect 502885 452434 502951 452437
rect 26068 452374 60076 452434
rect 499836 452432 502951 452434
rect 499836 452376 502890 452432
rect 502946 452376 502951 452432
rect 499836 452374 502951 452376
rect 26068 452372 26074 452374
rect 502885 452371 502951 452374
rect 502701 452162 502767 452165
rect 499836 452160 502767 452162
rect 499836 452104 502706 452160
rect 502762 452104 502767 452160
rect 499836 452102 502767 452104
rect 502701 452099 502767 452102
rect 28758 451828 28764 451892
rect 28828 451890 28834 451892
rect 502793 451890 502859 451893
rect 28828 451830 60076 451890
rect 499836 451888 502859 451890
rect 499836 451832 502798 451888
rect 502854 451832 502859 451888
rect 499836 451830 502859 451832
rect 28828 451828 28834 451830
rect 502793 451827 502859 451830
rect 502609 451618 502675 451621
rect 499836 451616 502675 451618
rect 499836 451560 502614 451616
rect 502670 451560 502675 451616
rect 499836 451558 502675 451560
rect 502609 451555 502675 451558
rect 48078 451284 48084 451348
rect 48148 451346 48154 451348
rect 500125 451346 500191 451349
rect 48148 451286 60076 451346
rect 499836 451344 500191 451346
rect 499836 451288 500130 451344
rect 500186 451288 500191 451344
rect 499836 451286 500191 451288
rect 48148 451284 48154 451286
rect 500125 451283 500191 451286
rect 500861 451210 500927 451213
rect 503621 451210 503687 451213
rect 500861 451208 503687 451210
rect 500861 451152 500866 451208
rect 500922 451152 503626 451208
rect 503682 451152 503687 451208
rect 500861 451150 503687 451152
rect 500861 451147 500927 451150
rect 503621 451147 503687 451150
rect 503621 451074 503687 451077
rect 499836 451072 503687 451074
rect 499836 451016 503626 451072
rect 503682 451016 503687 451072
rect 499836 451014 503687 451016
rect 503621 451011 503687 451014
rect 31518 450740 31524 450804
rect 31588 450802 31594 450804
rect 503621 450802 503687 450805
rect 31588 450742 60076 450802
rect 499836 450800 503687 450802
rect 499836 450744 503626 450800
rect 503682 450744 503687 450800
rect 499836 450742 503687 450744
rect 31588 450740 31594 450742
rect 503621 450739 503687 450742
rect 502701 450530 502767 450533
rect 499836 450528 502767 450530
rect 499836 450472 502706 450528
rect 502762 450472 502767 450528
rect 499836 450470 502767 450472
rect 502701 450467 502767 450470
rect 34278 450196 34284 450260
rect 34348 450258 34354 450260
rect 502885 450258 502951 450261
rect 34348 450198 60076 450258
rect 499836 450256 502951 450258
rect 499836 450200 502890 450256
rect 502946 450200 502951 450256
rect 499836 450198 502951 450200
rect 34348 450196 34354 450198
rect 502885 450195 502951 450198
rect 502609 449986 502675 449989
rect 499836 449984 502675 449986
rect 499836 449928 502614 449984
rect 502670 449928 502675 449984
rect 499836 449926 502675 449928
rect 502609 449923 502675 449926
rect -960 449578 480 449668
rect 54702 449652 54708 449716
rect 54772 449714 54778 449716
rect 503621 449714 503687 449717
rect 54772 449654 60076 449714
rect 499836 449712 503687 449714
rect 499836 449656 503626 449712
rect 503682 449656 503687 449712
rect 499836 449654 503687 449656
rect 54772 449652 54778 449654
rect 503621 449651 503687 449654
rect 3734 449578 3740 449580
rect -960 449518 3740 449578
rect -960 449428 480 449518
rect 3734 449516 3740 449518
rect 3804 449516 3810 449580
rect 503621 449442 503687 449445
rect 499836 449440 503687 449442
rect 499836 449384 503626 449440
rect 503682 449384 503687 449440
rect 499836 449382 503687 449384
rect 503621 449379 503687 449382
rect 32990 449108 32996 449172
rect 33060 449170 33066 449172
rect 502885 449170 502951 449173
rect 33060 449110 60076 449170
rect 499836 449168 502951 449170
rect 499836 449112 502890 449168
rect 502946 449112 502951 449168
rect 499836 449110 502951 449112
rect 33060 449108 33066 449110
rect 502885 449107 502951 449110
rect 502701 448898 502767 448901
rect 499836 448896 502767 448898
rect 499836 448840 502706 448896
rect 502762 448840 502767 448896
rect 499836 448838 502767 448840
rect 502701 448835 502767 448838
rect 57278 448564 57284 448628
rect 57348 448626 57354 448628
rect 502793 448626 502859 448629
rect 57348 448566 60076 448626
rect 499836 448624 502859 448626
rect 499836 448568 502798 448624
rect 502854 448568 502859 448624
rect 499836 448566 502859 448568
rect 57348 448564 57354 448566
rect 502793 448563 502859 448566
rect 503621 448354 503687 448357
rect 499836 448352 503687 448354
rect 499836 448296 503626 448352
rect 503682 448296 503687 448352
rect 499836 448294 503687 448296
rect 503621 448291 503687 448294
rect 31334 448020 31340 448084
rect 31404 448082 31410 448084
rect 502885 448082 502951 448085
rect 31404 448022 60076 448082
rect 499836 448080 502951 448082
rect 499836 448024 502890 448080
rect 502946 448024 502951 448080
rect 499836 448022 502951 448024
rect 31404 448020 31410 448022
rect 502885 448019 502951 448022
rect 502701 447810 502767 447813
rect 499836 447808 502767 447810
rect 499836 447752 502706 447808
rect 502762 447752 502767 447808
rect 499836 447750 502767 447752
rect 502701 447747 502767 447750
rect 53598 447476 53604 447540
rect 53668 447538 53674 447540
rect 502609 447538 502675 447541
rect 53668 447478 60076 447538
rect 499836 447536 502675 447538
rect 499836 447480 502614 447536
rect 502670 447480 502675 447536
rect 499836 447478 502675 447480
rect 53668 447476 53674 447478
rect 502609 447475 502675 447478
rect 508405 447266 508471 447269
rect 499836 447264 508471 447266
rect 499836 447208 508410 447264
rect 508466 447208 508471 447264
rect 499836 447206 508471 447208
rect 508405 447203 508471 447206
rect 59118 446932 59124 446996
rect 59188 446994 59194 446996
rect 512545 446994 512611 446997
rect 59188 446934 60076 446994
rect 499836 446992 512611 446994
rect 499836 446936 512550 446992
rect 512606 446936 512611 446992
rect 499836 446934 512611 446936
rect 59188 446932 59194 446934
rect 512545 446931 512611 446934
rect 512269 446722 512335 446725
rect 499836 446720 512335 446722
rect 499836 446664 512274 446720
rect 512330 446664 512335 446720
rect 499836 446662 512335 446664
rect 512269 446659 512335 446662
rect 58382 446388 58388 446452
rect 58452 446450 58458 446452
rect 512729 446450 512795 446453
rect 58452 446390 60076 446450
rect 499836 446448 512795 446450
rect 499836 446392 512734 446448
rect 512790 446392 512795 446448
rect 499836 446390 512795 446392
rect 58452 446388 58458 446390
rect 512729 446387 512795 446390
rect 519537 446178 519603 446181
rect 499836 446176 519603 446178
rect 499836 446120 519542 446176
rect 519598 446120 519603 446176
rect 499836 446118 519603 446120
rect 519537 446115 519603 446118
rect 59854 445844 59860 445908
rect 59924 445906 59930 445908
rect 507117 445906 507183 445909
rect 59924 445846 60076 445906
rect 499836 445904 507183 445906
rect 499836 445848 507122 445904
rect 507178 445848 507183 445904
rect 499836 445846 507183 445848
rect 59924 445844 59930 445846
rect 507117 445843 507183 445846
rect 512453 445634 512519 445637
rect 499836 445632 512519 445634
rect 499836 445576 512458 445632
rect 512514 445576 512519 445632
rect 499836 445574 512519 445576
rect 512453 445571 512519 445574
rect 52310 445300 52316 445364
rect 52380 445362 52386 445364
rect 503621 445362 503687 445365
rect 52380 445302 60076 445362
rect 499836 445360 503687 445362
rect 499836 445304 503626 445360
rect 503682 445304 503687 445360
rect 499836 445302 503687 445304
rect 52380 445300 52386 445302
rect 503621 445299 503687 445302
rect 507025 445090 507091 445093
rect 499836 445088 507091 445090
rect 499836 445032 507030 445088
rect 507086 445032 507091 445088
rect 499836 445030 507091 445032
rect 507025 445027 507091 445030
rect 41086 444756 41092 444820
rect 41156 444818 41162 444820
rect 534993 444818 535059 444821
rect 41156 444758 60076 444818
rect 499836 444816 535059 444818
rect 499836 444760 534998 444816
rect 535054 444760 535059 444816
rect 499836 444758 535059 444760
rect 41156 444756 41162 444758
rect 534993 444755 535059 444758
rect 583520 444668 584960 444908
rect 500125 444546 500191 444549
rect 499836 444544 500191 444546
rect 499836 444488 500130 444544
rect 500186 444488 500191 444544
rect 499836 444486 500191 444488
rect 500125 444483 500191 444486
rect 57830 444212 57836 444276
rect 57900 444274 57906 444276
rect 519445 444274 519511 444277
rect 57900 444214 60076 444274
rect 499836 444272 519511 444274
rect 499836 444216 519450 444272
rect 519506 444216 519511 444272
rect 499836 444214 519511 444216
rect 57900 444212 57906 444214
rect 519445 444211 519511 444214
rect 504173 444002 504239 444005
rect 499836 444000 504239 444002
rect 499836 443944 504178 444000
rect 504234 443944 504239 444000
rect 499836 443942 504239 443944
rect 504173 443939 504239 443942
rect 39614 443668 39620 443732
rect 39684 443730 39690 443732
rect 501505 443730 501571 443733
rect 39684 443670 60076 443730
rect 499836 443728 501571 443730
rect 499836 443672 501510 443728
rect 501566 443672 501571 443728
rect 499836 443670 501571 443672
rect 39684 443668 39690 443670
rect 501505 443667 501571 443670
rect 500125 443458 500191 443461
rect 499836 443456 500191 443458
rect 499836 443400 500130 443456
rect 500186 443400 500191 443456
rect 499836 443398 500191 443400
rect 500125 443395 500191 443398
rect 44766 443124 44772 443188
rect 44836 443186 44842 443188
rect 501321 443186 501387 443189
rect 44836 443126 60076 443186
rect 499836 443184 501387 443186
rect 499836 443128 501326 443184
rect 501382 443128 501387 443184
rect 499836 443126 501387 443128
rect 44836 443124 44842 443126
rect 501321 443123 501387 443126
rect 501137 442914 501203 442917
rect 499836 442912 501203 442914
rect 499836 442856 501142 442912
rect 501198 442856 501203 442912
rect 499836 442854 501203 442856
rect 501137 442851 501203 442854
rect 37406 442580 37412 442644
rect 37476 442642 37482 442644
rect 502057 442642 502123 442645
rect 37476 442582 60076 442642
rect 499836 442640 502123 442642
rect 499836 442584 502062 442640
rect 502118 442584 502123 442640
rect 499836 442582 502123 442584
rect 37476 442580 37482 442582
rect 502057 442579 502123 442582
rect 500125 442370 500191 442373
rect 499836 442368 500191 442370
rect 499836 442312 500130 442368
rect 500186 442312 500191 442368
rect 499836 442310 500191 442312
rect 500125 442307 500191 442310
rect 37038 442036 37044 442100
rect 37108 442098 37114 442100
rect 500217 442098 500283 442101
rect 37108 442038 60076 442098
rect 499836 442096 500283 442098
rect 499836 442040 500222 442096
rect 500278 442040 500283 442096
rect 499836 442038 500283 442040
rect 37108 442036 37114 442038
rect 500217 442035 500283 442038
rect 503621 441826 503687 441829
rect 499836 441824 503687 441826
rect 499836 441768 503626 441824
rect 503682 441768 503687 441824
rect 499836 441766 503687 441768
rect 503621 441763 503687 441766
rect 32806 441492 32812 441556
rect 32876 441554 32882 441556
rect 501229 441554 501295 441557
rect 32876 441494 60076 441554
rect 499836 441552 501295 441554
rect 499836 441496 501234 441552
rect 501290 441496 501295 441552
rect 499836 441494 501295 441496
rect 32876 441492 32882 441494
rect 501229 441491 501295 441494
rect 510981 441282 511047 441285
rect 499836 441280 511047 441282
rect 499836 441224 510986 441280
rect 511042 441224 511047 441280
rect 499836 441222 511047 441224
rect 510981 441219 511047 441222
rect 34094 440948 34100 441012
rect 34164 441010 34170 441012
rect 509601 441010 509667 441013
rect 34164 440950 60076 441010
rect 499836 441008 509667 441010
rect 499836 440952 509606 441008
rect 509662 440952 509667 441008
rect 499836 440950 509667 440952
rect 34164 440948 34170 440950
rect 509601 440947 509667 440950
rect 503621 440738 503687 440741
rect 499836 440736 503687 440738
rect 499836 440680 503626 440736
rect 503682 440680 503687 440736
rect 499836 440678 503687 440680
rect 503621 440675 503687 440678
rect 32622 440404 32628 440468
rect 32692 440466 32698 440468
rect 510889 440466 510955 440469
rect 32692 440406 60076 440466
rect 499836 440464 510955 440466
rect 499836 440408 510894 440464
rect 510950 440408 510955 440464
rect 499836 440406 510955 440408
rect 32692 440404 32698 440406
rect 510889 440403 510955 440406
rect 503621 440194 503687 440197
rect 499836 440192 503687 440194
rect 499836 440136 503626 440192
rect 503682 440136 503687 440192
rect 499836 440134 503687 440136
rect 503621 440131 503687 440134
rect 47526 439860 47532 439924
rect 47596 439922 47602 439924
rect 503621 439922 503687 439925
rect 47596 439862 60076 439922
rect 499836 439920 503687 439922
rect 499836 439864 503626 439920
rect 503682 439864 503687 439920
rect 499836 439862 503687 439864
rect 47596 439860 47602 439862
rect 503621 439859 503687 439862
rect 522021 439650 522087 439653
rect 499836 439648 522087 439650
rect 499836 439592 522026 439648
rect 522082 439592 522087 439648
rect 499836 439590 522087 439592
rect 522021 439587 522087 439590
rect 46606 439316 46612 439380
rect 46676 439378 46682 439380
rect 512085 439378 512151 439381
rect 46676 439318 60076 439378
rect 499836 439376 512151 439378
rect 499836 439320 512090 439376
rect 512146 439320 512151 439376
rect 499836 439318 512151 439320
rect 46676 439316 46682 439318
rect 512085 439315 512151 439318
rect 504081 439106 504147 439109
rect 499836 439104 504147 439106
rect 499836 439048 504086 439104
rect 504142 439048 504147 439104
rect 499836 439046 504147 439048
rect 504081 439043 504147 439046
rect 44950 438772 44956 438836
rect 45020 438834 45026 438836
rect 501045 438834 501111 438837
rect 45020 438774 60076 438834
rect 499836 438832 501111 438834
rect 499836 438776 501050 438832
rect 501106 438776 501111 438832
rect 499836 438774 501111 438776
rect 45020 438772 45026 438774
rect 501045 438771 501111 438774
rect 504265 438562 504331 438565
rect 499836 438560 504331 438562
rect 499836 438504 504270 438560
rect 504326 438504 504331 438560
rect 499836 438502 504331 438504
rect 504265 438499 504331 438502
rect 49049 438290 49115 438293
rect 504357 438290 504423 438293
rect 49049 438288 60076 438290
rect 49049 438232 49054 438288
rect 49110 438232 60076 438288
rect 49049 438230 60076 438232
rect 499836 438288 504423 438290
rect 499836 438232 504362 438288
rect 504418 438232 504423 438288
rect 499836 438230 504423 438232
rect 49049 438227 49115 438230
rect 504357 438227 504423 438230
rect 503621 438018 503687 438021
rect 499836 438016 503687 438018
rect 499836 437960 503626 438016
rect 503682 437960 503687 438016
rect 499836 437958 503687 437960
rect 503621 437955 503687 437958
rect 57513 437746 57579 437749
rect 503529 437746 503595 437749
rect 57513 437744 60076 437746
rect 57513 437688 57518 437744
rect 57574 437688 60076 437744
rect 57513 437686 60076 437688
rect 499836 437744 503595 437746
rect 499836 437688 503534 437744
rect 503590 437688 503595 437744
rect 499836 437686 503595 437688
rect 57513 437683 57579 437686
rect 503529 437683 503595 437686
rect 512361 437474 512427 437477
rect 499836 437472 512427 437474
rect 499836 437416 512366 437472
rect 512422 437416 512427 437472
rect 499836 437414 512427 437416
rect 512361 437411 512427 437414
rect 49141 437202 49207 437205
rect 503621 437202 503687 437205
rect 49141 437200 60076 437202
rect 49141 437144 49146 437200
rect 49202 437144 60076 437200
rect 49141 437142 60076 437144
rect 499836 437200 503687 437202
rect 499836 437144 503626 437200
rect 503682 437144 503687 437200
rect 499836 437142 503687 437144
rect 49141 437139 49207 437142
rect 503621 437139 503687 437142
rect 503621 436930 503687 436933
rect 499836 436928 503687 436930
rect 499836 436872 503626 436928
rect 503682 436872 503687 436928
rect 499836 436870 503687 436872
rect 503621 436867 503687 436870
rect -960 436508 480 436748
rect 48957 436658 49023 436661
rect 523585 436658 523651 436661
rect 48957 436656 60076 436658
rect 48957 436600 48962 436656
rect 49018 436600 60076 436656
rect 48957 436598 60076 436600
rect 499836 436656 523651 436658
rect 499836 436600 523590 436656
rect 523646 436600 523651 436656
rect 499836 436598 523651 436600
rect 48957 436595 49023 436598
rect 523585 436595 523651 436598
rect 524781 436386 524847 436389
rect 499836 436384 524847 436386
rect 499836 436328 524786 436384
rect 524842 436328 524847 436384
rect 499836 436326 524847 436328
rect 524781 436323 524847 436326
rect 49417 436114 49483 436117
rect 525190 436114 525196 436116
rect 49417 436112 60076 436114
rect 49417 436056 49422 436112
rect 49478 436056 60076 436112
rect 49417 436054 60076 436056
rect 499836 436054 525196 436114
rect 49417 436051 49483 436054
rect 525190 436052 525196 436054
rect 525260 436052 525266 436116
rect 520825 435842 520891 435845
rect 499836 435840 520891 435842
rect 499836 435784 520830 435840
rect 520886 435784 520891 435840
rect 499836 435782 520891 435784
rect 520825 435779 520891 435782
rect 50245 435570 50311 435573
rect 503621 435570 503687 435573
rect 50245 435568 60076 435570
rect 50245 435512 50250 435568
rect 50306 435512 60076 435568
rect 50245 435510 60076 435512
rect 499836 435568 503687 435570
rect 499836 435512 503626 435568
rect 503682 435512 503687 435568
rect 499836 435510 503687 435512
rect 50245 435507 50311 435510
rect 503621 435507 503687 435510
rect 519118 435298 519124 435300
rect 499836 435238 519124 435298
rect 519118 435236 519124 435238
rect 519188 435236 519194 435300
rect 42057 435026 42123 435029
rect 520222 435026 520228 435028
rect 42057 435024 60076 435026
rect 42057 434968 42062 435024
rect 42118 434968 60076 435024
rect 42057 434966 60076 434968
rect 499836 434966 520228 435026
rect 42057 434963 42123 434966
rect 520222 434964 520228 434966
rect 520292 434964 520298 435028
rect 503437 434754 503503 434757
rect 499836 434752 503503 434754
rect 499836 434696 503442 434752
rect 503498 434696 503503 434752
rect 499836 434694 503503 434696
rect 503437 434691 503503 434694
rect 51625 434482 51691 434485
rect 503621 434482 503687 434485
rect 51625 434480 60076 434482
rect 51625 434424 51630 434480
rect 51686 434424 60076 434480
rect 51625 434422 60076 434424
rect 499836 434480 503687 434482
rect 499836 434424 503626 434480
rect 503682 434424 503687 434480
rect 499836 434422 503687 434424
rect 51625 434419 51691 434422
rect 503621 434419 503687 434422
rect 502793 434210 502859 434213
rect 499836 434208 502859 434210
rect 499836 434152 502798 434208
rect 502854 434152 502859 434208
rect 499836 434150 502859 434152
rect 502793 434147 502859 434150
rect 51533 433938 51599 433941
rect 503529 433938 503595 433941
rect 51533 433936 60076 433938
rect 51533 433880 51538 433936
rect 51594 433880 60076 433936
rect 51533 433878 60076 433880
rect 499836 433936 503595 433938
rect 499836 433880 503534 433936
rect 503590 433880 503595 433936
rect 499836 433878 503595 433880
rect 51533 433875 51599 433878
rect 503529 433875 503595 433878
rect 503897 433666 503963 433669
rect 499836 433664 503963 433666
rect 499836 433608 503902 433664
rect 503958 433608 503963 433664
rect 499836 433606 503963 433608
rect 503897 433603 503963 433606
rect 49325 433394 49391 433397
rect 503437 433394 503503 433397
rect 49325 433392 60076 433394
rect 49325 433336 49330 433392
rect 49386 433336 60076 433392
rect 49325 433334 60076 433336
rect 499836 433392 503503 433394
rect 499836 433336 503442 433392
rect 503498 433336 503503 433392
rect 499836 433334 503503 433336
rect 49325 433331 49391 433334
rect 503437 433331 503503 433334
rect 503437 433122 503503 433125
rect 499836 433120 503503 433122
rect 499836 433064 503442 433120
rect 503498 433064 503503 433120
rect 499836 433062 503503 433064
rect 503437 433059 503503 433062
rect 49233 432850 49299 432853
rect 502609 432850 502675 432853
rect 49233 432848 60076 432850
rect 49233 432792 49238 432848
rect 49294 432792 60076 432848
rect 49233 432790 60076 432792
rect 499836 432848 502675 432850
rect 499836 432792 502614 432848
rect 502670 432792 502675 432848
rect 499836 432790 502675 432792
rect 49233 432787 49299 432790
rect 502609 432787 502675 432790
rect 503529 432578 503595 432581
rect 499836 432576 503595 432578
rect 499836 432520 503534 432576
rect 503590 432520 503595 432576
rect 499836 432518 503595 432520
rect 503529 432515 503595 432518
rect 25497 432306 25563 432309
rect 503621 432306 503687 432309
rect 25497 432304 60076 432306
rect 25497 432248 25502 432304
rect 25558 432248 60076 432304
rect 25497 432246 60076 432248
rect 499836 432304 503687 432306
rect 499836 432248 503626 432304
rect 503682 432248 503687 432304
rect 499836 432246 503687 432248
rect 25497 432243 25563 432246
rect 503621 432243 503687 432246
rect 503437 432034 503503 432037
rect 499836 432032 503503 432034
rect 499836 431976 503442 432032
rect 503498 431976 503503 432032
rect 499836 431974 503503 431976
rect 503437 431971 503503 431974
rect 39481 431762 39547 431765
rect 503621 431762 503687 431765
rect 39481 431760 60076 431762
rect 39481 431704 39486 431760
rect 39542 431704 60076 431760
rect 39481 431702 60076 431704
rect 499836 431760 503687 431762
rect 499836 431704 503626 431760
rect 503682 431704 503687 431760
rect 499836 431702 503687 431704
rect 39481 431699 39547 431702
rect 503621 431699 503687 431702
rect 580441 431626 580507 431629
rect 583520 431626 584960 431716
rect 580441 431624 584960 431626
rect 580441 431568 580446 431624
rect 580502 431568 584960 431624
rect 580441 431566 584960 431568
rect 580441 431563 580507 431566
rect 503529 431490 503595 431493
rect 499836 431488 503595 431490
rect 499836 431432 503534 431488
rect 503590 431432 503595 431488
rect 583520 431476 584960 431566
rect 499836 431430 503595 431432
rect 503529 431427 503595 431430
rect 55673 431218 55739 431221
rect 503437 431218 503503 431221
rect 55673 431216 60076 431218
rect 55673 431160 55678 431216
rect 55734 431160 60076 431216
rect 55673 431158 60076 431160
rect 499836 431216 503503 431218
rect 499836 431160 503442 431216
rect 503498 431160 503503 431216
rect 499836 431158 503503 431160
rect 55673 431155 55739 431158
rect 503437 431155 503503 431158
rect 502517 430946 502583 430949
rect 499836 430944 502583 430946
rect 499836 430888 502522 430944
rect 502578 430888 502583 430944
rect 499836 430886 502583 430888
rect 502517 430883 502583 430886
rect 50337 430674 50403 430677
rect 502701 430674 502767 430677
rect 50337 430672 60076 430674
rect 50337 430616 50342 430672
rect 50398 430616 60076 430672
rect 50337 430614 60076 430616
rect 499836 430672 502767 430674
rect 499836 430616 502706 430672
rect 502762 430616 502767 430672
rect 499836 430614 502767 430616
rect 50337 430611 50403 430614
rect 502701 430611 502767 430614
rect 503621 430402 503687 430405
rect 499836 430400 503687 430402
rect 499836 430344 503626 430400
rect 503682 430344 503687 430400
rect 499836 430342 503687 430344
rect 503621 430339 503687 430342
rect 58985 430130 59051 430133
rect 502609 430130 502675 430133
rect 58985 430128 60076 430130
rect 58985 430072 58990 430128
rect 59046 430072 60076 430128
rect 58985 430070 60076 430072
rect 499836 430128 502675 430130
rect 499836 430072 502614 430128
rect 502670 430072 502675 430128
rect 499836 430070 502675 430072
rect 58985 430067 59051 430070
rect 502609 430067 502675 430070
rect 503621 429992 503687 429997
rect 503621 429936 503626 429992
rect 503682 429936 503687 429992
rect 503621 429931 503687 429936
rect 503624 429858 503684 429931
rect 499836 429798 503684 429858
rect 36629 429586 36695 429589
rect 503529 429586 503595 429589
rect 36629 429584 60076 429586
rect 36629 429528 36634 429584
rect 36690 429528 60076 429584
rect 36629 429526 60076 429528
rect 499836 429584 503595 429586
rect 499836 429528 503534 429584
rect 503590 429528 503595 429584
rect 499836 429526 503595 429528
rect 36629 429523 36695 429526
rect 503529 429523 503595 429526
rect 503437 429314 503503 429317
rect 499836 429312 503503 429314
rect 499836 429256 503442 429312
rect 503498 429256 503503 429312
rect 499836 429254 503503 429256
rect 503437 429251 503503 429254
rect 58893 429042 58959 429045
rect 503621 429042 503687 429045
rect 58893 429040 60076 429042
rect 58893 428984 58898 429040
rect 58954 428984 60076 429040
rect 58893 428982 60076 428984
rect 499836 429040 503687 429042
rect 499836 428984 503626 429040
rect 503682 428984 503687 429040
rect 499836 428982 503687 428984
rect 58893 428979 58959 428982
rect 503621 428979 503687 428982
rect 503621 428770 503687 428773
rect 499836 428768 503687 428770
rect 499836 428712 503626 428768
rect 503682 428712 503687 428768
rect 499836 428710 503687 428712
rect 503621 428707 503687 428710
rect 57145 428498 57211 428501
rect 503621 428498 503687 428501
rect 57145 428496 60076 428498
rect 57145 428440 57150 428496
rect 57206 428440 60076 428496
rect 57145 428438 60076 428440
rect 499836 428496 503687 428498
rect 499836 428440 503626 428496
rect 503682 428440 503687 428496
rect 499836 428438 503687 428440
rect 57145 428435 57211 428438
rect 503621 428435 503687 428438
rect 502517 428226 502583 428229
rect 499836 428224 502583 428226
rect 499836 428168 502522 428224
rect 502578 428168 502583 428224
rect 499836 428166 502583 428168
rect 502517 428163 502583 428166
rect 59077 427954 59143 427957
rect 503621 427954 503687 427957
rect 59077 427952 60076 427954
rect 59077 427896 59082 427952
rect 59138 427896 60076 427952
rect 59077 427894 60076 427896
rect 499836 427952 503687 427954
rect 499836 427896 503626 427952
rect 503682 427896 503687 427952
rect 499836 427894 503687 427896
rect 59077 427891 59143 427894
rect 503621 427891 503687 427894
rect 502701 427682 502767 427685
rect 499836 427680 502767 427682
rect 499836 427624 502706 427680
rect 502762 427624 502767 427680
rect 499836 427622 502767 427624
rect 502701 427619 502767 427622
rect 32489 427410 32555 427413
rect 502793 427410 502859 427413
rect 32489 427408 60076 427410
rect 32489 427352 32494 427408
rect 32550 427352 60076 427408
rect 32489 427350 60076 427352
rect 499836 427408 502859 427410
rect 499836 427352 502798 427408
rect 502854 427352 502859 427408
rect 499836 427350 502859 427352
rect 32489 427347 32555 427350
rect 502793 427347 502859 427350
rect 503621 427138 503687 427141
rect 499836 427136 503687 427138
rect 499836 427080 503626 427136
rect 503682 427080 503687 427136
rect 499836 427078 503687 427080
rect 503621 427075 503687 427078
rect 533337 427138 533403 427141
rect 536373 427138 536439 427141
rect 533337 427136 536439 427138
rect 533337 427080 533342 427136
rect 533398 427080 536378 427136
rect 536434 427080 536439 427136
rect 533337 427078 536439 427080
rect 533337 427075 533403 427078
rect 536373 427075 536439 427078
rect 35249 426866 35315 426869
rect 503437 426866 503503 426869
rect 35249 426864 60076 426866
rect 35249 426808 35254 426864
rect 35310 426808 60076 426864
rect 35249 426806 60076 426808
rect 499836 426864 503503 426866
rect 499836 426808 503442 426864
rect 503498 426808 503503 426864
rect 499836 426806 503503 426808
rect 35249 426803 35315 426806
rect 503437 426803 503503 426806
rect 503529 426594 503595 426597
rect 499836 426592 503595 426594
rect 499836 426536 503534 426592
rect 503590 426536 503595 426592
rect 499836 426534 503595 426536
rect 503529 426531 503595 426534
rect 50153 426322 50219 426325
rect 503621 426322 503687 426325
rect 50153 426320 60076 426322
rect 50153 426264 50158 426320
rect 50214 426264 60076 426320
rect 50153 426262 60076 426264
rect 499836 426320 503687 426322
rect 499836 426264 503626 426320
rect 503682 426264 503687 426320
rect 499836 426262 503687 426264
rect 50153 426259 50219 426262
rect 503621 426259 503687 426262
rect 515673 426050 515739 426053
rect 499836 426048 515739 426050
rect 499836 425992 515678 426048
rect 515734 425992 515739 426048
rect 499836 425990 515739 425992
rect 515673 425987 515739 425990
rect 47669 425778 47735 425781
rect 503437 425778 503503 425781
rect 47669 425776 60076 425778
rect 47669 425720 47674 425776
rect 47730 425720 60076 425776
rect 47669 425718 60076 425720
rect 499836 425776 503503 425778
rect 499836 425720 503442 425776
rect 503498 425720 503503 425776
rect 499836 425718 503503 425720
rect 47669 425715 47735 425718
rect 503437 425715 503503 425718
rect 502885 425506 502951 425509
rect 499836 425504 502951 425506
rect 499836 425448 502890 425504
rect 502946 425448 502951 425504
rect 499836 425446 502951 425448
rect 502885 425443 502951 425446
rect 53189 425234 53255 425237
rect 503529 425234 503595 425237
rect 53189 425232 60076 425234
rect 53189 425176 53194 425232
rect 53250 425176 60076 425232
rect 53189 425174 60076 425176
rect 499836 425232 503595 425234
rect 499836 425176 503534 425232
rect 503590 425176 503595 425232
rect 499836 425174 503595 425176
rect 53189 425171 53255 425174
rect 503529 425171 503595 425174
rect 503621 424962 503687 424965
rect 499836 424960 503687 424962
rect 499836 424904 503626 424960
rect 503682 424904 503687 424960
rect 499836 424902 503687 424904
rect 503621 424899 503687 424902
rect 47761 424690 47827 424693
rect 517881 424690 517947 424693
rect 47761 424688 60076 424690
rect 47761 424632 47766 424688
rect 47822 424632 60076 424688
rect 47761 424630 60076 424632
rect 499836 424688 517947 424690
rect 499836 424632 517886 424688
rect 517942 424632 517947 424688
rect 499836 424630 517947 424632
rect 47761 424627 47827 424630
rect 517881 424627 517947 424630
rect 503621 424418 503687 424421
rect 499836 424416 503687 424418
rect 499836 424360 503626 424416
rect 503682 424360 503687 424416
rect 499836 424358 503687 424360
rect 503621 424355 503687 424358
rect 50429 424146 50495 424149
rect 503529 424146 503595 424149
rect 50429 424144 60076 424146
rect 50429 424088 50434 424144
rect 50490 424088 60076 424144
rect 50429 424086 60076 424088
rect 499836 424144 503595 424146
rect 499836 424088 503534 424144
rect 503590 424088 503595 424144
rect 499836 424086 503595 424088
rect 50429 424083 50495 424086
rect 503529 424083 503595 424086
rect 503437 423874 503503 423877
rect 499836 423872 503503 423874
rect 499836 423816 503442 423872
rect 503498 423816 503503 423872
rect 499836 423814 503503 423816
rect 503437 423811 503503 423814
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 59169 423602 59235 423605
rect 503621 423602 503687 423605
rect 59169 423600 60076 423602
rect 59169 423544 59174 423600
rect 59230 423544 60076 423600
rect 59169 423542 60076 423544
rect 499836 423600 503687 423602
rect 499836 423544 503626 423600
rect 503682 423544 503687 423600
rect 499836 423542 503687 423544
rect 59169 423539 59235 423542
rect 503621 423539 503687 423542
rect 502609 423330 502675 423333
rect 499836 423328 502675 423330
rect 499836 423272 502614 423328
rect 502670 423272 502675 423328
rect 499836 423270 502675 423272
rect 502609 423267 502675 423270
rect 32673 423058 32739 423061
rect 502425 423058 502491 423061
rect 32673 423056 60076 423058
rect 32673 423000 32678 423056
rect 32734 423000 60076 423056
rect 32673 422998 60076 423000
rect 499836 423056 502491 423058
rect 499836 423000 502430 423056
rect 502486 423000 502491 423056
rect 499836 422998 502491 423000
rect 32673 422995 32739 422998
rect 502425 422995 502491 422998
rect 502517 422786 502583 422789
rect 499836 422784 502583 422786
rect 499836 422728 502522 422784
rect 502578 422728 502583 422784
rect 499836 422726 502583 422728
rect 502517 422723 502583 422726
rect 50521 422514 50587 422517
rect 502701 422514 502767 422517
rect 50521 422512 60076 422514
rect 50521 422456 50526 422512
rect 50582 422456 60076 422512
rect 50521 422454 60076 422456
rect 499836 422512 502767 422514
rect 499836 422456 502706 422512
rect 502762 422456 502767 422512
rect 499836 422454 502767 422456
rect 50521 422451 50587 422454
rect 502701 422451 502767 422454
rect 32581 421970 32647 421973
rect 32581 421968 60076 421970
rect 32581 421912 32586 421968
rect 32642 421912 60076 421968
rect 32581 421910 60076 421912
rect 32581 421907 32647 421910
rect 35157 421426 35223 421429
rect 35157 421424 60076 421426
rect 35157 421368 35162 421424
rect 35218 421368 60076 421424
rect 35157 421366 60076 421368
rect 35157 421363 35223 421366
rect 26969 420882 27035 420885
rect 26969 420880 60076 420882
rect 26969 420824 26974 420880
rect 27030 420824 60076 420880
rect 26969 420822 60076 420824
rect 26969 420819 27035 420822
rect 31201 420338 31267 420341
rect 31201 420336 60076 420338
rect 31201 420280 31206 420336
rect 31262 420280 60076 420336
rect 31201 420278 60076 420280
rect 31201 420275 31267 420278
rect 41965 419794 42031 419797
rect 41965 419792 60076 419794
rect 41965 419736 41970 419792
rect 42026 419736 60076 419792
rect 41965 419734 60076 419736
rect 41965 419731 42031 419734
rect 40493 419250 40559 419253
rect 40493 419248 60076 419250
rect 40493 419192 40498 419248
rect 40554 419192 60076 419248
rect 40493 419190 60076 419192
rect 40493 419187 40559 419190
rect 46381 418706 46447 418709
rect 46381 418704 60076 418706
rect 46381 418648 46386 418704
rect 46442 418648 60076 418704
rect 46381 418646 60076 418648
rect 46381 418643 46447 418646
rect 544326 418236 544332 418300
rect 544396 418298 544402 418300
rect 583520 418298 584960 418388
rect 544396 418238 584960 418298
rect 544396 418236 544402 418238
rect 46289 418162 46355 418165
rect 46289 418160 60076 418162
rect 46289 418104 46294 418160
rect 46350 418104 60076 418160
rect 583520 418148 584960 418238
rect 46289 418102 60076 418104
rect 46289 418099 46355 418102
rect 51717 417618 51783 417621
rect 51717 417616 60076 417618
rect 51717 417560 51722 417616
rect 51778 417560 60076 417616
rect 51717 417558 60076 417560
rect 51717 417555 51783 417558
rect 41270 417012 41276 417076
rect 41340 417074 41346 417076
rect 41340 417014 60076 417074
rect 41340 417012 41346 417014
rect 39246 416468 39252 416532
rect 39316 416530 39322 416532
rect 39316 416470 60076 416530
rect 39316 416468 39322 416470
rect 39062 415924 39068 415988
rect 39132 415986 39138 415988
rect 39132 415926 60076 415986
rect 39132 415924 39138 415926
rect 42374 415380 42380 415444
rect 42444 415442 42450 415444
rect 42444 415382 60076 415442
rect 42444 415380 42450 415382
rect 30230 414836 30236 414900
rect 30300 414898 30306 414900
rect 30300 414838 60076 414898
rect 30300 414836 30306 414838
rect 38878 414292 38884 414356
rect 38948 414354 38954 414356
rect 38948 414294 60076 414354
rect 38948 414292 38954 414294
rect 44398 413748 44404 413812
rect 44468 413810 44474 413812
rect 44468 413750 60076 413810
rect 44468 413748 44474 413750
rect 36537 413266 36603 413269
rect 36537 413264 60076 413266
rect 36537 413208 36542 413264
rect 36598 413208 60076 413264
rect 36537 413206 60076 413208
rect 36537 413203 36603 413206
rect 54385 412722 54451 412725
rect 54385 412720 60076 412722
rect 54385 412664 54390 412720
rect 54446 412664 60076 412720
rect 54385 412662 60076 412664
rect 54385 412659 54451 412662
rect 35341 412178 35407 412181
rect 35341 412176 60076 412178
rect 35341 412120 35346 412176
rect 35402 412120 60076 412176
rect 35341 412118 60076 412120
rect 35341 412115 35407 412118
rect 54661 411634 54727 411637
rect 54661 411632 60076 411634
rect 54661 411576 54666 411632
rect 54722 411576 60076 411632
rect 54661 411574 60076 411576
rect 54661 411571 54727 411574
rect 55765 411090 55831 411093
rect 55765 411088 60076 411090
rect 55765 411032 55770 411088
rect 55826 411032 60076 411088
rect 55765 411030 60076 411032
rect 55765 411027 55831 411030
rect -960 410546 480 410636
rect 3918 410546 3924 410548
rect -960 410486 3924 410546
rect -960 410396 480 410486
rect 3918 410484 3924 410486
rect 3988 410484 3994 410548
rect 27245 410546 27311 410549
rect 27245 410544 60076 410546
rect 27245 410488 27250 410544
rect 27306 410488 60076 410544
rect 27245 410486 60076 410488
rect 27245 410483 27311 410486
rect 28441 410002 28507 410005
rect 28441 410000 60076 410002
rect 28441 409944 28446 410000
rect 28502 409944 60076 410000
rect 28441 409942 60076 409944
rect 28441 409939 28507 409942
rect 55949 409458 56015 409461
rect 55949 409456 60076 409458
rect 55949 409400 55954 409456
rect 56010 409400 60076 409456
rect 55949 409398 60076 409400
rect 55949 409395 56015 409398
rect 28349 408914 28415 408917
rect 28349 408912 60076 408914
rect 28349 408856 28354 408912
rect 28410 408856 60076 408912
rect 28349 408854 60076 408856
rect 28349 408851 28415 408854
rect 34237 408370 34303 408373
rect 34237 408368 60076 408370
rect 34237 408312 34242 408368
rect 34298 408312 60076 408368
rect 34237 408310 60076 408312
rect 34237 408307 34303 408310
rect 52177 407826 52243 407829
rect 508497 407826 508563 407829
rect 533337 407826 533403 407829
rect 52177 407824 60076 407826
rect 52177 407768 52182 407824
rect 52238 407768 60076 407824
rect 52177 407766 60076 407768
rect 508497 407824 533403 407826
rect 508497 407768 508502 407824
rect 508558 407768 533342 407824
rect 533398 407768 533403 407824
rect 508497 407766 533403 407768
rect 52177 407763 52243 407766
rect 508497 407763 508563 407766
rect 533337 407763 533403 407766
rect 51901 407282 51967 407285
rect 51901 407280 60076 407282
rect 51901 407224 51906 407280
rect 51962 407224 60076 407280
rect 51901 407222 60076 407224
rect 51901 407219 51967 407222
rect 56041 406738 56107 406741
rect 56041 406736 60076 406738
rect 56041 406680 56046 406736
rect 56102 406680 60076 406736
rect 56041 406678 60076 406680
rect 56041 406675 56107 406678
rect 38377 406194 38443 406197
rect 38377 406192 60076 406194
rect 38377 406136 38382 406192
rect 38438 406136 60076 406192
rect 38377 406134 60076 406136
rect 38377 406131 38443 406134
rect 40585 405650 40651 405653
rect 40585 405648 60076 405650
rect 40585 405592 40590 405648
rect 40646 405592 60076 405648
rect 40585 405590 60076 405592
rect 40585 405587 40651 405590
rect 36997 405106 37063 405109
rect 36997 405104 60076 405106
rect 36997 405048 37002 405104
rect 37058 405048 60076 405104
rect 36997 405046 60076 405048
rect 36997 405043 37063 405046
rect 500677 404970 500743 404973
rect 532877 404970 532943 404973
rect 583520 404970 584960 405060
rect 500677 404968 584960 404970
rect 500677 404912 500682 404968
rect 500738 404912 532882 404968
rect 532938 404912 584960 404968
rect 500677 404910 584960 404912
rect 500677 404907 500743 404910
rect 532877 404907 532943 404910
rect 583520 404820 584960 404910
rect 38193 404562 38259 404565
rect 38193 404560 60076 404562
rect 38193 404504 38198 404560
rect 38254 404504 60076 404560
rect 38193 404502 60076 404504
rect 38193 404499 38259 404502
rect 36721 404018 36787 404021
rect 36721 404016 60076 404018
rect 36721 403960 36726 404016
rect 36782 403960 60076 404016
rect 36721 403958 60076 403960
rect 36721 403955 36787 403958
rect 36813 403474 36879 403477
rect 36813 403472 60076 403474
rect 36813 403416 36818 403472
rect 36874 403416 60076 403472
rect 36813 403414 60076 403416
rect 36813 403411 36879 403414
rect 36905 402930 36971 402933
rect 36905 402928 60076 402930
rect 36905 402872 36910 402928
rect 36966 402872 60076 402928
rect 36905 402870 60076 402872
rect 36905 402867 36971 402870
rect 39389 402386 39455 402389
rect 39389 402384 60076 402386
rect 39389 402328 39394 402384
rect 39450 402328 60076 402384
rect 39389 402326 60076 402328
rect 39389 402323 39455 402326
rect 40677 401842 40743 401845
rect 40677 401840 60076 401842
rect 40677 401784 40682 401840
rect 40738 401784 60076 401840
rect 40677 401782 60076 401784
rect 40677 401779 40743 401782
rect 33961 401298 34027 401301
rect 33961 401296 60076 401298
rect 33961 401240 33966 401296
rect 34022 401240 60076 401296
rect 33961 401238 60076 401240
rect 33961 401235 34027 401238
rect 27061 400754 27127 400757
rect 27061 400752 60076 400754
rect 27061 400696 27066 400752
rect 27122 400696 60076 400752
rect 27061 400694 60076 400696
rect 27061 400691 27127 400694
rect 35433 400210 35499 400213
rect 35433 400208 60076 400210
rect 35433 400152 35438 400208
rect 35494 400152 60076 400208
rect 35433 400150 60076 400152
rect 35433 400147 35499 400150
rect 35525 399666 35591 399669
rect 35525 399664 60076 399666
rect 35525 399608 35530 399664
rect 35586 399608 60076 399664
rect 35525 399606 60076 399608
rect 35525 399603 35591 399606
rect 34145 399122 34211 399125
rect 34145 399120 60076 399122
rect 34145 399064 34150 399120
rect 34206 399064 60076 399120
rect 34145 399062 60076 399064
rect 34145 399059 34211 399062
rect 34053 398578 34119 398581
rect 34053 398576 60076 398578
rect 34053 398520 34058 398576
rect 34114 398520 60076 398576
rect 34053 398518 60076 398520
rect 34053 398515 34119 398518
rect 2814 398108 2820 398172
rect 2884 398170 2890 398172
rect 4061 398170 4127 398173
rect 2884 398168 4127 398170
rect 2884 398112 4066 398168
rect 4122 398112 4127 398168
rect 2884 398110 4127 398112
rect 2884 398108 2890 398110
rect 4061 398107 4127 398110
rect 35617 398034 35683 398037
rect 35617 398032 60076 398034
rect 35617 397976 35622 398032
rect 35678 397976 60076 398032
rect 35617 397974 60076 397976
rect 35617 397971 35683 397974
rect -960 397490 480 397580
rect 3550 397490 3556 397492
rect -960 397430 3556 397490
rect -960 397340 480 397430
rect 3550 397428 3556 397430
rect 3620 397428 3626 397492
rect 39297 397490 39363 397493
rect 39297 397488 60076 397490
rect 39297 397432 39302 397488
rect 39358 397432 60076 397488
rect 39297 397430 60076 397432
rect 39297 397427 39363 397430
rect 38285 396946 38351 396949
rect 38285 396944 60076 396946
rect 38285 396888 38290 396944
rect 38346 396888 60076 396944
rect 38285 396886 60076 396888
rect 38285 396883 38351 396886
rect 39573 396402 39639 396405
rect 39573 396400 60076 396402
rect 39573 396344 39578 396400
rect 39634 396344 60076 396400
rect 39573 396342 60076 396344
rect 39573 396339 39639 396342
rect 27429 395858 27495 395861
rect 27429 395856 60076 395858
rect 27429 395800 27434 395856
rect 27490 395800 60076 395856
rect 27429 395798 60076 395800
rect 27429 395795 27495 395798
rect 35801 395314 35867 395317
rect 35801 395312 60076 395314
rect 35801 395256 35806 395312
rect 35862 395256 60076 395312
rect 35801 395254 60076 395256
rect 35801 395251 35867 395254
rect 46841 394770 46907 394773
rect 46841 394768 60076 394770
rect 46841 394712 46846 394768
rect 46902 394712 60076 394768
rect 46841 394710 60076 394712
rect 46841 394707 46907 394710
rect 505369 394634 505435 394637
rect 508497 394634 508563 394637
rect 505369 394632 508563 394634
rect 505369 394576 505374 394632
rect 505430 394576 508502 394632
rect 508558 394576 508563 394632
rect 505369 394574 508563 394576
rect 505369 394571 505435 394574
rect 508497 394571 508563 394574
rect 28257 394226 28323 394229
rect 28257 394224 60076 394226
rect 28257 394168 28262 394224
rect 28318 394168 60076 394224
rect 28257 394166 60076 394168
rect 28257 394163 28323 394166
rect 26785 393682 26851 393685
rect 26785 393680 60076 393682
rect 26785 393624 26790 393680
rect 26846 393624 60076 393680
rect 26785 393622 60076 393624
rect 26785 393619 26851 393622
rect 31661 393138 31727 393141
rect 31661 393136 60076 393138
rect 31661 393080 31666 393136
rect 31722 393080 60076 393136
rect 31661 393078 60076 393080
rect 31661 393075 31727 393078
rect 33777 392594 33843 392597
rect 33777 392592 60076 392594
rect 33777 392536 33782 392592
rect 33838 392536 60076 392592
rect 33777 392534 60076 392536
rect 33777 392531 33843 392534
rect 33041 392050 33107 392053
rect 33041 392048 60076 392050
rect 33041 391992 33046 392048
rect 33102 391992 60076 392048
rect 33041 391990 60076 391992
rect 33041 391987 33107 391990
rect 499573 391914 499639 391917
rect 500585 391914 500651 391917
rect 499573 391912 500651 391914
rect 499573 391856 499578 391912
rect 499634 391856 500590 391912
rect 500646 391856 500651 391912
rect 499573 391854 500651 391856
rect 499573 391851 499639 391854
rect 500585 391851 500651 391854
rect 583520 391628 584960 391868
rect 30281 391506 30347 391509
rect 30281 391504 60076 391506
rect 30281 391448 30286 391504
rect 30342 391448 60076 391504
rect 30281 391446 60076 391448
rect 30281 391443 30347 391446
rect 30189 390962 30255 390965
rect 30189 390960 60076 390962
rect 30189 390904 30194 390960
rect 30250 390904 60076 390960
rect 30189 390902 60076 390904
rect 30189 390899 30255 390902
rect 59905 390690 59971 390693
rect 60917 390690 60983 390693
rect 59905 390688 60983 390690
rect 59905 390632 59910 390688
rect 59966 390632 60922 390688
rect 60978 390632 60983 390688
rect 59905 390630 60983 390632
rect 59905 390627 59971 390630
rect 60917 390627 60983 390630
rect 498285 390690 498351 390693
rect 501965 390690 502031 390693
rect 498285 390688 502031 390690
rect 498285 390632 498290 390688
rect 498346 390632 501970 390688
rect 502026 390632 502031 390688
rect 498285 390630 502031 390632
rect 498285 390627 498351 390630
rect 501965 390627 502031 390630
rect 323577 390418 323643 390421
rect 505369 390418 505435 390421
rect 323577 390416 505435 390418
rect 323577 390360 323582 390416
rect 323638 390360 505374 390416
rect 505430 390360 505435 390416
rect 323577 390358 505435 390360
rect 323577 390355 323643 390358
rect 505369 390355 505435 390358
rect 316585 390282 316651 390285
rect 316585 390280 325710 390282
rect 316585 390224 316590 390280
rect 316646 390224 325710 390280
rect 316585 390222 325710 390224
rect 316585 390219 316651 390222
rect 321829 390146 321895 390149
rect 325650 390146 325710 390222
rect 357934 390220 357940 390284
rect 358004 390282 358010 390284
rect 543222 390282 543228 390284
rect 358004 390222 543228 390282
rect 358004 390220 358010 390222
rect 543222 390220 543228 390222
rect 543292 390220 543298 390284
rect 528737 390146 528803 390149
rect 321829 390144 323226 390146
rect 321829 390088 321834 390144
rect 321890 390088 323226 390144
rect 321829 390086 323226 390088
rect 325650 390144 528803 390146
rect 325650 390088 528742 390144
rect 528798 390088 528803 390144
rect 325650 390086 528803 390088
rect 321829 390083 321895 390086
rect 323166 390010 323226 390086
rect 528737 390083 528803 390086
rect 501086 390010 501092 390012
rect 323166 389950 501092 390010
rect 501086 389948 501092 389950
rect 501156 389948 501162 390012
rect 224769 389874 224835 389877
rect 510705 389874 510771 389877
rect 224769 389872 510771 389874
rect 224769 389816 224774 389872
rect 224830 389816 510710 389872
rect 510766 389816 510771 389872
rect 224769 389814 510771 389816
rect 224769 389811 224835 389814
rect 510705 389811 510771 389814
rect 542905 389194 542971 389197
rect 543222 389194 543228 389196
rect 542905 389192 543228 389194
rect 542905 389136 542910 389192
rect 542966 389136 543228 389192
rect 542905 389134 543228 389136
rect 542905 389131 542971 389134
rect 543222 389132 543228 389134
rect 543292 389132 543298 389196
rect 60917 389058 60983 389061
rect 66897 389058 66963 389061
rect 60917 389056 66963 389058
rect 60917 389000 60922 389056
rect 60978 389000 66902 389056
rect 66958 389000 66963 389056
rect 60917 388998 66963 389000
rect 60917 388995 60983 388998
rect 66897 388995 66963 388998
rect 304349 389058 304415 389061
rect 500677 389058 500743 389061
rect 304349 389056 500743 389058
rect 304349 389000 304354 389056
rect 304410 389000 500682 389056
rect 500738 389000 500743 389056
rect 304349 388998 500743 389000
rect 304349 388995 304415 388998
rect 500677 388995 500743 388998
rect 318057 388922 318123 388925
rect 500493 388922 500559 388925
rect 318057 388920 500559 388922
rect 318057 388864 318062 388920
rect 318118 388864 500498 388920
rect 500554 388864 500559 388920
rect 318057 388862 500559 388864
rect 318057 388859 318123 388862
rect 500493 388859 500559 388862
rect 398925 388786 398991 388789
rect 546677 388786 546743 388789
rect 398925 388784 546743 388786
rect 398925 388728 398930 388784
rect 398986 388728 546682 388784
rect 546738 388728 546743 388784
rect 398925 388726 546743 388728
rect 398925 388723 398991 388726
rect 546677 388723 546743 388726
rect 345606 388588 345612 388652
rect 345676 388650 345682 388652
rect 538806 388650 538812 388652
rect 345676 388590 538812 388650
rect 345676 388588 345682 388590
rect 538806 388588 538812 388590
rect 538876 388588 538882 388652
rect 238661 388514 238727 388517
rect 538305 388514 538371 388517
rect 238661 388512 538371 388514
rect 238661 388456 238666 388512
rect 238722 388456 538310 388512
rect 538366 388456 538371 388512
rect 238661 388454 538371 388456
rect 238661 388451 238727 388454
rect 538305 388451 538371 388454
rect 238477 388378 238543 388381
rect 544285 388378 544351 388381
rect 238477 388376 544351 388378
rect 238477 388320 238482 388376
rect 238538 388320 544290 388376
rect 544346 388320 544351 388376
rect 238477 388318 544351 388320
rect 238477 388315 238543 388318
rect 544285 388315 544351 388318
rect 400213 388242 400279 388245
rect 548057 388242 548123 388245
rect 400213 388240 548123 388242
rect 400213 388184 400218 388240
rect 400274 388184 548062 388240
rect 548118 388184 548123 388240
rect 400213 388182 548123 388184
rect 400213 388179 400279 388182
rect 548057 388179 548123 388182
rect 233141 388106 233207 388109
rect 349797 388106 349863 388109
rect 233141 388104 349863 388106
rect 233141 388048 233146 388104
rect 233202 388048 349802 388104
rect 349858 388048 349863 388104
rect 233141 388046 349863 388048
rect 233141 388043 233207 388046
rect 349797 388043 349863 388046
rect 499941 388106 500007 388109
rect 500350 388106 500356 388108
rect 499941 388104 500356 388106
rect 499941 388048 499946 388104
rect 500002 388048 500356 388104
rect 499941 388046 500356 388048
rect 499941 388043 500007 388046
rect 500350 388044 500356 388046
rect 500420 388044 500426 388108
rect 227621 387970 227687 387973
rect 346301 387970 346367 387973
rect 227621 387968 346367 387970
rect 227621 387912 227626 387968
rect 227682 387912 346306 387968
rect 346362 387912 346367 387968
rect 227621 387910 346367 387912
rect 227621 387907 227687 387910
rect 346301 387907 346367 387910
rect 349654 387908 349660 387972
rect 349724 387970 349730 387972
rect 400305 387970 400371 387973
rect 349724 387968 400371 387970
rect 349724 387912 400310 387968
rect 400366 387912 400371 387968
rect 349724 387910 400371 387912
rect 349724 387908 349730 387910
rect 400305 387907 400371 387910
rect 231761 387834 231827 387837
rect 398833 387834 398899 387837
rect 231761 387832 398899 387834
rect 231761 387776 231766 387832
rect 231822 387776 398838 387832
rect 398894 387776 398899 387832
rect 231761 387774 398899 387776
rect 231761 387771 231827 387774
rect 398833 387771 398899 387774
rect 272885 387698 272951 387701
rect 279601 387698 279667 387701
rect 272885 387696 279667 387698
rect 272885 387640 272890 387696
rect 272946 387640 279606 387696
rect 279662 387640 279667 387696
rect 272885 387638 279667 387640
rect 272885 387635 272951 387638
rect 279601 387635 279667 387638
rect 480897 387698 480963 387701
rect 505093 387698 505159 387701
rect 480897 387696 505159 387698
rect 480897 387640 480902 387696
rect 480958 387640 505098 387696
rect 505154 387640 505159 387696
rect 480897 387638 505159 387640
rect 480897 387635 480963 387638
rect 505093 387635 505159 387638
rect 353293 387426 353359 387429
rect 360009 387426 360075 387429
rect 353293 387424 360075 387426
rect 353293 387368 353298 387424
rect 353354 387368 360014 387424
rect 360070 387368 360075 387424
rect 353293 387366 360075 387368
rect 353293 387363 353359 387366
rect 360009 387363 360075 387366
rect 491937 387426 492003 387429
rect 499481 387426 499547 387429
rect 491937 387424 499547 387426
rect 491937 387368 491942 387424
rect 491998 387368 499486 387424
rect 499542 387368 499547 387424
rect 491937 387366 499547 387368
rect 491937 387363 492003 387366
rect 499481 387363 499547 387366
rect 351545 387290 351611 387293
rect 357341 387290 357407 387293
rect 400213 387290 400279 387293
rect 351545 387288 400279 387290
rect 351545 387232 351550 387288
rect 351606 387232 357346 387288
rect 357402 387232 400218 387288
rect 400274 387232 400279 387288
rect 351545 387230 400279 387232
rect 351545 387227 351611 387230
rect 357341 387227 357407 387230
rect 400213 387227 400279 387230
rect 486141 387290 486207 387293
rect 500953 387290 501019 387293
rect 486141 387288 501019 387290
rect 486141 387232 486146 387288
rect 486202 387232 500958 387288
rect 501014 387232 501019 387288
rect 486141 387230 501019 387232
rect 486141 387227 486207 387230
rect 500953 387227 501019 387230
rect 262397 387154 262463 387157
rect 280061 387154 280127 387157
rect 262397 387152 280127 387154
rect 262397 387096 262402 387152
rect 262458 387096 280066 387152
rect 280122 387096 280127 387152
rect 262397 387094 280127 387096
rect 262397 387091 262463 387094
rect 280061 387091 280127 387094
rect 359825 387154 359891 387157
rect 417969 387154 418035 387157
rect 359825 387152 418035 387154
rect 359825 387096 359830 387152
rect 359886 387096 417974 387152
rect 418030 387096 418035 387152
rect 359825 387094 418035 387096
rect 359825 387091 359891 387094
rect 417969 387091 418035 387094
rect 484393 387154 484459 387157
rect 499757 387154 499823 387157
rect 484393 387152 499823 387154
rect 484393 387096 484398 387152
rect 484454 387096 499762 387152
rect 499818 387096 499823 387152
rect 484393 387094 499823 387096
rect 484393 387091 484459 387094
rect 499757 387091 499823 387094
rect 225689 387018 225755 387021
rect 279417 387018 279483 387021
rect 225689 387016 279483 387018
rect 225689 386960 225694 387016
rect 225750 386960 279422 387016
rect 279478 386960 279483 387016
rect 225689 386958 279483 386960
rect 225689 386955 225755 386958
rect 279417 386955 279483 386958
rect 350073 387018 350139 387021
rect 353937 387018 354003 387021
rect 398925 387018 398991 387021
rect 350073 387016 398991 387018
rect 350073 386960 350078 387016
rect 350134 386960 353942 387016
rect 353998 386960 398930 387016
rect 398986 386960 398991 387016
rect 350073 386958 398991 386960
rect 350073 386955 350139 386958
rect 353937 386955 354003 386958
rect 398925 386955 398991 386958
rect 403617 387018 403683 387021
rect 465165 387018 465231 387021
rect 403617 387016 465231 387018
rect 403617 386960 403622 387016
rect 403678 386960 465170 387016
rect 465226 386960 465231 387016
rect 403617 386958 465231 386960
rect 403617 386955 403683 386958
rect 465165 386955 465231 386958
rect 485865 387018 485931 387021
rect 502609 387018 502675 387021
rect 485865 387016 502675 387018
rect 485865 386960 485870 387016
rect 485926 386960 502614 387016
rect 502670 386960 502675 387016
rect 485865 386958 502675 386960
rect 485865 386955 485931 386958
rect 502609 386955 502675 386958
rect 283373 386882 283439 386885
rect 286685 386882 286751 386885
rect 283373 386880 286751 386882
rect 283373 386824 283378 386880
rect 283434 386824 286690 386880
rect 286746 386824 286751 386880
rect 283373 386822 286751 386824
rect 283373 386819 283439 386822
rect 286685 386819 286751 386822
rect 361614 386820 361620 386884
rect 361684 386882 361690 386884
rect 362033 386882 362099 386885
rect 361684 386880 362099 386882
rect 361684 386824 362038 386880
rect 362094 386824 362099 386880
rect 361684 386822 362099 386824
rect 361684 386820 361690 386822
rect 362033 386819 362099 386822
rect 362902 386820 362908 386884
rect 362972 386882 362978 386884
rect 363781 386882 363847 386885
rect 362972 386880 363847 386882
rect 362972 386824 363786 386880
rect 363842 386824 363847 386880
rect 362972 386822 363847 386824
rect 362972 386820 362978 386822
rect 363781 386819 363847 386822
rect 359641 386746 359707 386749
rect 360142 386746 360148 386748
rect 359641 386744 360148 386746
rect 359641 386688 359646 386744
rect 359702 386688 360148 386744
rect 359641 386686 360148 386688
rect 359641 386683 359707 386686
rect 360142 386684 360148 386686
rect 360212 386684 360218 386748
rect 360009 386610 360075 386613
rect 404261 386610 404327 386613
rect 360009 386608 404327 386610
rect 360009 386552 360014 386608
rect 360070 386552 404266 386608
rect 404322 386552 404327 386608
rect 360009 386550 404327 386552
rect 360009 386547 360075 386550
rect 404261 386547 404327 386550
rect 360193 386474 360259 386477
rect 360326 386474 360332 386476
rect 360193 386472 360332 386474
rect 360193 386416 360198 386472
rect 360254 386416 360332 386472
rect 360193 386414 360332 386416
rect 360193 386411 360259 386414
rect 360326 386412 360332 386414
rect 360396 386412 360402 386476
rect 265893 386338 265959 386341
rect 288157 386338 288223 386341
rect 265893 386336 288223 386338
rect 265893 386280 265898 386336
rect 265954 386280 288162 386336
rect 288218 386280 288223 386336
rect 265893 386278 288223 386280
rect 265893 386275 265959 386278
rect 288157 386275 288223 386278
rect 312537 386338 312603 386341
rect 537477 386338 537543 386341
rect 312537 386336 537543 386338
rect 312537 386280 312542 386336
rect 312598 386280 537482 386336
rect 537538 386280 537543 386336
rect 312537 386278 537543 386280
rect 312537 386275 312603 386278
rect 537477 386275 537543 386278
rect 216949 386202 217015 386205
rect 322381 386202 322447 386205
rect 216949 386200 322447 386202
rect 216949 386144 216954 386200
rect 217010 386144 322386 386200
rect 322442 386144 322447 386200
rect 216949 386142 322447 386144
rect 216949 386139 217015 386142
rect 322381 386139 322447 386142
rect 404261 386202 404327 386205
rect 546493 386202 546559 386205
rect 404261 386200 546559 386202
rect 404261 386144 404266 386200
rect 404322 386144 546498 386200
rect 546554 386144 546559 386200
rect 404261 386142 546559 386144
rect 404261 386139 404327 386142
rect 546493 386139 546559 386142
rect 134793 386066 134859 386069
rect 307017 386066 307083 386069
rect 134793 386064 307083 386066
rect 134793 386008 134798 386064
rect 134854 386008 307022 386064
rect 307078 386008 307083 386064
rect 134793 386006 307083 386008
rect 134793 386003 134859 386006
rect 307017 386003 307083 386006
rect 431217 386066 431283 386069
rect 502517 386066 502583 386069
rect 431217 386064 502583 386066
rect 431217 386008 431222 386064
rect 431278 386008 502522 386064
rect 502578 386008 502583 386064
rect 431217 386006 502583 386008
rect 431217 386003 431283 386006
rect 502517 386003 502583 386006
rect 265065 385930 265131 385933
rect 458173 385930 458239 385933
rect 265065 385928 458239 385930
rect 265065 385872 265070 385928
rect 265126 385872 458178 385928
rect 458234 385872 458239 385928
rect 265065 385870 458239 385872
rect 265065 385867 265131 385870
rect 458173 385867 458239 385870
rect 491293 385930 491359 385933
rect 498101 385930 498167 385933
rect 491293 385928 498167 385930
rect 491293 385872 491298 385928
rect 491354 385872 498106 385928
rect 498162 385872 498167 385928
rect 491293 385870 498167 385872
rect 491293 385867 491359 385870
rect 498101 385867 498167 385870
rect 96337 385794 96403 385797
rect 300117 385794 300183 385797
rect 96337 385792 300183 385794
rect 96337 385736 96342 385792
rect 96398 385736 300122 385792
rect 300178 385736 300183 385792
rect 96337 385734 300183 385736
rect 96337 385731 96403 385734
rect 300117 385731 300183 385734
rect 349838 385732 349844 385796
rect 349908 385794 349914 385796
rect 542629 385794 542695 385797
rect 349908 385792 542695 385794
rect 349908 385736 542634 385792
rect 542690 385736 542695 385792
rect 349908 385734 542695 385736
rect 349908 385732 349914 385734
rect 542629 385731 542695 385734
rect 282177 385658 282243 385661
rect 540237 385658 540303 385661
rect 282177 385656 540303 385658
rect 282177 385600 282182 385656
rect 282238 385600 540242 385656
rect 540298 385600 540303 385656
rect 282177 385598 540303 385600
rect 282177 385595 282243 385598
rect 540237 385595 540303 385598
rect 66897 384978 66963 384981
rect 68921 384978 68987 384981
rect 66897 384976 68987 384978
rect 66897 384920 66902 384976
rect 66958 384920 68926 384976
rect 68982 384920 68987 384976
rect 66897 384918 68987 384920
rect 66897 384915 66963 384918
rect 68921 384915 68987 384918
rect 80605 384978 80671 384981
rect 234613 384978 234679 384981
rect 379513 384978 379579 384981
rect 80605 384976 234679 384978
rect 80605 384920 80610 384976
rect 80666 384920 234618 384976
rect 234674 384920 234679 384976
rect 80605 384918 234679 384920
rect 80605 384915 80671 384918
rect 234613 384915 234679 384918
rect 238710 384976 379579 384978
rect 238710 384920 379518 384976
rect 379574 384920 379579 384976
rect 238710 384918 379579 384920
rect 235809 384842 235875 384845
rect 238710 384842 238770 384918
rect 379513 384915 379579 384918
rect 235809 384840 238770 384842
rect 235809 384784 235814 384840
rect 235870 384784 238770 384840
rect 235809 384782 238770 384784
rect 281625 384842 281691 384845
rect 292113 384842 292179 384845
rect 281625 384840 292179 384842
rect 281625 384784 281630 384840
rect 281686 384784 292118 384840
rect 292174 384784 292179 384840
rect 281625 384782 292179 384784
rect 235809 384779 235875 384782
rect 281625 384779 281691 384782
rect 292113 384779 292179 384782
rect 356646 384780 356652 384844
rect 356716 384842 356722 384844
rect 543774 384842 543780 384844
rect 356716 384782 543780 384842
rect 356716 384780 356722 384782
rect 543774 384780 543780 384782
rect 543844 384780 543850 384844
rect 152273 384706 152339 384709
rect 286501 384706 286567 384709
rect 152273 384704 286567 384706
rect 152273 384648 152278 384704
rect 152334 384648 286506 384704
rect 286562 384648 286567 384704
rect 152273 384646 286567 384648
rect 152273 384643 152339 384646
rect 286501 384643 286567 384646
rect 351126 384644 351132 384708
rect 351196 384706 351202 384708
rect 546534 384706 546540 384708
rect 351196 384646 546540 384706
rect 351196 384644 351202 384646
rect 546534 384644 546540 384646
rect 546604 384644 546610 384708
rect 143533 384570 143599 384573
rect 318149 384570 318215 384573
rect 143533 384568 318215 384570
rect -960 384284 480 384524
rect 143533 384512 143538 384568
rect 143594 384512 318154 384568
rect 318210 384512 318215 384568
rect 143533 384510 318215 384512
rect 143533 384507 143599 384510
rect 318149 384507 318215 384510
rect 346894 384508 346900 384572
rect 346964 384570 346970 384572
rect 550950 384570 550956 384572
rect 346964 384510 550956 384570
rect 346964 384508 346970 384510
rect 550950 384508 550956 384510
rect 551020 384508 551026 384572
rect 231669 384434 231735 384437
rect 487889 384434 487955 384437
rect 231669 384432 487955 384434
rect 231669 384376 231674 384432
rect 231730 384376 487894 384432
rect 487950 384376 487955 384432
rect 231669 384374 487955 384376
rect 231669 384371 231735 384374
rect 487889 384371 487955 384374
rect 231577 384298 231643 384301
rect 489637 384298 489703 384301
rect 231577 384296 489703 384298
rect 231577 384240 231582 384296
rect 231638 384240 489642 384296
rect 489698 384240 489703 384296
rect 231577 384238 489703 384240
rect 231577 384235 231643 384238
rect 489637 384235 489703 384238
rect 497457 384298 497523 384301
rect 502425 384298 502491 384301
rect 497457 384296 502491 384298
rect 497457 384240 497462 384296
rect 497518 384240 502430 384296
rect 502486 384240 502491 384296
rect 497457 384238 502491 384240
rect 497457 384235 497523 384238
rect 502425 384235 502491 384238
rect 233049 384162 233115 384165
rect 369025 384162 369091 384165
rect 233049 384160 369091 384162
rect 233049 384104 233054 384160
rect 233110 384104 369030 384160
rect 369086 384104 369091 384160
rect 233049 384102 369091 384104
rect 233049 384099 233115 384102
rect 369025 384099 369091 384102
rect 354622 383964 354628 384028
rect 354692 384026 354698 384028
rect 355961 384026 356027 384029
rect 354692 384024 356027 384026
rect 354692 383968 355966 384024
rect 356022 383968 356027 384024
rect 354692 383966 356027 383968
rect 354692 383964 354698 383966
rect 355961 383963 356027 383966
rect 353886 383828 353892 383892
rect 353956 383890 353962 383892
rect 357341 383890 357407 383893
rect 353956 383888 357407 383890
rect 353956 383832 357346 383888
rect 357402 383832 357407 383888
rect 353956 383830 357407 383832
rect 353956 383828 353962 383830
rect 357341 383827 357407 383830
rect 230381 383754 230447 383757
rect 282085 383754 282151 383757
rect 230381 383752 282151 383754
rect 230381 383696 230386 383752
rect 230442 383696 282090 383752
rect 282146 383696 282151 383752
rect 230381 383694 282151 383696
rect 230381 383691 230447 383694
rect 282085 383691 282151 383694
rect 183737 383346 183803 383349
rect 292021 383346 292087 383349
rect 183737 383344 292087 383346
rect 183737 383288 183742 383344
rect 183798 383288 292026 383344
rect 292082 383288 292087 383344
rect 183737 383286 292087 383288
rect 183737 383283 183803 383286
rect 292021 383283 292087 383286
rect 232773 383210 232839 383213
rect 416221 383210 416287 383213
rect 232773 383208 416287 383210
rect 232773 383152 232778 383208
rect 232834 383152 416226 383208
rect 416282 383152 416287 383208
rect 232773 383150 416287 383152
rect 232773 383147 232839 383150
rect 416221 383147 416287 383150
rect 471237 383210 471303 383213
rect 502701 383210 502767 383213
rect 471237 383208 502767 383210
rect 471237 383152 471242 383208
rect 471298 383152 502706 383208
rect 502762 383152 502767 383208
rect 471237 383150 502767 383152
rect 471237 383147 471303 383150
rect 502701 383147 502767 383150
rect 136541 383074 136607 383077
rect 294689 383074 294755 383077
rect 136541 383072 294755 383074
rect 136541 383016 136546 383072
rect 136602 383016 294694 383072
rect 294750 383016 294755 383072
rect 136541 383014 294755 383016
rect 136541 383011 136607 383014
rect 294689 383011 294755 383014
rect 358118 383012 358124 383076
rect 358188 383074 358194 383076
rect 542537 383074 542603 383077
rect 358188 383072 542603 383074
rect 358188 383016 542542 383072
rect 542598 383016 542603 383072
rect 358188 383014 542603 383016
rect 358188 383012 358194 383014
rect 542537 383011 542603 383014
rect 3734 382876 3740 382940
rect 3804 382938 3810 382940
rect 137134 382938 137140 382940
rect 3804 382878 137140 382938
rect 3804 382876 3810 382878
rect 137134 382876 137140 382878
rect 137204 382876 137210 382940
rect 229001 382938 229067 382941
rect 509417 382938 509483 382941
rect 229001 382936 509483 382938
rect 229001 382880 229006 382936
rect 229062 382880 509422 382936
rect 509478 382880 509483 382936
rect 229001 382878 509483 382880
rect 229001 382875 229067 382878
rect 509417 382875 509483 382878
rect 239673 382258 239739 382261
rect 321093 382258 321159 382261
rect 239673 382256 321159 382258
rect 239673 382200 239678 382256
rect 239734 382200 321098 382256
rect 321154 382200 321159 382256
rect 239673 382198 321159 382200
rect 239673 382195 239739 382198
rect 321093 382195 321159 382198
rect 356830 382196 356836 382260
rect 356900 382258 356906 382260
rect 542445 382258 542511 382261
rect 356900 382256 542511 382258
rect 356900 382200 542450 382256
rect 542506 382200 542511 382256
rect 356900 382198 542511 382200
rect 356900 382196 356906 382198
rect 542445 382195 542511 382198
rect 266905 382122 266971 382125
rect 461669 382122 461735 382125
rect 266905 382120 461735 382122
rect 266905 382064 266910 382120
rect 266966 382064 461674 382120
rect 461730 382064 461735 382120
rect 266905 382062 461735 382064
rect 266905 382059 266971 382062
rect 461669 382059 461735 382062
rect 69197 381986 69263 381989
rect 71773 381986 71839 381989
rect 69197 381984 71839 381986
rect 69197 381928 69202 381984
rect 69258 381928 71778 381984
rect 71834 381928 71839 381984
rect 69197 381926 71839 381928
rect 69197 381923 69263 381926
rect 71773 381923 71839 381926
rect 180241 381986 180307 381989
rect 296161 381986 296227 381989
rect 180241 381984 296227 381986
rect 180241 381928 180246 381984
rect 180302 381928 296166 381984
rect 296222 381928 296227 381984
rect 180241 381926 296227 381928
rect 180241 381923 180307 381926
rect 296161 381923 296227 381926
rect 355174 381924 355180 381988
rect 355244 381986 355250 381988
rect 550030 381986 550036 381988
rect 355244 381926 550036 381986
rect 355244 381924 355250 381926
rect 550030 381924 550036 381926
rect 550100 381924 550106 381988
rect 133045 381850 133111 381853
rect 289169 381850 289235 381853
rect 133045 381848 289235 381850
rect 133045 381792 133050 381848
rect 133106 381792 289174 381848
rect 289230 381792 289235 381848
rect 133045 381790 289235 381792
rect 133045 381787 133111 381790
rect 289169 381787 289235 381790
rect 338614 381788 338620 381852
rect 338684 381850 338690 381852
rect 550766 381850 550772 381852
rect 338684 381790 550772 381850
rect 338684 381788 338690 381790
rect 550766 381788 550772 381790
rect 550836 381788 550842 381852
rect 223481 381714 223547 381717
rect 507945 381714 508011 381717
rect 223481 381712 508011 381714
rect 223481 381656 223486 381712
rect 223542 381656 507950 381712
rect 508006 381656 508011 381712
rect 223481 381654 508011 381656
rect 223481 381651 223547 381654
rect 507945 381651 508011 381654
rect 231485 381578 231551 381581
rect 535637 381578 535703 381581
rect 231485 381576 535703 381578
rect 231485 381520 231490 381576
rect 231546 381520 535642 381576
rect 535698 381520 535703 381576
rect 231485 381518 535703 381520
rect 231485 381515 231551 381518
rect 535637 381515 535703 381518
rect 234337 381442 234403 381445
rect 398741 381442 398807 381445
rect 234337 381440 398807 381442
rect 234337 381384 234342 381440
rect 234398 381384 398746 381440
rect 398802 381384 398807 381440
rect 234337 381382 398807 381384
rect 234337 381379 234403 381382
rect 398741 381379 398807 381382
rect 230197 381170 230263 381173
rect 240041 381170 240107 381173
rect 230197 381168 240107 381170
rect 230197 381112 230202 381168
rect 230258 381112 240046 381168
rect 240102 381112 240107 381168
rect 230197 381110 240107 381112
rect 230197 381107 230263 381110
rect 240041 381107 240107 381110
rect 231393 381034 231459 381037
rect 266353 381034 266419 381037
rect 231393 381032 266419 381034
rect 231393 380976 231398 381032
rect 231454 380976 266358 381032
rect 266414 380976 266419 381032
rect 231393 380974 266419 380976
rect 231393 380971 231459 380974
rect 266353 380971 266419 380974
rect 490925 381034 490991 381037
rect 491937 381034 492003 381037
rect 490925 381032 492003 381034
rect 490925 380976 490930 381032
rect 490986 380976 491942 381032
rect 491998 380976 492003 381032
rect 490925 380974 492003 380976
rect 490925 380971 490991 380974
rect 491937 380971 492003 380974
rect 192477 380898 192543 380901
rect 320909 380898 320975 380901
rect 192477 380896 320975 380898
rect 192477 380840 192482 380896
rect 192538 380840 320914 380896
rect 320970 380840 320975 380896
rect 192477 380838 320975 380840
rect 192477 380835 192543 380838
rect 320909 380835 320975 380838
rect 237281 380762 237347 380765
rect 390001 380762 390067 380765
rect 237281 380760 390067 380762
rect 237281 380704 237286 380760
rect 237342 380704 390006 380760
rect 390062 380704 390067 380760
rect 237281 380702 390067 380704
rect 237281 380699 237347 380702
rect 390001 380699 390067 380702
rect 263225 380626 263291 380629
rect 454677 380626 454743 380629
rect 263225 380624 454743 380626
rect 263225 380568 263230 380624
rect 263286 380568 454682 380624
rect 454738 380568 454743 380624
rect 263225 380566 454743 380568
rect 263225 380563 263291 380566
rect 454677 380563 454743 380566
rect 70117 380490 70183 380493
rect 291837 380490 291903 380493
rect 70117 380488 291903 380490
rect 70117 380432 70122 380488
rect 70178 380432 291842 380488
rect 291898 380432 291903 380488
rect 70117 380430 291903 380432
rect 70117 380427 70183 380430
rect 291837 380427 291903 380430
rect 73613 380354 73679 380357
rect 304257 380354 304323 380357
rect 73613 380352 304323 380354
rect 73613 380296 73618 380352
rect 73674 380296 304262 380352
rect 304318 380296 304323 380352
rect 73613 380294 304323 380296
rect 73613 380291 73679 380294
rect 304257 380291 304323 380294
rect 71773 380218 71839 380221
rect 77569 380218 77635 380221
rect 71773 380216 77635 380218
rect 71773 380160 71778 380216
rect 71834 380160 77574 380216
rect 77630 380160 77635 380216
rect 71773 380158 77635 380160
rect 71773 380155 71839 380158
rect 77569 380155 77635 380158
rect 239806 380156 239812 380220
rect 239876 380218 239882 380220
rect 580206 380218 580212 380220
rect 239876 380158 580212 380218
rect 239876 380156 239882 380158
rect 580206 380156 580212 380158
rect 580276 380156 580282 380220
rect 169753 379402 169819 379405
rect 305729 379402 305795 379405
rect 169753 379400 305795 379402
rect 169753 379344 169758 379400
rect 169814 379344 305734 379400
rect 305790 379344 305795 379400
rect 169753 379342 305795 379344
rect 169753 379339 169819 379342
rect 305729 379339 305795 379342
rect 355542 379340 355548 379404
rect 355612 379402 355618 379404
rect 538622 379402 538628 379404
rect 355612 379342 538628 379402
rect 355612 379340 355618 379342
rect 538622 379340 538628 379342
rect 538692 379340 538698 379404
rect 547638 379340 547644 379404
rect 547708 379340 547714 379404
rect 122557 379266 122623 379269
rect 286317 379266 286383 379269
rect 122557 379264 286383 379266
rect 122557 379208 122562 379264
rect 122618 379208 286322 379264
rect 286378 379208 286383 379264
rect 122557 379206 286383 379208
rect 122557 379203 122623 379206
rect 286317 379203 286383 379206
rect 352966 379204 352972 379268
rect 353036 379266 353042 379268
rect 547646 379266 547706 379340
rect 353036 379206 547706 379266
rect 353036 379204 353042 379206
rect 238569 379130 238635 379133
rect 523861 379130 523927 379133
rect 238569 379128 523927 379130
rect 238569 379072 238574 379128
rect 238630 379072 523866 379128
rect 523922 379072 523927 379128
rect 238569 379070 523927 379072
rect 238569 379067 238635 379070
rect 523861 379067 523927 379070
rect 230105 378994 230171 378997
rect 518157 378994 518223 378997
rect 230105 378992 518223 378994
rect 230105 378936 230110 378992
rect 230166 378936 518162 378992
rect 518218 378936 518223 378992
rect 230105 378934 518223 378936
rect 230105 378931 230171 378934
rect 518157 378931 518223 378934
rect 228909 378858 228975 378861
rect 534165 378858 534231 378861
rect 228909 378856 534231 378858
rect 228909 378800 228914 378856
rect 228970 378800 534170 378856
rect 534226 378800 534231 378856
rect 228909 378798 534231 378800
rect 228909 378795 228975 378798
rect 534165 378795 534231 378798
rect 231301 378722 231367 378725
rect 536925 378722 536991 378725
rect 231301 378720 536991 378722
rect 231301 378664 231306 378720
rect 231362 378664 536930 378720
rect 536986 378664 536991 378720
rect 231301 378662 536991 378664
rect 231301 378659 231367 378662
rect 536925 378659 536991 378662
rect 233601 378586 233667 378589
rect 395245 378586 395311 378589
rect 233601 378584 395311 378586
rect 233601 378528 233606 378584
rect 233662 378528 395250 378584
rect 395306 378528 395311 378584
rect 233601 378526 395311 378528
rect 233601 378523 233667 378526
rect 395245 378523 395311 378526
rect 487337 378586 487403 378589
rect 491201 378586 491267 378589
rect 487337 378584 491267 378586
rect 487337 378528 487342 378584
rect 487398 378528 491206 378584
rect 491262 378528 491267 378584
rect 487337 378526 491267 378528
rect 487337 378523 487403 378526
rect 491201 378523 491267 378526
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 181989 378042 182055 378045
rect 294873 378042 294939 378045
rect 181989 378040 294939 378042
rect 181989 377984 181994 378040
rect 182050 377984 294878 378040
rect 294934 377984 294939 378040
rect 181989 377982 294939 377984
rect 181989 377979 182055 377982
rect 294873 377979 294939 377982
rect 487245 378042 487311 378045
rect 490925 378042 490991 378045
rect 487245 378040 490991 378042
rect 487245 377984 487250 378040
rect 487306 377984 490930 378040
rect 490986 377984 490991 378040
rect 487245 377982 490991 377984
rect 487245 377979 487311 377982
rect 490925 377979 490991 377982
rect 235809 377906 235875 377909
rect 376017 377906 376083 377909
rect 235809 377904 376083 377906
rect 235809 377848 235814 377904
rect 235870 377848 376022 377904
rect 376078 377848 376083 377904
rect 235809 377846 376083 377848
rect 235809 377843 235875 377846
rect 376017 377843 376083 377846
rect 235625 377770 235691 377773
rect 386505 377770 386571 377773
rect 235625 377768 386571 377770
rect 235625 377712 235630 377768
rect 235686 377712 386510 377768
rect 386566 377712 386571 377768
rect 235625 377710 386571 377712
rect 235625 377707 235691 377710
rect 386505 377707 386571 377710
rect 129549 377634 129615 377637
rect 293217 377634 293283 377637
rect 129549 377632 293283 377634
rect 129549 377576 129554 377632
rect 129610 377576 293222 377632
rect 293278 377576 293283 377632
rect 129549 377574 293283 377576
rect 129549 377571 129615 377574
rect 293217 377571 293283 377574
rect 234470 377436 234476 377500
rect 234540 377498 234546 377500
rect 414473 377498 414539 377501
rect 234540 377496 414539 377498
rect 234540 377440 414478 377496
rect 414534 377440 414539 377496
rect 234540 377438 414539 377440
rect 234540 377436 234546 377438
rect 414473 377435 414539 377438
rect 228817 377362 228883 377365
rect 531497 377362 531563 377365
rect 228817 377360 531563 377362
rect 228817 377304 228822 377360
rect 228878 377304 531502 377360
rect 531558 377304 531563 377360
rect 228817 377302 531563 377304
rect 228817 377299 228883 377302
rect 531497 377299 531563 377302
rect 77569 377090 77635 377093
rect 80697 377090 80763 377093
rect 77569 377088 80763 377090
rect 77569 377032 77574 377088
rect 77630 377032 80702 377088
rect 80758 377032 80763 377088
rect 77569 377030 80763 377032
rect 77569 377027 77635 377030
rect 80697 377027 80763 377030
rect 235717 376682 235783 376685
rect 383009 376682 383075 376685
rect 235717 376680 383075 376682
rect 235717 376624 235722 376680
rect 235778 376624 383014 376680
rect 383070 376624 383075 376680
rect 235717 376622 383075 376624
rect 235717 376619 235783 376622
rect 383009 376619 383075 376622
rect 485405 376682 485471 376685
rect 487337 376682 487403 376685
rect 485405 376680 487403 376682
rect 485405 376624 485410 376680
rect 485466 376624 487342 376680
rect 487398 376624 487403 376680
rect 485405 376622 487403 376624
rect 485405 376619 485471 376622
rect 487337 376619 487403 376622
rect 141785 376546 141851 376549
rect 295977 376546 296043 376549
rect 141785 376544 296043 376546
rect 141785 376488 141790 376544
rect 141846 376488 295982 376544
rect 296038 376488 296043 376544
rect 141785 376486 296043 376488
rect 141785 376483 141851 376486
rect 295977 376483 296043 376486
rect 354070 376484 354076 376548
rect 354140 376546 354146 376548
rect 550582 376546 550588 376548
rect 354140 376486 550588 376546
rect 354140 376484 354146 376486
rect 550582 376484 550588 376486
rect 550652 376484 550658 376548
rect 227529 376410 227595 376413
rect 528001 376410 528067 376413
rect 227529 376408 528067 376410
rect 227529 376352 227534 376408
rect 227590 376352 528006 376408
rect 528062 376352 528067 376408
rect 227529 376350 528067 376352
rect 227529 376347 227595 376350
rect 528001 376347 528067 376350
rect 223389 376274 223455 376277
rect 528645 376274 528711 376277
rect 223389 376272 528711 376274
rect 223389 376216 223394 376272
rect 223450 376216 528650 376272
rect 528706 376216 528711 376272
rect 223389 376214 528711 376216
rect 223389 376211 223455 376214
rect 528645 376211 528711 376214
rect 228725 376138 228791 376141
rect 534073 376138 534139 376141
rect 228725 376136 534139 376138
rect 228725 376080 228730 376136
rect 228786 376080 534078 376136
rect 534134 376080 534139 376136
rect 228725 376078 534139 376080
rect 228725 376075 228791 376078
rect 534073 376075 534139 376078
rect 226241 376002 226307 376005
rect 532693 376002 532759 376005
rect 226241 376000 532759 376002
rect 226241 375944 226246 376000
rect 226302 375944 532698 376000
rect 532754 375944 532759 376000
rect 226241 375942 532759 375944
rect 226241 375939 226307 375942
rect 532693 375939 532759 375942
rect 195973 375866 196039 375869
rect 309869 375866 309935 375869
rect 195973 375864 309935 375866
rect 195973 375808 195978 375864
rect 196034 375808 309874 375864
rect 309930 375808 309935 375864
rect 195973 375806 309935 375808
rect 195973 375803 196039 375806
rect 309869 375803 309935 375806
rect 485773 375866 485839 375869
rect 487245 375866 487311 375869
rect 485773 375864 487311 375866
rect 485773 375808 485778 375864
rect 485834 375808 487250 375864
rect 487306 375808 487311 375864
rect 485773 375806 487311 375808
rect 485773 375803 485839 375806
rect 487245 375803 487311 375806
rect 230013 375458 230079 375461
rect 234613 375458 234679 375461
rect 230013 375456 234679 375458
rect 230013 375400 230018 375456
rect 230074 375400 234618 375456
rect 234674 375400 234679 375456
rect 230013 375398 234679 375400
rect 230013 375395 230079 375398
rect 234613 375395 234679 375398
rect 357198 375396 357204 375460
rect 357268 375458 357274 375460
rect 485957 375458 486023 375461
rect 357268 375456 486023 375458
rect 357268 375400 485962 375456
rect 486018 375400 486023 375456
rect 357268 375398 486023 375400
rect 357268 375396 357274 375398
rect 485957 375395 486023 375398
rect 234429 375322 234495 375325
rect 290733 375322 290799 375325
rect 234429 375320 290799 375322
rect 234429 375264 234434 375320
rect 234490 375264 290738 375320
rect 290794 375264 290799 375320
rect 234429 375262 290799 375264
rect 234429 375259 234495 375262
rect 290733 375259 290799 375262
rect 171501 375186 171567 375189
rect 284886 375186 284892 375188
rect 171501 375184 284892 375186
rect 171501 375128 171506 375184
rect 171562 375128 284892 375184
rect 171501 375126 284892 375128
rect 171501 375123 171567 375126
rect 284886 375124 284892 375126
rect 284956 375124 284962 375188
rect 178493 375050 178559 375053
rect 307201 375050 307267 375053
rect 178493 375048 307267 375050
rect 178493 374992 178498 375048
rect 178554 374992 307206 375048
rect 307262 374992 307267 375048
rect 178493 374990 307267 374992
rect 178493 374987 178559 374990
rect 307201 374987 307267 374990
rect 234153 374914 234219 374917
rect 400489 374914 400555 374917
rect 234153 374912 400555 374914
rect 234153 374856 234158 374912
rect 234214 374856 400494 374912
rect 400550 374856 400555 374912
rect 234153 374854 400555 374856
rect 234153 374851 234219 374854
rect 400489 374851 400555 374854
rect 282126 374716 282132 374780
rect 282196 374778 282202 374780
rect 538254 374778 538260 374780
rect 282196 374718 538260 374778
rect 282196 374716 282202 374718
rect 538254 374716 538260 374718
rect 538324 374716 538330 374780
rect 236729 374642 236795 374645
rect 529381 374642 529447 374645
rect 236729 374640 529447 374642
rect 236729 374584 236734 374640
rect 236790 374584 529386 374640
rect 529442 374584 529447 374640
rect 236729 374582 529447 374584
rect 236729 374579 236795 374582
rect 529381 374579 529447 374582
rect 235533 373962 235599 373965
rect 381261 373962 381327 373965
rect 235533 373960 381327 373962
rect 235533 373904 235538 373960
rect 235594 373904 381266 373960
rect 381322 373904 381327 373960
rect 235533 373902 381327 373904
rect 235533 373899 235599 373902
rect 381261 373899 381327 373902
rect 140037 373826 140103 373829
rect 290457 373826 290523 373829
rect 140037 373824 290523 373826
rect 140037 373768 140042 373824
rect 140098 373768 290462 373824
rect 290518 373768 290523 373824
rect 140037 373766 290523 373768
rect 140037 373763 140103 373766
rect 290457 373763 290523 373766
rect 277025 373690 277091 373693
rect 504725 373690 504791 373693
rect 277025 373688 504791 373690
rect 277025 373632 277030 373688
rect 277086 373632 504730 373688
rect 504786 373632 504791 373688
rect 277025 373630 504791 373632
rect 277025 373627 277091 373630
rect 504725 373627 504791 373630
rect 78857 373554 78923 373557
rect 315389 373554 315455 373557
rect 78857 373552 315455 373554
rect 78857 373496 78862 373552
rect 78918 373496 315394 373552
rect 315450 373496 315455 373552
rect 78857 373494 315455 373496
rect 78857 373491 78923 373494
rect 315389 373491 315455 373494
rect 264145 373418 264211 373421
rect 280889 373418 280955 373421
rect 264145 373416 280955 373418
rect 264145 373360 264150 373416
rect 264206 373360 280894 373416
rect 280950 373360 280955 373416
rect 264145 373358 280955 373360
rect 264145 373355 264211 373358
rect 280889 373355 280955 373358
rect 282310 373356 282316 373420
rect 282380 373418 282386 373420
rect 541014 373418 541020 373420
rect 282380 373358 541020 373418
rect 282380 373356 282386 373358
rect 541014 373356 541020 373358
rect 541084 373356 541090 373420
rect 226149 373282 226215 373285
rect 535453 373282 535519 373285
rect 226149 373280 535519 373282
rect 226149 373224 226154 373280
rect 226210 373224 535458 373280
rect 535514 373224 535519 373280
rect 226149 373222 535519 373224
rect 226149 373219 226215 373222
rect 535453 373219 535519 373222
rect 232681 373146 232747 373149
rect 358261 373146 358327 373149
rect 232681 373144 358327 373146
rect 232681 373088 232686 373144
rect 232742 373088 358266 373144
rect 358322 373088 358327 373144
rect 232681 373086 358327 373088
rect 232681 373083 232747 373086
rect 358261 373083 358327 373086
rect 236821 372738 236887 372741
rect 276013 372738 276079 372741
rect 236821 372736 276079 372738
rect 236821 372680 236826 372736
rect 236882 372680 276018 372736
rect 276074 372680 276079 372736
rect 236821 372678 276079 372680
rect 236821 372675 236887 372678
rect 276013 372675 276079 372678
rect 482277 372738 482343 372741
rect 485773 372738 485839 372741
rect 482277 372736 485839 372738
rect 482277 372680 482282 372736
rect 482338 372680 485778 372736
rect 485834 372680 485839 372736
rect 482277 372678 485839 372680
rect 482277 372675 482343 372678
rect 485773 372675 485839 372678
rect 236177 372466 236243 372469
rect 294965 372466 295031 372469
rect 236177 372464 295031 372466
rect 236177 372408 236182 372464
rect 236238 372408 294970 372464
rect 295026 372408 295031 372464
rect 236177 372406 295031 372408
rect 236177 372403 236243 372406
rect 294965 372403 295031 372406
rect 211705 372330 211771 372333
rect 284937 372330 285003 372333
rect 211705 372328 285003 372330
rect 211705 372272 211710 372328
rect 211766 372272 284942 372328
rect 284998 372272 285003 372328
rect 211705 372270 285003 372272
rect 211705 372267 211771 372270
rect 284937 372267 285003 372270
rect 234245 372194 234311 372197
rect 391749 372194 391815 372197
rect 234245 372192 391815 372194
rect 234245 372136 234250 372192
rect 234306 372136 391754 372192
rect 391810 372136 391815 372192
rect 234245 372134 391815 372136
rect 234245 372131 234311 372134
rect 391749 372131 391815 372134
rect 185485 372058 185551 372061
rect 301589 372058 301655 372061
rect 185485 372056 301655 372058
rect 185485 372000 185490 372056
rect 185546 372000 301594 372056
rect 301650 372000 301655 372056
rect 185485 371998 301655 372000
rect 185485 371995 185551 371998
rect 301589 371995 301655 371998
rect 351310 371996 351316 372060
rect 351380 372058 351386 372060
rect 543222 372058 543228 372060
rect 351380 371998 543228 372058
rect 351380 371996 351386 371998
rect 543222 371996 543228 371998
rect 543292 371996 543298 372060
rect 282361 371922 282427 371925
rect 540145 371922 540211 371925
rect 282361 371920 540211 371922
rect 282361 371864 282366 371920
rect 282422 371864 540150 371920
rect 540206 371864 540211 371920
rect 282361 371862 540211 371864
rect 282361 371859 282427 371862
rect 540145 371859 540211 371862
rect 482829 371786 482895 371789
rect 485405 371786 485471 371789
rect 482829 371784 485471 371786
rect 482829 371728 482834 371784
rect 482890 371728 485410 371784
rect 485466 371728 485471 371784
rect 482829 371726 485471 371728
rect 482829 371723 482895 371726
rect 485405 371723 485471 371726
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 542353 371378 542419 371381
rect 542670 371378 542676 371380
rect 542353 371376 542676 371378
rect 542353 371320 542358 371376
rect 542414 371320 542676 371376
rect 542353 371318 542676 371320
rect 542353 371315 542419 371318
rect 542670 371316 542676 371318
rect 542740 371316 542746 371380
rect 276657 371242 276723 371245
rect 287830 371242 287836 371244
rect 276657 371240 287836 371242
rect 276657 371184 276662 371240
rect 276718 371184 287836 371240
rect 276657 371182 287836 371184
rect 276657 371179 276723 371182
rect 287830 371180 287836 371182
rect 287900 371180 287906 371244
rect 229185 371106 229251 371109
rect 305913 371106 305979 371109
rect 229185 371104 305979 371106
rect 229185 371048 229190 371104
rect 229246 371048 305918 371104
rect 305974 371048 305979 371104
rect 229185 371046 305979 371048
rect 229185 371043 229251 371046
rect 305913 371043 305979 371046
rect 176745 370970 176811 370973
rect 288065 370970 288131 370973
rect 176745 370968 288131 370970
rect 176745 370912 176750 370968
rect 176806 370912 288070 370968
rect 288126 370912 288131 370968
rect 176745 370910 288131 370912
rect 176745 370907 176811 370910
rect 288065 370907 288131 370910
rect 127801 370834 127867 370837
rect 291929 370834 291995 370837
rect 127801 370832 291995 370834
rect 127801 370776 127806 370832
rect 127862 370776 291934 370832
rect 291990 370776 291995 370832
rect 127801 370774 291995 370776
rect 127801 370771 127867 370774
rect 291929 370771 291995 370774
rect 233877 370698 233943 370701
rect 405733 370698 405799 370701
rect 233877 370696 405799 370698
rect 233877 370640 233882 370696
rect 233938 370640 405738 370696
rect 405794 370640 405799 370696
rect 233877 370638 405799 370640
rect 233877 370635 233943 370638
rect 405733 370635 405799 370638
rect 282678 370500 282684 370564
rect 282748 370562 282754 370564
rect 541198 370562 541204 370564
rect 282748 370502 541204 370562
rect 282748 370500 282754 370502
rect 541198 370500 541204 370502
rect 541268 370500 541274 370564
rect 478873 369882 478939 369885
rect 482829 369882 482895 369885
rect 478873 369880 482895 369882
rect 478873 369824 478878 369880
rect 478934 369824 482834 369880
rect 482890 369824 482895 369880
rect 478873 369822 482895 369824
rect 478873 369819 478939 369822
rect 482829 369819 482895 369822
rect 223941 369474 224007 369477
rect 303245 369474 303311 369477
rect 223941 369472 303311 369474
rect 223941 369416 223946 369472
rect 224002 369416 303250 369472
rect 303306 369416 303311 369472
rect 223941 369414 303311 369416
rect 223941 369411 224007 369414
rect 303245 369411 303311 369414
rect 194225 369338 194291 369341
rect 297449 369338 297515 369341
rect 194225 369336 297515 369338
rect 194225 369280 194230 369336
rect 194286 369280 297454 369336
rect 297510 369280 297515 369336
rect 194225 369278 297515 369280
rect 194225 369275 194291 369278
rect 297449 369275 297515 369278
rect 234061 369202 234127 369205
rect 393497 369202 393563 369205
rect 234061 369200 393563 369202
rect 234061 369144 234066 369200
rect 234122 369144 393502 369200
rect 393558 369144 393563 369200
rect 234061 369142 393563 369144
rect 234061 369139 234127 369142
rect 393497 369139 393563 369142
rect 237925 369066 237991 369069
rect 280797 369066 280863 369069
rect 237925 369064 280863 369066
rect 237925 369008 237930 369064
rect 237986 369008 280802 369064
rect 280858 369008 280863 369064
rect 237925 369006 280863 369008
rect 237925 369003 237991 369006
rect 280797 369003 280863 369006
rect 282494 369004 282500 369068
rect 282564 369066 282570 369068
rect 539358 369066 539364 369068
rect 282564 369006 539364 369066
rect 282564 369004 282570 369006
rect 539358 369004 539364 369006
rect 539428 369004 539434 369068
rect 204713 368250 204779 368253
rect 319621 368250 319687 368253
rect 204713 368248 319687 368250
rect 204713 368192 204718 368248
rect 204774 368192 319626 368248
rect 319682 368192 319687 368248
rect 204713 368190 319687 368192
rect 204713 368187 204779 368190
rect 319621 368187 319687 368190
rect 234521 368114 234587 368117
rect 370773 368114 370839 368117
rect 234521 368112 370839 368114
rect 234521 368056 234526 368112
rect 234582 368056 370778 368112
rect 370834 368056 370839 368112
rect 234521 368054 370839 368056
rect 234521 368051 234587 368054
rect 370773 368051 370839 368054
rect 166257 367978 166323 367981
rect 314193 367978 314259 367981
rect 166257 367976 314259 367978
rect 166257 367920 166262 367976
rect 166318 367920 314198 367976
rect 314254 367920 314259 367976
rect 166257 367918 314259 367920
rect 166257 367915 166323 367918
rect 314193 367915 314259 367918
rect 232589 367842 232655 367845
rect 412725 367842 412791 367845
rect 232589 367840 412791 367842
rect 232589 367784 232594 367840
rect 232650 367784 412730 367840
rect 412786 367784 412791 367840
rect 232589 367782 412791 367784
rect 232589 367779 232655 367782
rect 412725 367779 412791 367782
rect 81433 367706 81499 367709
rect 88149 367706 88215 367709
rect 81433 367704 88215 367706
rect 81433 367648 81438 367704
rect 81494 367648 88154 367704
rect 88210 367648 88215 367704
rect 81433 367646 88215 367648
rect 81433 367643 81499 367646
rect 88149 367643 88215 367646
rect 119061 367706 119127 367709
rect 298737 367706 298803 367709
rect 119061 367704 298803 367706
rect 119061 367648 119066 367704
rect 119122 367648 298742 367704
rect 298798 367648 298803 367704
rect 119061 367646 298803 367648
rect 119061 367643 119127 367646
rect 298737 367643 298803 367646
rect 352782 367644 352788 367708
rect 352852 367706 352858 367708
rect 542854 367706 542860 367708
rect 352852 367646 542860 367706
rect 352852 367644 352858 367646
rect 542854 367644 542860 367646
rect 542924 367644 542930 367708
rect 476389 367026 476455 367029
rect 478873 367026 478939 367029
rect 476389 367024 478939 367026
rect 476389 366968 476394 367024
rect 476450 366968 478878 367024
rect 478934 366968 478939 367024
rect 476389 366966 478939 366968
rect 476389 366963 476455 366966
rect 478873 366963 478939 366966
rect 213453 366754 213519 366757
rect 299013 366754 299079 366757
rect 213453 366752 299079 366754
rect 213453 366696 213458 366752
rect 213514 366696 299018 366752
rect 299074 366696 299079 366752
rect 213453 366694 299079 366696
rect 213453 366691 213519 366694
rect 299013 366691 299079 366694
rect 168005 366618 168071 366621
rect 323669 366618 323735 366621
rect 168005 366616 323735 366618
rect 168005 366560 168010 366616
rect 168066 366560 323674 366616
rect 323730 366560 323735 366616
rect 168005 366558 323735 366560
rect 168005 366555 168071 366558
rect 323669 366555 323735 366558
rect 234286 366420 234292 366484
rect 234356 366482 234362 366484
rect 410977 366482 411043 366485
rect 234356 366480 411043 366482
rect 234356 366424 410982 366480
rect 411038 366424 411043 366480
rect 234356 366422 411043 366424
rect 234356 366420 234362 366422
rect 410977 366419 411043 366422
rect 120809 366346 120875 366349
rect 302969 366346 303035 366349
rect 120809 366344 303035 366346
rect 120809 366288 120814 366344
rect 120870 366288 302974 366344
rect 303030 366288 303035 366344
rect 120809 366286 303035 366288
rect 120809 366283 120875 366286
rect 302969 366283 303035 366286
rect 88149 365802 88215 365805
rect 94497 365802 94563 365805
rect 88149 365800 94563 365802
rect 88149 365744 88154 365800
rect 88210 365744 94502 365800
rect 94558 365744 94563 365800
rect 88149 365742 94563 365744
rect 88149 365739 88215 365742
rect 94497 365739 94563 365742
rect 202965 365666 203031 365669
rect 311433 365666 311499 365669
rect 202965 365664 311499 365666
rect 202965 365608 202970 365664
rect 203026 365608 311438 365664
rect 311494 365608 311499 365664
rect 202965 365606 311499 365608
rect 202965 365603 203031 365606
rect 311433 365603 311499 365606
rect 237189 365530 237255 365533
rect 384757 365530 384823 365533
rect 237189 365528 384823 365530
rect 237189 365472 237194 365528
rect 237250 365472 384762 365528
rect 384818 365472 384823 365528
rect 237189 365470 384823 365472
rect 237189 365467 237255 365470
rect 384757 365467 384823 365470
rect 154021 365394 154087 365397
rect 298921 365394 298987 365397
rect 154021 365392 298987 365394
rect 154021 365336 154026 365392
rect 154082 365336 298926 365392
rect 298982 365336 298987 365392
rect 154021 365334 298987 365336
rect 154021 365331 154087 365334
rect 298921 365331 298987 365334
rect 357014 365332 357020 365396
rect 357084 365394 357090 365396
rect 543406 365394 543412 365396
rect 357084 365334 543412 365394
rect 357084 365332 357090 365334
rect 543406 365332 543412 365334
rect 543476 365332 543482 365396
rect 106825 365258 106891 365261
rect 286409 365258 286475 365261
rect 106825 365256 286475 365258
rect 106825 365200 106830 365256
rect 106886 365200 286414 365256
rect 286470 365200 286475 365256
rect 106825 365198 286475 365200
rect 106825 365195 106891 365198
rect 286409 365195 286475 365198
rect 354254 365196 354260 365260
rect 354324 365258 354330 365260
rect 542670 365258 542676 365260
rect 354324 365198 542676 365258
rect 354324 365196 354330 365198
rect 542670 365196 542676 365198
rect 542740 365196 542746 365260
rect 264145 365122 264211 365125
rect 456425 365122 456491 365125
rect 264145 365120 456491 365122
rect 264145 365064 264150 365120
rect 264206 365064 456430 365120
rect 456486 365064 456491 365120
rect 264145 365062 456491 365064
rect 264145 365059 264211 365062
rect 456425 365059 456491 365062
rect 580206 365060 580212 365124
rect 580276 365122 580282 365124
rect 583520 365122 584960 365212
rect 580276 365062 584960 365122
rect 580276 365060 580282 365062
rect 234102 364924 234108 364988
rect 234172 364986 234178 364988
rect 516961 364986 517027 364989
rect 234172 364984 517027 364986
rect 234172 364928 516966 364984
rect 517022 364928 517027 364984
rect 583520 364972 584960 365062
rect 234172 364926 517027 364928
rect 234172 364924 234178 364926
rect 516961 364923 517027 364926
rect 227437 364306 227503 364309
rect 300485 364306 300551 364309
rect 227437 364304 300551 364306
rect 227437 364248 227442 364304
rect 227498 364248 300490 364304
rect 300546 364248 300551 364304
rect 227437 364246 300551 364248
rect 227437 364243 227503 364246
rect 300485 364243 300551 364246
rect 159265 364170 159331 364173
rect 303153 364170 303219 364173
rect 159265 364168 303219 364170
rect 159265 364112 159270 364168
rect 159326 364112 303158 364168
rect 303214 364112 303219 364168
rect 159265 364110 303219 364112
rect 159265 364107 159331 364110
rect 303153 364107 303219 364110
rect 235073 364034 235139 364037
rect 396993 364034 397059 364037
rect 235073 364032 397059 364034
rect 235073 363976 235078 364032
rect 235134 363976 396998 364032
rect 397054 363976 397059 364032
rect 235073 363974 397059 363976
rect 235073 363971 235139 363974
rect 396993 363971 397059 363974
rect 265985 363898 266051 363901
rect 459921 363898 459987 363901
rect 265985 363896 459987 363898
rect 265985 363840 265990 363896
rect 266046 363840 459926 363896
rect 459982 363840 459987 363896
rect 265985 363838 459987 363840
rect 265985 363835 266051 363838
rect 459921 363835 459987 363838
rect 238293 363762 238359 363765
rect 522481 363762 522547 363765
rect 238293 363760 522547 363762
rect 238293 363704 238298 363760
rect 238354 363704 522486 363760
rect 522542 363704 522547 363760
rect 238293 363702 522547 363704
rect 238293 363699 238359 363702
rect 522481 363699 522547 363702
rect 46013 363626 46079 363629
rect 341609 363626 341675 363629
rect 46013 363624 341675 363626
rect 46013 363568 46018 363624
rect 46074 363568 341614 363624
rect 341670 363568 341675 363624
rect 46013 363566 341675 363568
rect 46013 363563 46079 363566
rect 341609 363563 341675 363566
rect 355358 363564 355364 363628
rect 355428 363626 355434 363628
rect 543038 363626 543044 363628
rect 355428 363566 543044 363626
rect 355428 363564 355434 363566
rect 543038 363564 543044 363566
rect 543108 363564 543114 363628
rect 482277 363218 482343 363221
rect 480210 363216 482343 363218
rect 480210 363160 482282 363216
rect 482338 363160 482343 363216
rect 480210 363158 482343 363160
rect 209957 362946 210023 362949
rect 293493 362946 293559 362949
rect 209957 362944 293559 362946
rect 209957 362888 209962 362944
rect 210018 362888 293498 362944
rect 293554 362888 293559 362944
rect 209957 362886 293559 362888
rect 209957 362883 210023 362886
rect 293493 362883 293559 362886
rect 479517 362946 479583 362949
rect 480210 362946 480270 363158
rect 482277 363155 482343 363158
rect 479517 362944 480270 362946
rect 479517 362888 479522 362944
rect 479578 362888 480270 362944
rect 479517 362886 480270 362888
rect 479517 362883 479583 362886
rect 232957 362810 233023 362813
rect 367277 362810 367343 362813
rect 232957 362808 367343 362810
rect 232957 362752 232962 362808
rect 233018 362752 367282 362808
rect 367338 362752 367343 362808
rect 232957 362750 367343 362752
rect 232957 362747 233023 362750
rect 367277 362747 367343 362750
rect 235441 362674 235507 362677
rect 377765 362674 377831 362677
rect 235441 362672 377831 362674
rect 235441 362616 235446 362672
rect 235502 362616 377770 362672
rect 377826 362616 377831 362672
rect 235441 362614 377831 362616
rect 235441 362611 235507 362614
rect 377765 362611 377831 362614
rect 161013 362538 161079 362541
rect 304441 362538 304507 362541
rect 161013 362536 304507 362538
rect 161013 362480 161018 362536
rect 161074 362480 304446 362536
rect 304502 362480 304507 362536
rect 161013 362478 304507 362480
rect 161013 362475 161079 362478
rect 304441 362475 304507 362478
rect 282637 362402 282703 362405
rect 540053 362402 540119 362405
rect 282637 362400 540119 362402
rect 282637 362344 282642 362400
rect 282698 362344 540058 362400
rect 540114 362344 540119 362400
rect 282637 362342 540119 362344
rect 282637 362339 282703 362342
rect 540053 362339 540119 362342
rect 239622 362204 239628 362268
rect 239692 362266 239698 362268
rect 580390 362266 580396 362268
rect 239692 362206 580396 362266
rect 239692 362204 239698 362206
rect 580390 362204 580396 362206
rect 580460 362204 580466 362268
rect 473261 362130 473327 362133
rect 476389 362130 476455 362133
rect 473261 362128 476455 362130
rect 473261 362072 473266 362128
rect 473322 362072 476394 362128
rect 476450 362072 476455 362128
rect 473261 362070 476455 362072
rect 473261 362067 473327 362070
rect 476389 362067 476455 362070
rect 208209 361586 208275 361589
rect 318241 361586 318307 361589
rect 208209 361584 318307 361586
rect 208209 361528 208214 361584
rect 208270 361528 318246 361584
rect 318302 361528 318307 361584
rect 208209 361526 318307 361528
rect 208209 361523 208275 361526
rect 318241 361523 318307 361526
rect 157517 361450 157583 361453
rect 300301 361450 300367 361453
rect 157517 361448 300367 361450
rect 157517 361392 157522 361448
rect 157578 361392 300306 361448
rect 300362 361392 300367 361448
rect 157517 361390 300367 361392
rect 157517 361387 157583 361390
rect 300301 361387 300367 361390
rect 233785 361314 233851 361317
rect 402237 361314 402303 361317
rect 233785 361312 402303 361314
rect 233785 361256 233790 361312
rect 233846 361256 402242 361312
rect 402298 361256 402303 361312
rect 233785 361254 402303 361256
rect 233785 361251 233851 361254
rect 402237 361251 402303 361254
rect 239489 361178 239555 361181
rect 525241 361178 525307 361181
rect 239489 361176 525307 361178
rect 239489 361120 239494 361176
rect 239550 361120 525246 361176
rect 525302 361120 525307 361176
rect 239489 361118 525307 361120
rect 239489 361115 239555 361118
rect 525241 361115 525307 361118
rect 239438 360980 239444 361044
rect 239508 361042 239514 361044
rect 580574 361042 580580 361044
rect 239508 360982 580580 361042
rect 239508 360980 239514 360982
rect 580574 360980 580580 360982
rect 580644 360980 580650 361044
rect 43662 360844 43668 360908
rect 43732 360906 43738 360908
rect 501045 360906 501111 360909
rect 43732 360904 501111 360906
rect 43732 360848 501050 360904
rect 501106 360848 501111 360904
rect 43732 360846 501111 360848
rect 43732 360844 43738 360846
rect 501045 360843 501111 360846
rect 251909 360770 251975 360773
rect 350441 360770 350507 360773
rect 251909 360768 350507 360770
rect 251909 360712 251914 360768
rect 251970 360712 350446 360768
rect 350502 360712 350507 360768
rect 251909 360710 350507 360712
rect 251909 360707 251975 360710
rect 350441 360707 350507 360710
rect 467833 360226 467899 360229
rect 473261 360226 473327 360229
rect 467833 360224 473327 360226
rect 467833 360168 467838 360224
rect 467894 360168 473266 360224
rect 473322 360168 473327 360224
rect 467833 360166 473327 360168
rect 467833 360163 467899 360166
rect 473261 360163 473327 360166
rect 248505 360090 248571 360093
rect 426709 360090 426775 360093
rect 248505 360088 426775 360090
rect 248505 360032 248510 360088
rect 248566 360032 426714 360088
rect 426770 360032 426775 360088
rect 248505 360030 426775 360032
rect 248505 360027 248571 360030
rect 426709 360027 426775 360030
rect 249425 359954 249491 359957
rect 428457 359954 428523 359957
rect 249425 359952 428523 359954
rect 249425 359896 249430 359952
rect 249486 359896 428462 359952
rect 428518 359896 428523 359952
rect 249425 359894 428523 359896
rect 249425 359891 249491 359894
rect 428457 359891 428523 359894
rect 252185 359818 252251 359821
rect 262949 359818 263015 359821
rect 431953 359818 432019 359821
rect 252185 359816 262874 359818
rect 252185 359760 252190 359816
rect 252246 359760 262874 359816
rect 252185 359758 262874 359760
rect 252185 359755 252251 359758
rect 77109 359682 77175 359685
rect 252369 359682 252435 359685
rect 77109 359680 252435 359682
rect 77109 359624 77114 359680
rect 77170 359624 252374 359680
rect 252430 359624 252435 359680
rect 77109 359622 252435 359624
rect 77109 359619 77175 359622
rect 252369 359619 252435 359622
rect 252645 359682 252711 359685
rect 262673 359682 262739 359685
rect 252645 359680 262739 359682
rect 252645 359624 252650 359680
rect 252706 359624 262678 359680
rect 262734 359624 262739 359680
rect 252645 359622 262739 359624
rect 262814 359682 262874 359758
rect 262949 359816 432019 359818
rect 262949 359760 262954 359816
rect 263010 359760 431958 359816
rect 432014 359760 432019 359816
rect 262949 359758 432019 359760
rect 262949 359755 263015 359758
rect 431953 359755 432019 359758
rect 433701 359682 433767 359685
rect 262814 359680 433767 359682
rect 262814 359624 433706 359680
rect 433762 359624 433767 359680
rect 262814 359622 433767 359624
rect 252645 359619 252711 359622
rect 262673 359619 262739 359622
rect 433701 359619 433767 359622
rect 242985 359546 243051 359549
rect 482645 359546 482711 359549
rect 242985 359544 482711 359546
rect 242985 359488 242990 359544
rect 243046 359488 482650 359544
rect 482706 359488 482711 359544
rect 242985 359486 482711 359488
rect 242985 359483 243051 359486
rect 482645 359483 482711 359486
rect 232865 359410 232931 359413
rect 365529 359410 365595 359413
rect 232865 359408 365595 359410
rect 232865 359352 232870 359408
rect 232926 359352 365534 359408
rect 365590 359352 365595 359408
rect 232865 359350 365595 359352
rect 232865 359347 232931 359350
rect 365529 359347 365595 359350
rect 421557 359410 421623 359413
rect 480897 359410 480963 359413
rect 421557 359408 480963 359410
rect 421557 359352 421562 359408
rect 421618 359352 480902 359408
rect 480958 359352 480963 359408
rect 421557 359350 480963 359352
rect 421557 359347 421623 359350
rect 480897 359347 480963 359350
rect 247585 359274 247651 359277
rect 424961 359274 425027 359277
rect 247585 359272 425027 359274
rect 247585 359216 247590 359272
rect 247646 359216 424966 359272
rect 425022 359216 425027 359272
rect 247585 359214 425027 359216
rect 247585 359211 247651 359214
rect 424961 359211 425027 359214
rect 82353 359138 82419 359141
rect 252461 359138 252527 359141
rect 82353 359136 252527 359138
rect 82353 359080 82358 359136
rect 82414 359080 252466 359136
rect 252522 359080 252527 359136
rect 82353 359078 252527 359080
rect 82353 359075 82419 359078
rect 252461 359075 252527 359078
rect 251265 359002 251331 359005
rect 252645 359002 252711 359005
rect 251265 359000 252711 359002
rect 251265 358944 251270 359000
rect 251326 358944 252650 359000
rect 252706 358944 252711 359000
rect 251265 358942 252711 358944
rect 251265 358939 251331 358942
rect 252645 358939 252711 358942
rect 4061 358730 4127 358733
rect 271781 358730 271847 358733
rect 4061 358728 271847 358730
rect 4061 358672 4066 358728
rect 4122 358672 271786 358728
rect 271842 358672 271847 358728
rect 4061 358670 271847 358672
rect 4061 358667 4127 358670
rect 271781 358667 271847 358670
rect 246757 358594 246823 358597
rect 423213 358594 423279 358597
rect 246757 358592 423279 358594
rect -960 358458 480 358548
rect 246757 358536 246762 358592
rect 246818 358536 423218 358592
rect 423274 358536 423279 358592
rect 246757 358534 423279 358536
rect 246757 358531 246823 358534
rect 423213 358531 423279 358534
rect 271781 358458 271847 358461
rect -960 358456 271847 358458
rect -960 358400 271786 358456
rect 271842 358400 271847 358456
rect -960 358398 271847 358400
rect -960 358308 480 358398
rect 271781 358395 271847 358398
rect 269665 358322 269731 358325
rect 466913 358322 466979 358325
rect 269665 358320 466979 358322
rect 269665 358264 269670 358320
rect 269726 358264 466918 358320
rect 466974 358264 466979 358320
rect 269665 358262 466979 358264
rect 269665 358259 269731 358262
rect 466913 358259 466979 358262
rect 270585 358186 270651 358189
rect 468661 358186 468727 358189
rect 270585 358184 468727 358186
rect 270585 358128 270590 358184
rect 270646 358128 468666 358184
rect 468722 358128 468727 358184
rect 270585 358126 468727 358128
rect 270585 358123 270651 358126
rect 468661 358123 468727 358126
rect 271505 358050 271571 358053
rect 470409 358050 470475 358053
rect 271505 358048 470475 358050
rect 271505 357992 271510 358048
rect 271566 357992 470414 358048
rect 470470 357992 470475 358048
rect 271505 357990 470475 357992
rect 271505 357987 271571 357990
rect 470409 357987 470475 357990
rect 245745 357914 245811 357917
rect 421465 357914 421531 357917
rect 245745 357912 421531 357914
rect 245745 357856 245750 357912
rect 245806 357856 421470 357912
rect 421526 357856 421531 357912
rect 245745 357854 421531 357856
rect 245745 357851 245811 357854
rect 421465 357851 421531 357854
rect 268745 357778 268811 357781
rect 403617 357778 403683 357781
rect 268745 357776 403683 357778
rect 268745 357720 268750 357776
rect 268806 357720 403622 357776
rect 403678 357720 403683 357776
rect 268745 357718 403683 357720
rect 268745 357715 268811 357718
rect 403617 357715 403683 357718
rect 246665 357642 246731 357645
rect 280981 357642 281047 357645
rect 246665 357640 281047 357642
rect 246665 357584 246670 357640
rect 246726 357584 280986 357640
rect 281042 357584 281047 357640
rect 246665 357582 281047 357584
rect 246665 357579 246731 357582
rect 280981 357579 281047 357582
rect 282913 357508 282979 357509
rect 282862 357444 282868 357508
rect 282932 357506 282979 357508
rect 282932 357504 283024 357506
rect 282974 357448 283024 357504
rect 282932 357446 283024 357448
rect 282932 357444 282979 357446
rect 282913 357443 282979 357444
rect 254945 357370 255011 357373
rect 438945 357370 439011 357373
rect 254945 357368 439011 357370
rect 254945 357312 254950 357368
rect 255006 357312 438950 357368
rect 439006 357312 439011 357368
rect 254945 357310 439011 357312
rect 254945 357307 255011 357310
rect 438945 357307 439011 357310
rect 255865 357234 255931 357237
rect 440693 357234 440759 357237
rect 255865 357232 440759 357234
rect 255865 357176 255870 357232
rect 255926 357176 440698 357232
rect 440754 357176 440759 357232
rect 255865 357174 440759 357176
rect 255865 357171 255931 357174
rect 440693 357171 440759 357174
rect 256785 357098 256851 357101
rect 442441 357098 442507 357101
rect 256785 357096 442507 357098
rect 256785 357040 256790 357096
rect 256846 357040 442446 357096
rect 442502 357040 442507 357096
rect 256785 357038 442507 357040
rect 256785 357035 256851 357038
rect 442441 357035 442507 357038
rect 257705 356962 257771 356965
rect 444189 356962 444255 356965
rect 257705 356960 444255 356962
rect 257705 356904 257710 356960
rect 257766 356904 444194 356960
rect 444250 356904 444255 356960
rect 257705 356902 444255 356904
rect 257705 356899 257771 356902
rect 444189 356899 444255 356902
rect 258625 356826 258691 356829
rect 445937 356826 446003 356829
rect 258625 356824 446003 356826
rect 258625 356768 258630 356824
rect 258686 356768 445942 356824
rect 445998 356768 446003 356824
rect 258625 356766 446003 356768
rect 258625 356763 258691 356766
rect 445937 356763 446003 356766
rect 259545 356690 259611 356693
rect 447685 356690 447751 356693
rect 259545 356688 447751 356690
rect 259545 356632 259550 356688
rect 259606 356632 447690 356688
rect 447746 356632 447751 356688
rect 259545 356630 447751 356632
rect 259545 356627 259611 356630
rect 447685 356627 447751 356630
rect 254025 356554 254091 356557
rect 437197 356554 437263 356557
rect 254025 356552 437263 356554
rect 254025 356496 254030 356552
rect 254086 356496 437202 356552
rect 437258 356496 437263 356552
rect 254025 356494 437263 356496
rect 254025 356491 254091 356494
rect 437197 356491 437263 356494
rect 3366 355948 3372 356012
rect 3436 356010 3442 356012
rect 238385 356010 238451 356013
rect 3436 356008 238451 356010
rect 3436 355952 238390 356008
rect 238446 355952 238451 356008
rect 3436 355950 238451 355952
rect 3436 355948 3442 355950
rect 238385 355947 238451 355950
rect 276381 356010 276447 356013
rect 358445 356010 358511 356013
rect 276381 356008 358511 356010
rect 276381 355952 276386 356008
rect 276442 355952 358450 356008
rect 358506 355952 358511 356008
rect 276381 355950 358511 355952
rect 276381 355947 276447 355950
rect 358445 355947 358511 355950
rect 460933 356010 460999 356013
rect 467833 356010 467899 356013
rect 460933 356008 467899 356010
rect 460933 355952 460938 356008
rect 460994 355952 467838 356008
rect 467894 355952 467899 356008
rect 460933 355950 467899 355952
rect 460933 355947 460999 355950
rect 467833 355947 467899 355950
rect 529933 356010 529999 356013
rect 530526 356010 530532 356012
rect 529933 356008 530532 356010
rect 529933 355952 529938 356008
rect 529994 355952 530532 356008
rect 529933 355950 530532 355952
rect 529933 355947 529999 355950
rect 530526 355948 530532 355950
rect 530596 355948 530602 356012
rect 532693 356010 532759 356013
rect 533286 356010 533292 356012
rect 532693 356008 533292 356010
rect 532693 355952 532698 356008
rect 532754 355952 533292 356008
rect 532693 355950 533292 355952
rect 532693 355947 532759 355950
rect 533286 355948 533292 355950
rect 533356 355948 533362 356012
rect 534073 356010 534139 356013
rect 534574 356010 534580 356012
rect 534073 356008 534580 356010
rect 534073 355952 534078 356008
rect 534134 355952 534580 356008
rect 534073 355950 534580 355952
rect 534073 355947 534139 355950
rect 534574 355948 534580 355950
rect 534644 355948 534650 356012
rect 233693 355874 233759 355877
rect 407481 355874 407547 355877
rect 233693 355872 407547 355874
rect 233693 355816 233698 355872
rect 233754 355816 407486 355872
rect 407542 355816 407547 355872
rect 233693 355814 407547 355816
rect 233693 355811 233759 355814
rect 407481 355811 407547 355814
rect 267825 355738 267891 355741
rect 463417 355738 463483 355741
rect 267825 355736 463483 355738
rect 267825 355680 267830 355736
rect 267886 355680 463422 355736
rect 463478 355680 463483 355736
rect 267825 355678 463483 355680
rect 267825 355675 267891 355678
rect 463417 355675 463483 355678
rect 71865 355602 71931 355605
rect 287697 355602 287763 355605
rect 71865 355600 287763 355602
rect 71865 355544 71870 355600
rect 71926 355544 287702 355600
rect 287758 355544 287763 355600
rect 71865 355542 287763 355544
rect 71865 355539 71931 355542
rect 287697 355539 287763 355542
rect 238201 355466 238267 355469
rect 526621 355466 526687 355469
rect 238201 355464 526687 355466
rect 238201 355408 238206 355464
rect 238262 355408 526626 355464
rect 526682 355408 526687 355464
rect 238201 355406 526687 355408
rect 238201 355403 238267 355406
rect 526621 355403 526687 355406
rect 239397 355330 239463 355333
rect 532141 355330 532207 355333
rect 239397 355328 532207 355330
rect 239397 355272 239402 355328
rect 239458 355272 532146 355328
rect 532202 355272 532207 355328
rect 239397 355270 532207 355272
rect 239397 355267 239463 355270
rect 532141 355267 532207 355270
rect 235073 355194 235139 355197
rect 372521 355194 372587 355197
rect 235073 355192 372587 355194
rect 235073 355136 235078 355192
rect 235134 355136 372526 355192
rect 372582 355136 372587 355192
rect 235073 355134 372587 355136
rect 235073 355131 235139 355134
rect 372521 355131 372587 355134
rect 237097 355058 237163 355061
rect 276013 355058 276079 355061
rect 284293 355060 284359 355061
rect 284293 355058 284340 355060
rect 237097 355056 276079 355058
rect 237097 355000 237102 355056
rect 237158 355000 276018 355056
rect 276074 355000 276079 355056
rect 237097 354998 276079 355000
rect 284248 355056 284340 355058
rect 284248 355000 284298 355056
rect 284248 354998 284340 355000
rect 237097 354995 237163 354998
rect 276013 354995 276079 354998
rect 284293 354996 284340 354998
rect 284404 354996 284410 355060
rect 284293 354995 284359 354996
rect 238109 354922 238175 354925
rect 269021 354922 269087 354925
rect 238109 354920 269087 354922
rect 238109 354864 238114 354920
rect 238170 354864 269026 354920
rect 269082 354864 269087 354920
rect 238109 354862 269087 354864
rect 238109 354859 238175 354862
rect 269021 354859 269087 354862
rect 31150 354588 31156 354652
rect 31220 354650 31226 354652
rect 239397 354650 239463 354653
rect 31220 354648 239463 354650
rect 31220 354592 239402 354648
rect 239458 354592 239463 354648
rect 31220 354590 239463 354592
rect 31220 354588 31226 354590
rect 239397 354587 239463 354590
rect 31385 354514 31451 354517
rect 237005 354514 237071 354517
rect 31385 354512 237071 354514
rect 31385 354456 31390 354512
rect 31446 354456 237010 354512
rect 237066 354456 237071 354512
rect 31385 354454 237071 354456
rect 31385 354451 31451 354454
rect 237005 354451 237071 354454
rect 31017 354378 31083 354381
rect 237097 354378 237163 354381
rect 31017 354376 237163 354378
rect 31017 354320 31022 354376
rect 31078 354320 237102 354376
rect 237158 354320 237163 354376
rect 31017 354318 237163 354320
rect 31017 354315 31083 354318
rect 237097 354315 237163 354318
rect 239673 354378 239739 354381
rect 504214 354378 504220 354380
rect 239673 354376 504220 354378
rect 239673 354320 239678 354376
rect 239734 354320 504220 354376
rect 239673 354318 504220 354320
rect 239673 354315 239739 354318
rect 504214 354316 504220 354318
rect 504284 354316 504290 354380
rect 236637 354242 236703 354245
rect 506974 354242 506980 354244
rect 236637 354240 506980 354242
rect 236637 354184 236642 354240
rect 236698 354184 506980 354240
rect 236637 354182 506980 354184
rect 236637 354179 236703 354182
rect 506974 354180 506980 354182
rect 507044 354180 507050 354244
rect 236545 354106 236611 354109
rect 508681 354106 508747 354109
rect 236545 354104 508747 354106
rect 236545 354048 236550 354104
rect 236606 354048 508686 354104
rect 508742 354048 508747 354104
rect 236545 354046 508747 354048
rect 236545 354043 236611 354046
rect 508681 354043 508747 354046
rect 3918 353908 3924 353972
rect 3988 353970 3994 353972
rect 283046 353970 283052 353972
rect 3988 353910 283052 353970
rect 3988 353908 3994 353910
rect 283046 353908 283052 353910
rect 283116 353908 283122 353972
rect 235758 353772 235764 353836
rect 235828 353834 235834 353836
rect 409229 353834 409295 353837
rect 235828 353832 409295 353834
rect 235828 353776 409234 353832
rect 409290 353776 409295 353832
rect 235828 353774 409295 353776
rect 235828 353772 235834 353774
rect 409229 353771 409295 353774
rect 235257 353698 235323 353701
rect 374269 353698 374335 353701
rect 235257 353696 374335 353698
rect 235257 353640 235262 353696
rect 235318 353640 374274 353696
rect 374330 353640 374335 353696
rect 235257 353638 374335 353640
rect 235257 353635 235323 353638
rect 374269 353635 374335 353638
rect 231158 353500 231164 353564
rect 231228 353562 231234 353564
rect 285806 353562 285812 353564
rect 231228 353502 285812 353562
rect 231228 353500 231234 353502
rect 285806 353500 285812 353502
rect 285876 353500 285882 353564
rect 239254 353364 239260 353428
rect 239324 353426 239330 353428
rect 240041 353426 240107 353429
rect 239324 353424 240107 353426
rect 239324 353368 240046 353424
rect 240102 353368 240107 353424
rect 239324 353366 240107 353368
rect 239324 353364 239330 353366
rect 240041 353363 240107 353366
rect 43069 353290 43135 353293
rect 235349 353290 235415 353293
rect 43069 353288 235415 353290
rect 43069 353232 43074 353288
rect 43130 353232 235354 353288
rect 235410 353232 235415 353288
rect 43069 353230 235415 353232
rect 43069 353227 43135 353230
rect 235349 353227 235415 353230
rect 199469 353154 199535 353157
rect 329097 353154 329163 353157
rect 199469 353152 329163 353154
rect 199469 353096 199474 353152
rect 199530 353096 329102 353152
rect 329158 353096 329163 353152
rect 199469 353094 329163 353096
rect 199469 353091 199535 353094
rect 329097 353091 329163 353094
rect 148777 353018 148843 353021
rect 301497 353018 301563 353021
rect 148777 353016 301563 353018
rect 148777 352960 148782 353016
rect 148838 352960 301502 353016
rect 301558 352960 301563 353016
rect 148777 352958 301563 352960
rect 148777 352955 148843 352958
rect 301497 352955 301563 352958
rect 235073 352882 235139 352885
rect 388253 352882 388319 352885
rect 235073 352880 388319 352882
rect 235073 352824 235078 352880
rect 235134 352824 388258 352880
rect 388314 352824 388319 352880
rect 235073 352822 388319 352824
rect 235073 352819 235139 352822
rect 388253 352819 388319 352822
rect 105077 352746 105143 352749
rect 289445 352746 289511 352749
rect 105077 352744 289511 352746
rect 105077 352688 105082 352744
rect 105138 352688 289450 352744
rect 289506 352688 289511 352744
rect 105077 352686 289511 352688
rect 105077 352683 105143 352686
rect 289445 352683 289511 352686
rect 401961 352746 402027 352749
rect 497457 352746 497523 352749
rect 401961 352744 497523 352746
rect 401961 352688 401966 352744
rect 402022 352688 497462 352744
rect 497518 352688 497523 352744
rect 401961 352686 497523 352688
rect 401961 352683 402027 352686
rect 497457 352683 497523 352686
rect 50838 352548 50844 352612
rect 50908 352610 50914 352612
rect 347589 352610 347655 352613
rect 421557 352610 421623 352613
rect 50908 352608 347655 352610
rect 50908 352552 347594 352608
rect 347650 352552 347655 352608
rect 50908 352550 347655 352552
rect 50908 352548 50914 352550
rect 347589 352547 347655 352550
rect 373950 352608 421623 352610
rect 373950 352552 421562 352608
rect 421618 352552 421623 352608
rect 373950 352550 421623 352552
rect 230933 352474 230999 352477
rect 296253 352474 296319 352477
rect 230933 352472 296319 352474
rect 230933 352416 230938 352472
rect 230994 352416 296258 352472
rect 296314 352416 296319 352472
rect 230933 352414 296319 352416
rect 230933 352411 230999 352414
rect 296253 352411 296319 352414
rect 373950 351933 374010 352550
rect 421557 352547 421623 352550
rect 457897 352610 457963 352613
rect 471237 352610 471303 352613
rect 457897 352608 471303 352610
rect 457897 352552 457902 352608
rect 457958 352552 471242 352608
rect 471298 352552 471303 352608
rect 457897 352550 471303 352552
rect 457897 352547 457963 352550
rect 471237 352547 471303 352550
rect 429929 352066 429995 352069
rect 431217 352066 431283 352069
rect 429929 352064 431283 352066
rect 429929 352008 429934 352064
rect 429990 352008 431222 352064
rect 431278 352008 431283 352064
rect 429929 352006 431283 352008
rect 429929 352003 429995 352006
rect 431217 352003 431283 352006
rect 224861 351930 224927 351933
rect 283097 351930 283163 351933
rect 224861 351928 283163 351930
rect 224861 351872 224866 351928
rect 224922 351872 283102 351928
rect 283158 351872 283163 351928
rect 224861 351870 283163 351872
rect 224861 351867 224927 351870
rect 283097 351867 283163 351870
rect 358721 351930 358787 351933
rect 373950 351930 374059 351933
rect 358721 351928 374059 351930
rect 358721 351872 358726 351928
rect 358782 351872 373998 351928
rect 374054 351872 374059 351928
rect 358721 351870 374059 351872
rect 358721 351867 358787 351870
rect 373993 351867 374059 351870
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 75361 351794 75427 351797
rect 222101 351794 222167 351797
rect 75361 351792 222167 351794
rect 75361 351736 75366 351792
rect 75422 351736 222106 351792
rect 222162 351736 222167 351792
rect 583520 351780 584960 351870
rect 75361 351734 222167 351736
rect 75361 351731 75427 351734
rect 222101 351731 222167 351734
rect 112069 351658 112135 351661
rect 224217 351658 224283 351661
rect 112069 351656 224283 351658
rect 112069 351600 112074 351656
rect 112130 351600 224222 351656
rect 224278 351600 224283 351656
rect 112069 351598 224283 351600
rect 112069 351595 112135 351598
rect 224217 351595 224283 351598
rect 224677 351522 224743 351525
rect 287145 351522 287211 351525
rect 224677 351520 287211 351522
rect 224677 351464 224682 351520
rect 224738 351464 287150 351520
rect 287206 351464 287211 351520
rect 224677 351462 287211 351464
rect 224677 351459 224743 351462
rect 287145 351459 287211 351462
rect 222009 351386 222075 351389
rect 280429 351386 280495 351389
rect 222009 351384 280495 351386
rect 222009 351328 222014 351384
rect 222070 351328 280434 351384
rect 280490 351328 280495 351384
rect 222009 351326 280495 351328
rect 222009 351323 222075 351326
rect 280429 351323 280495 351326
rect 201217 351250 201283 351253
rect 308581 351250 308647 351253
rect 201217 351248 308647 351250
rect 201217 351192 201222 351248
rect 201278 351192 308586 351248
rect 308642 351192 308647 351248
rect 201217 351190 308647 351192
rect 201217 351187 201283 351190
rect 308581 351187 308647 351190
rect 229921 351116 229987 351117
rect 229870 351114 229876 351116
rect 229830 351054 229876 351114
rect 229940 351112 229987 351116
rect 229982 351056 229987 351112
rect 229870 351052 229876 351054
rect 229940 351052 229987 351056
rect 229921 351051 229987 351052
rect 282821 351114 282887 351117
rect 539685 351114 539751 351117
rect 282821 351112 539751 351114
rect 282821 351056 282826 351112
rect 282882 351056 539690 351112
rect 539746 351056 539751 351112
rect 282821 351054 539751 351056
rect 282821 351051 282887 351054
rect 539685 351051 539751 351054
rect 218789 350978 218855 350981
rect 304993 350978 305059 350981
rect 218789 350976 305059 350978
rect 218789 350920 218794 350976
rect 218850 350920 304998 350976
rect 305054 350920 305059 350976
rect 218789 350918 305059 350920
rect 218789 350915 218855 350918
rect 304993 350915 305059 350918
rect 218973 350842 219039 350845
rect 306373 350842 306439 350845
rect 218973 350840 306439 350842
rect 218973 350784 218978 350840
rect 219034 350784 306378 350840
rect 306434 350784 306439 350840
rect 218973 350782 306439 350784
rect 218973 350779 219039 350782
rect 306373 350779 306439 350782
rect 211797 350706 211863 350709
rect 302601 350706 302667 350709
rect 211797 350704 302667 350706
rect 211797 350648 211802 350704
rect 211858 350648 302606 350704
rect 302662 350648 302667 350704
rect 211797 350646 302667 350648
rect 211797 350643 211863 350646
rect 302601 350643 302667 350646
rect 476113 350706 476179 350709
rect 479517 350706 479583 350709
rect 476113 350704 479583 350706
rect 476113 350648 476118 350704
rect 476174 350648 479522 350704
rect 479578 350648 479583 350704
rect 476113 350646 479583 350648
rect 476113 350643 476179 350646
rect 479517 350643 479583 350646
rect 94497 350570 94563 350573
rect 95877 350570 95943 350573
rect 94497 350568 95943 350570
rect 94497 350512 94502 350568
rect 94558 350512 95882 350568
rect 95938 350512 95943 350568
rect 94497 350510 95943 350512
rect 94497 350507 94563 350510
rect 95877 350507 95943 350510
rect 209037 350570 209103 350573
rect 301129 350570 301195 350573
rect 209037 350568 301195 350570
rect 209037 350512 209042 350568
rect 209098 350512 301134 350568
rect 301190 350512 301195 350568
rect 209037 350510 301195 350512
rect 209037 350507 209103 350510
rect 301129 350507 301195 350510
rect 30097 350434 30163 350437
rect 226333 350434 226399 350437
rect 30097 350432 226399 350434
rect 30097 350376 30102 350432
rect 30158 350376 226338 350432
rect 226394 350376 226399 350432
rect 30097 350374 226399 350376
rect 30097 350371 30163 350374
rect 226333 350371 226399 350374
rect 222193 350162 222259 350165
rect 315481 350162 315547 350165
rect 222193 350160 315547 350162
rect 222193 350104 222198 350160
rect 222254 350104 315486 350160
rect 315542 350104 315547 350160
rect 222193 350102 315547 350104
rect 222193 350099 222259 350102
rect 315481 350099 315547 350102
rect 174997 350026 175063 350029
rect 293401 350026 293467 350029
rect 174997 350024 293467 350026
rect 174997 349968 175002 350024
rect 175058 349968 293406 350024
rect 293462 349968 293467 350024
rect 174997 349966 293467 349968
rect 174997 349963 175063 349966
rect 293401 349963 293467 349966
rect 126053 349890 126119 349893
rect 300209 349890 300275 349893
rect 126053 349888 300275 349890
rect 126053 349832 126058 349888
rect 126114 349832 300214 349888
rect 300270 349832 300275 349888
rect 126053 349830 300275 349832
rect 126053 349827 126119 349830
rect 300209 349827 300275 349830
rect 346209 349890 346275 349893
rect 460841 349890 460907 349893
rect 346209 349888 460907 349890
rect 346209 349832 346214 349888
rect 346270 349832 460846 349888
rect 460902 349832 460907 349888
rect 346209 349830 460907 349832
rect 346209 349827 346275 349830
rect 460841 349827 460907 349830
rect 99833 349754 99899 349757
rect 287881 349754 287947 349757
rect 99833 349752 287947 349754
rect 99833 349696 99838 349752
rect 99894 349696 287886 349752
rect 287942 349696 287947 349752
rect 99833 349694 287947 349696
rect 99833 349691 99899 349694
rect 287881 349691 287947 349694
rect 353293 349754 353359 349757
rect 476113 349754 476179 349757
rect 353293 349752 476179 349754
rect 353293 349696 353298 349752
rect 353354 349696 476118 349752
rect 476174 349696 476179 349752
rect 353293 349694 476179 349696
rect 353293 349691 353359 349694
rect 476113 349691 476179 349694
rect 227345 349618 227411 349621
rect 288525 349618 288591 349621
rect 227345 349616 288591 349618
rect 227345 349560 227350 349616
rect 227406 349560 288530 349616
rect 288586 349560 288591 349616
rect 227345 349558 288591 349560
rect 227345 349555 227411 349558
rect 288525 349555 288591 349558
rect 227161 349482 227227 349485
rect 284753 349482 284819 349485
rect 227161 349480 284819 349482
rect 227161 349424 227166 349480
rect 227222 349424 284758 349480
rect 284814 349424 284819 349480
rect 227161 349422 284819 349424
rect 227161 349419 227227 349422
rect 284753 349419 284819 349422
rect 226977 349346 227043 349349
rect 287053 349346 287119 349349
rect 226977 349344 287119 349346
rect 226977 349288 226982 349344
rect 227038 349288 287058 349344
rect 287114 349288 287119 349344
rect 226977 349286 287119 349288
rect 226977 349283 227043 349286
rect 287053 349283 287119 349286
rect 234981 349210 235047 349213
rect 298093 349212 298159 349213
rect 235206 349210 235212 349212
rect 234981 349208 235212 349210
rect 234981 349152 234986 349208
rect 235042 349152 235212 349208
rect 234981 349150 235212 349152
rect 234981 349147 235047 349150
rect 235206 349148 235212 349150
rect 235276 349148 235282 349212
rect 298093 349210 298140 349212
rect 298048 349208 298140 349210
rect 298048 349152 298098 349208
rect 298048 349150 298140 349152
rect 298093 349148 298140 349150
rect 298204 349148 298210 349212
rect 298093 349147 298159 349148
rect 212257 349074 212323 349077
rect 249701 349074 249767 349077
rect 212257 349072 249767 349074
rect 212257 349016 212262 349072
rect 212318 349016 249706 349072
rect 249762 349016 249767 349072
rect 212257 349014 249767 349016
rect 212257 349011 212323 349014
rect 249701 349011 249767 349014
rect 282913 349074 282979 349077
rect 361614 349074 361620 349076
rect 282913 349072 361620 349074
rect 282913 349016 282918 349072
rect 282974 349016 361620 349072
rect 282913 349014 361620 349016
rect 282913 349011 282979 349014
rect 361614 349012 361620 349014
rect 361684 349012 361690 349076
rect 94589 348938 94655 348941
rect 220721 348938 220787 348941
rect 94589 348936 220787 348938
rect 94589 348880 94594 348936
rect 94650 348880 220726 348936
rect 220782 348880 220787 348936
rect 94589 348878 220787 348880
rect 94589 348875 94655 348878
rect 220721 348875 220787 348878
rect 284293 348938 284359 348941
rect 362902 348938 362908 348940
rect 284293 348936 362908 348938
rect 284293 348880 284298 348936
rect 284354 348880 362908 348936
rect 284293 348878 362908 348880
rect 284293 348875 284359 348878
rect 362902 348876 362908 348878
rect 362972 348876 362978 348940
rect 113817 348802 113883 348805
rect 222101 348802 222167 348805
rect 113817 348800 222167 348802
rect 113817 348744 113822 348800
rect 113878 348744 222106 348800
rect 222162 348744 222167 348800
rect 113817 348742 222167 348744
rect 113817 348739 113883 348742
rect 222101 348739 222167 348742
rect 258901 348802 258967 348805
rect 259637 348802 259703 348805
rect 258901 348800 259703 348802
rect 258901 348744 258906 348800
rect 258962 348744 259642 348800
rect 259698 348744 259703 348800
rect 258901 348742 259703 348744
rect 258901 348739 258967 348742
rect 259637 348739 259703 348742
rect 150525 348666 150591 348669
rect 224217 348666 224283 348669
rect 150525 348664 224283 348666
rect 150525 348608 150530 348664
rect 150586 348608 224222 348664
rect 224278 348608 224283 348664
rect 150525 348606 224283 348608
rect 150525 348603 150591 348606
rect 224217 348603 224283 348606
rect 227069 348666 227135 348669
rect 283281 348666 283347 348669
rect 227069 348664 283347 348666
rect 227069 348608 227074 348664
rect 227130 348608 283286 348664
rect 283342 348608 283347 348664
rect 227069 348606 283347 348608
rect 227069 348603 227135 348606
rect 283281 348603 283347 348606
rect 187233 348530 187299 348533
rect 226425 348530 226491 348533
rect 187233 348528 226491 348530
rect 187233 348472 187238 348528
rect 187294 348472 226430 348528
rect 226486 348472 226491 348528
rect 187233 348470 226491 348472
rect 187233 348467 187299 348470
rect 226425 348467 226491 348470
rect 248321 348530 248387 348533
rect 327809 348530 327875 348533
rect 248321 348528 327875 348530
rect 248321 348472 248326 348528
rect 248382 348472 327814 348528
rect 327870 348472 327875 348528
rect 248321 348470 327875 348472
rect 248321 348467 248387 348470
rect 327809 348467 327875 348470
rect 212073 348394 212139 348397
rect 259361 348394 259427 348397
rect 212073 348392 259427 348394
rect 212073 348336 212078 348392
rect 212134 348336 259366 348392
rect 259422 348336 259427 348392
rect 212073 348334 259427 348336
rect 212073 348331 212139 348334
rect 259361 348331 259427 348334
rect 259637 348394 259703 348397
rect 351177 348394 351243 348397
rect 259637 348392 351243 348394
rect 259637 348336 259642 348392
rect 259698 348336 351182 348392
rect 351238 348336 351243 348392
rect 259637 348334 351243 348336
rect 259637 348331 259703 348334
rect 351177 348331 351243 348334
rect 68369 348258 68435 348261
rect 212441 348258 212507 348261
rect 68369 348256 212507 348258
rect 68369 348200 68374 348256
rect 68430 348200 212446 348256
rect 212502 348200 212507 348256
rect 68369 348198 212507 348200
rect 68369 348195 68435 348198
rect 212441 348195 212507 348198
rect 224401 348258 224467 348261
rect 284661 348258 284727 348261
rect 224401 348256 284727 348258
rect 224401 348200 224406 348256
rect 224462 348200 284666 348256
rect 284722 348200 284727 348256
rect 224401 348198 284727 348200
rect 224401 348195 224467 348198
rect 284661 348195 284727 348198
rect 220077 348122 220143 348125
rect 290089 348122 290155 348125
rect 220077 348120 290155 348122
rect 220077 348064 220082 348120
rect 220138 348064 290094 348120
rect 290150 348064 290155 348120
rect 220077 348062 290155 348064
rect 220077 348059 220143 348062
rect 290089 348059 290155 348062
rect 211889 347986 211955 347989
rect 226333 347986 226399 347989
rect 211889 347984 226399 347986
rect 211889 347928 211894 347984
rect 211950 347928 226338 347984
rect 226394 347928 226399 347984
rect 211889 347926 226399 347928
rect 211889 347923 211955 347926
rect 226333 347923 226399 347926
rect 227478 347924 227484 347988
rect 227548 347986 227554 347988
rect 299422 347986 299428 347988
rect 227548 347926 299428 347986
rect 227548 347924 227554 347926
rect 299422 347924 299428 347926
rect 299492 347924 299498 347988
rect 71681 347850 71747 347853
rect 212257 347850 212323 347853
rect 71681 347848 212323 347850
rect 71681 347792 71686 347848
rect 71742 347792 212262 347848
rect 212318 347792 212323 347848
rect 71681 347790 212323 347792
rect 71681 347787 71747 347790
rect 212257 347787 212323 347790
rect 221549 347850 221615 347853
rect 226517 347850 226583 347853
rect 221549 347848 226583 347850
rect 221549 347792 221554 347848
rect 221610 347792 226522 347848
rect 226578 347792 226583 347848
rect 221549 347790 226583 347792
rect 221549 347787 221615 347790
rect 226517 347787 226583 347790
rect 226926 347788 226932 347852
rect 226996 347850 227002 347852
rect 299606 347850 299612 347852
rect 226996 347790 299612 347850
rect 226996 347788 227002 347790
rect 299606 347788 299612 347790
rect 299676 347788 299682 347852
rect 357249 347850 357315 347853
rect 531405 347850 531471 347853
rect 357249 347848 531471 347850
rect 357249 347792 357254 347848
rect 357310 347792 531410 347848
rect 531466 347792 531471 347848
rect 357249 347790 531471 347792
rect 357249 347787 357315 347790
rect 531405 347787 531471 347790
rect 85849 347714 85915 347717
rect 220721 347714 220787 347717
rect 85849 347712 220787 347714
rect 85849 347656 85854 347712
rect 85910 347656 220726 347712
rect 220782 347656 220787 347712
rect 85849 347654 220787 347656
rect 85849 347651 85915 347654
rect 220721 347651 220787 347654
rect 98085 347578 98151 347581
rect 223297 347578 223363 347581
rect 98085 347576 223363 347578
rect 98085 347520 98090 347576
rect 98146 347520 223302 347576
rect 223358 347520 223363 347576
rect 98085 347518 223363 347520
rect 98085 347515 98151 347518
rect 223297 347515 223363 347518
rect 223430 347516 223436 347580
rect 223500 347578 223506 347580
rect 288566 347578 288572 347580
rect 223500 347518 288572 347578
rect 223500 347516 223506 347518
rect 288566 347516 288572 347518
rect 288636 347516 288642 347580
rect 124305 347442 124371 347445
rect 225045 347442 225111 347445
rect 124305 347440 225111 347442
rect 124305 347384 124310 347440
rect 124366 347384 225050 347440
rect 225106 347384 225111 347440
rect 124305 347382 225111 347384
rect 124305 347379 124371 347382
rect 225045 347379 225111 347382
rect 267641 347442 267707 347445
rect 300577 347442 300643 347445
rect 267641 347440 300643 347442
rect 267641 347384 267646 347440
rect 267702 347384 300582 347440
rect 300638 347384 300643 347440
rect 267641 347382 300643 347384
rect 267641 347379 267707 347382
rect 300577 347379 300643 347382
rect 220445 347306 220511 347309
rect 283649 347306 283715 347309
rect 220445 347304 283715 347306
rect 220445 347248 220450 347304
rect 220506 347248 283654 347304
rect 283710 347248 283715 347304
rect 220445 347246 283715 347248
rect 220445 347243 220511 347246
rect 283649 347243 283715 347246
rect 218697 347170 218763 347173
rect 285213 347170 285279 347173
rect 218697 347168 285279 347170
rect 218697 347112 218702 347168
rect 218758 347112 285218 347168
rect 285274 347112 285279 347168
rect 218697 347110 285279 347112
rect 218697 347107 218763 347110
rect 285213 347107 285279 347110
rect 337377 347170 337443 347173
rect 353293 347170 353359 347173
rect 337377 347168 353359 347170
rect 337377 347112 337382 347168
rect 337438 347112 353298 347168
rect 353354 347112 353359 347168
rect 337377 347110 353359 347112
rect 337377 347107 337443 347110
rect 353293 347107 353359 347110
rect 173249 347034 173315 347037
rect 224953 347034 225019 347037
rect 173249 347032 225019 347034
rect 173249 346976 173254 347032
rect 173310 346976 224958 347032
rect 225014 346976 225019 347032
rect 173249 346974 225019 346976
rect 173249 346971 173315 346974
rect 224953 346971 225019 346974
rect 225781 347034 225847 347037
rect 243537 347034 243603 347037
rect 225781 347032 243603 347034
rect 225781 346976 225786 347032
rect 225842 346976 243542 347032
rect 243598 346976 243603 347032
rect 225781 346974 243603 346976
rect 225781 346971 225847 346974
rect 243537 346971 243603 346974
rect 244089 347034 244155 347037
rect 359825 347034 359891 347037
rect 244089 347032 359891 347034
rect 244089 346976 244094 347032
rect 244150 346976 359830 347032
rect 359886 346976 359891 347032
rect 244089 346974 359891 346976
rect 244089 346971 244155 346974
rect 359825 346971 359891 346974
rect 224350 346836 224356 346900
rect 224420 346898 224426 346900
rect 278998 346898 279004 346900
rect 224420 346838 279004 346898
rect 224420 346836 224426 346838
rect 278998 346836 279004 346838
rect 279068 346836 279074 346900
rect 227110 346700 227116 346764
rect 227180 346762 227186 346764
rect 291326 346762 291332 346764
rect 227180 346702 291332 346762
rect 227180 346700 227186 346702
rect 291326 346700 291332 346702
rect 291396 346700 291402 346764
rect 214782 346564 214788 346628
rect 214852 346626 214858 346628
rect 224217 346626 224283 346629
rect 214852 346624 224283 346626
rect 214852 346568 224222 346624
rect 224278 346568 224283 346624
rect 214852 346566 224283 346568
rect 214852 346564 214858 346566
rect 224217 346563 224283 346566
rect 48078 346428 48084 346492
rect 48148 346490 48154 346492
rect 266353 346490 266419 346493
rect 48148 346488 266419 346490
rect 48148 346432 266358 346488
rect 266414 346432 266419 346488
rect 48148 346430 266419 346432
rect 48148 346428 48154 346430
rect 266353 346427 266419 346430
rect 84101 346354 84167 346357
rect 220721 346354 220787 346357
rect 84101 346352 220787 346354
rect 84101 346296 84106 346352
rect 84162 346296 220726 346352
rect 220782 346296 220787 346352
rect 84101 346294 220787 346296
rect 84101 346291 84167 346294
rect 220721 346291 220787 346294
rect 220997 346354 221063 346357
rect 220997 346352 223498 346354
rect 220997 346296 221002 346352
rect 221058 346296 223498 346352
rect 220997 346294 223498 346296
rect 220997 346291 221063 346294
rect 87597 346218 87663 346221
rect 223205 346218 223271 346221
rect 87597 346216 223271 346218
rect 87597 346160 87602 346216
rect 87658 346160 223210 346216
rect 223266 346160 223271 346216
rect 87597 346158 223271 346160
rect 87597 346155 87663 346158
rect 223205 346155 223271 346158
rect 101581 346082 101647 346085
rect 223113 346082 223179 346085
rect 101581 346080 223179 346082
rect 101581 346024 101586 346080
rect 101642 346024 223118 346080
rect 223174 346024 223179 346080
rect 101581 346022 223179 346024
rect 223438 346082 223498 346294
rect 226190 346156 226196 346220
rect 226260 346218 226266 346220
rect 290774 346218 290780 346220
rect 226260 346158 290780 346218
rect 226260 346156 226266 346158
rect 290774 346156 290780 346158
rect 290844 346156 290850 346220
rect 274633 346082 274699 346085
rect 295057 346082 295123 346085
rect 503621 346082 503687 346085
rect 223438 346022 229110 346082
rect 101581 346019 101647 346022
rect 223113 346019 223179 346022
rect 220261 345946 220327 345949
rect 220997 345946 221063 345949
rect 220261 345944 221063 345946
rect 220261 345888 220266 345944
rect 220322 345888 221002 345944
rect 221058 345888 221063 345944
rect 220261 345886 221063 345888
rect 220261 345883 220327 345886
rect 220997 345883 221063 345886
rect 223021 345946 223087 345949
rect 229050 345946 229110 346022
rect 274633 346080 295123 346082
rect 274633 346024 274638 346080
rect 274694 346024 295062 346080
rect 295118 346024 295123 346080
rect 274633 346022 295123 346024
rect 274633 346019 274699 346022
rect 295057 346019 295123 346022
rect 499806 346080 503687 346082
rect 499806 346024 503626 346080
rect 503682 346024 503687 346080
rect 499806 346022 503687 346024
rect 253105 345946 253171 345949
rect 223021 345944 223498 345946
rect 223021 345888 223026 345944
rect 223082 345888 223498 345944
rect 223021 345886 223498 345888
rect 229050 345944 253171 345946
rect 229050 345888 253110 345944
rect 253166 345888 253171 345944
rect 229050 345886 253171 345888
rect 223021 345883 223087 345886
rect 138289 345810 138355 345813
rect 223297 345810 223363 345813
rect 138289 345808 223363 345810
rect 138289 345752 138294 345808
rect 138350 345752 223302 345808
rect 223358 345752 223363 345808
rect 138289 345750 223363 345752
rect 223438 345810 223498 345886
rect 253105 345883 253171 345886
rect 260649 345946 260715 345949
rect 292297 345946 292363 345949
rect 260649 345944 292363 345946
rect 260649 345888 260654 345944
rect 260710 345888 292302 345944
rect 292358 345888 292363 345944
rect 260649 345886 292363 345888
rect 260649 345883 260715 345886
rect 292297 345883 292363 345886
rect 244273 345810 244339 345813
rect 223438 345808 244339 345810
rect 223438 345752 244278 345808
rect 244334 345752 244339 345808
rect 223438 345750 244339 345752
rect 138289 345747 138355 345750
rect 223297 345747 223363 345750
rect 244273 345747 244339 345750
rect 253657 345810 253723 345813
rect 286777 345810 286843 345813
rect 253657 345808 286843 345810
rect 253657 345752 253662 345808
rect 253718 345752 286782 345808
rect 286838 345752 286843 345808
rect 253657 345750 286843 345752
rect 253657 345747 253723 345750
rect 286777 345747 286843 345750
rect 360142 345748 360148 345812
rect 360212 345810 360218 345812
rect 360469 345810 360535 345813
rect 360212 345808 360535 345810
rect 360212 345752 360474 345808
rect 360530 345752 360535 345808
rect 360212 345750 360535 345752
rect 360212 345748 360218 345750
rect 360469 345747 360535 345750
rect 499806 345712 499866 346022
rect 503621 346019 503687 346022
rect 217542 345612 217548 345676
rect 217612 345674 217618 345676
rect 274633 345674 274699 345677
rect 217612 345672 274699 345674
rect 217612 345616 274638 345672
rect 274694 345616 274699 345672
rect 217612 345614 274699 345616
rect 217612 345612 217618 345614
rect 274633 345611 274699 345614
rect 280153 345674 280219 345677
rect 280654 345674 280660 345676
rect 280153 345672 280660 345674
rect 280153 345616 280158 345672
rect 280214 345616 280660 345672
rect 280153 345614 280660 345616
rect 280153 345611 280219 345614
rect 280654 345612 280660 345614
rect 280724 345612 280730 345676
rect 284293 345674 284359 345677
rect 284518 345674 284524 345676
rect 284293 345672 284524 345674
rect 284293 345616 284298 345672
rect 284354 345616 284524 345672
rect 284293 345614 284524 345616
rect 284293 345611 284359 345614
rect 284518 345612 284524 345614
rect 284588 345612 284594 345676
rect 188981 345538 189047 345541
rect 226333 345538 226399 345541
rect 188981 345536 226399 345538
rect -960 345402 480 345492
rect 188981 345480 188986 345536
rect 189042 345480 226338 345536
rect 226394 345480 226399 345536
rect 188981 345478 226399 345480
rect 188981 345475 189047 345478
rect 226333 345475 226399 345478
rect 228214 345476 228220 345540
rect 228284 345538 228290 345540
rect 287646 345538 287652 345540
rect 228284 345478 287652 345538
rect 228284 345476 228290 345478
rect 287646 345476 287652 345478
rect 287716 345476 287722 345540
rect 4102 345402 4108 345404
rect -960 345342 4108 345402
rect -960 345252 480 345342
rect 4102 345340 4108 345342
rect 4172 345340 4178 345404
rect 222694 345340 222700 345404
rect 222764 345402 222770 345404
rect 225873 345402 225939 345405
rect 222764 345400 225939 345402
rect 222764 345344 225878 345400
rect 225934 345344 225939 345400
rect 222764 345342 225939 345344
rect 222764 345340 222770 345342
rect 225873 345339 225939 345342
rect 227294 345340 227300 345404
rect 227364 345402 227370 345404
rect 288382 345402 288388 345404
rect 227364 345342 288388 345402
rect 227364 345340 227370 345342
rect 288382 345340 288388 345342
rect 288452 345340 288458 345404
rect 212165 345266 212231 345269
rect 296989 345266 297055 345269
rect 212165 345264 297055 345266
rect 212165 345208 212170 345264
rect 212226 345208 296994 345264
rect 297050 345208 297055 345264
rect 212165 345206 297055 345208
rect 212165 345203 212231 345206
rect 296989 345203 297055 345206
rect 62021 345130 62087 345133
rect 216673 345130 216739 345133
rect 62021 345128 216739 345130
rect 62021 345072 62026 345128
rect 62082 345072 216678 345128
rect 216734 345072 216739 345128
rect 62021 345070 216739 345072
rect 62021 345067 62087 345070
rect 216673 345067 216739 345070
rect 222837 345130 222903 345133
rect 227713 345130 227779 345133
rect 222837 345128 227779 345130
rect 222837 345072 222842 345128
rect 222898 345072 227718 345128
rect 227774 345072 227779 345128
rect 222837 345070 227779 345072
rect 222837 345067 222903 345070
rect 227713 345067 227779 345070
rect 244825 345130 244891 345133
rect 260741 345130 260807 345133
rect 244825 345128 260807 345130
rect 244825 345072 244830 345128
rect 244886 345072 260746 345128
rect 260802 345072 260807 345128
rect 244825 345070 260807 345072
rect 244825 345067 244891 345070
rect 260741 345067 260807 345070
rect 339401 345130 339467 345133
rect 346209 345130 346275 345133
rect 339401 345128 346275 345130
rect 339401 345072 339406 345128
rect 339462 345072 346214 345128
rect 346270 345072 346275 345128
rect 339401 345070 346275 345072
rect 339401 345067 339467 345070
rect 346209 345067 346275 345070
rect 89345 344994 89411 344997
rect 214557 344994 214623 344997
rect 89345 344992 214623 344994
rect 89345 344936 89350 344992
rect 89406 344936 214562 344992
rect 214618 344936 214623 344992
rect 89345 344934 214623 344936
rect 89345 344931 89411 344934
rect 214557 344931 214623 344934
rect 217358 344932 217364 344996
rect 217428 344994 217434 344996
rect 255313 344994 255379 344997
rect 217428 344992 255379 344994
rect 217428 344936 255318 344992
rect 255374 344936 255379 344992
rect 217428 344934 255379 344936
rect 217428 344932 217434 344934
rect 255313 344931 255379 344934
rect 108573 344858 108639 344861
rect 216673 344858 216739 344861
rect 108573 344856 216739 344858
rect 108573 344800 108578 344856
rect 108634 344800 216678 344856
rect 216734 344800 216739 344856
rect 108573 344798 216739 344800
rect 108573 344795 108639 344798
rect 216673 344795 216739 344798
rect 218646 344796 218652 344860
rect 218716 344858 218722 344860
rect 306414 344858 306420 344860
rect 218716 344798 306420 344858
rect 218716 344796 218722 344798
rect 306414 344796 306420 344798
rect 306484 344796 306490 344860
rect 213177 344722 213243 344725
rect 251081 344722 251147 344725
rect 213177 344720 251147 344722
rect 213177 344664 213182 344720
rect 213238 344664 251086 344720
rect 251142 344664 251147 344720
rect 213177 344662 251147 344664
rect 213177 344659 213243 344662
rect 251081 344659 251147 344662
rect 145281 344586 145347 344589
rect 224217 344586 224283 344589
rect 145281 344584 224283 344586
rect 145281 344528 145286 344584
rect 145342 344528 224222 344584
rect 224278 344528 224283 344584
rect 145281 344526 224283 344528
rect 145281 344523 145347 344526
rect 224217 344523 224283 344526
rect 271137 344586 271203 344589
rect 285305 344586 285371 344589
rect 271137 344584 285371 344586
rect 271137 344528 271142 344584
rect 271198 344528 285310 344584
rect 285366 344528 285371 344584
rect 271137 344526 285371 344528
rect 271137 344523 271203 344526
rect 285305 344523 285371 344526
rect 197721 344450 197787 344453
rect 235993 344450 236059 344453
rect 197721 344448 236059 344450
rect 197721 344392 197726 344448
rect 197782 344392 235998 344448
rect 236054 344392 236059 344448
rect 197721 344390 236059 344392
rect 197721 344387 197787 344390
rect 235993 344387 236059 344390
rect 243169 344450 243235 344453
rect 292205 344450 292271 344453
rect 243169 344448 292271 344450
rect 243169 344392 243174 344448
rect 243230 344392 292210 344448
rect 292266 344392 292271 344448
rect 243169 344390 292271 344392
rect 243169 344387 243235 344390
rect 292205 344387 292271 344390
rect 131297 344314 131363 344317
rect 218053 344314 218119 344317
rect 131297 344312 218119 344314
rect 131297 344256 131302 344312
rect 131358 344256 218058 344312
rect 218114 344256 218119 344312
rect 131297 344254 218119 344256
rect 131297 344251 131363 344254
rect 218053 344251 218119 344254
rect 250161 344314 250227 344317
rect 345657 344314 345723 344317
rect 250161 344312 345723 344314
rect 250161 344256 250166 344312
rect 250222 344256 345662 344312
rect 345718 344256 345723 344312
rect 250161 344254 345723 344256
rect 250161 344251 250227 344254
rect 345657 344251 345723 344254
rect 214741 344178 214807 344181
rect 271781 344178 271847 344181
rect 214741 344176 271847 344178
rect 214741 344120 214746 344176
rect 214802 344120 271786 344176
rect 271842 344120 271847 344176
rect 214741 344118 271847 344120
rect 214741 344115 214807 344118
rect 271781 344115 271847 344118
rect 212349 344042 212415 344045
rect 281073 344042 281139 344045
rect 212349 344040 281139 344042
rect 212349 343984 212354 344040
rect 212410 343984 281078 344040
rect 281134 343984 281139 344040
rect 212349 343982 281139 343984
rect 212349 343979 212415 343982
rect 281073 343979 281139 343982
rect 224534 343844 224540 343908
rect 224604 343906 224610 343908
rect 303654 343906 303660 343908
rect 224604 343846 303660 343906
rect 224604 343844 224610 343846
rect 303654 343844 303660 343846
rect 303724 343844 303730 343908
rect 236361 343770 236427 343773
rect 243537 343770 243603 343773
rect 279509 343770 279575 343773
rect 236361 343768 243603 343770
rect 236361 343712 236366 343768
rect 236422 343712 243542 343768
rect 243598 343712 243603 343768
rect 236361 343710 243603 343712
rect 236361 343707 236427 343710
rect 243537 343707 243603 343710
rect 255270 343768 279575 343770
rect 255270 343712 279514 343768
rect 279570 343712 279575 343768
rect 255270 343710 279575 343712
rect 92841 343634 92907 343637
rect 214373 343634 214439 343637
rect 92841 343632 214439 343634
rect 92841 343576 92846 343632
rect 92902 343576 214378 343632
rect 214434 343576 214439 343632
rect 92841 343574 214439 343576
rect 92841 343571 92907 343574
rect 214373 343571 214439 343574
rect 215109 343634 215175 343637
rect 244273 343634 244339 343637
rect 215109 343632 244339 343634
rect 215109 343576 215114 343632
rect 215170 343576 244278 343632
rect 244334 343576 244339 343632
rect 215109 343574 244339 343576
rect 215109 343571 215175 343574
rect 244273 343571 244339 343574
rect 103329 343498 103395 343501
rect 214465 343498 214531 343501
rect 103329 343496 214531 343498
rect 103329 343440 103334 343496
rect 103390 343440 214470 343496
rect 214526 343440 214531 343496
rect 103329 343438 214531 343440
rect 103329 343435 103395 343438
rect 214465 343435 214531 343438
rect 117313 343362 117379 343365
rect 214649 343362 214715 343365
rect 117313 343360 214715 343362
rect 117313 343304 117318 343360
rect 117374 343304 214654 343360
rect 214710 343304 214715 343360
rect 117313 343302 214715 343304
rect 117313 343299 117379 343302
rect 214649 343299 214715 343302
rect 162761 343226 162827 343229
rect 214557 343226 214623 343229
rect 162761 343224 214623 343226
rect 162761 343168 162766 343224
rect 162822 343168 214562 343224
rect 214618 343168 214623 343224
rect 162761 343166 214623 343168
rect 162761 343163 162827 343166
rect 214557 343163 214623 343166
rect 212441 343090 212507 343093
rect 255270 343090 255330 343710
rect 279509 343707 279575 343710
rect 255405 343226 255471 343229
rect 299197 343226 299263 343229
rect 255405 343224 299263 343226
rect 255405 343168 255410 343224
rect 255466 343168 299202 343224
rect 299258 343168 299263 343224
rect 255405 343166 299263 343168
rect 255405 343163 255471 343166
rect 299197 343163 299263 343166
rect 212441 343088 255330 343090
rect 212441 343032 212446 343088
rect 212502 343032 255330 343088
rect 212441 343030 255330 343032
rect 333513 343090 333579 343093
rect 339401 343090 339467 343093
rect 333513 343088 339467 343090
rect 333513 343032 333518 343088
rect 333574 343032 339406 343088
rect 339462 343032 339467 343088
rect 333513 343030 339467 343032
rect 212441 343027 212507 343030
rect 333513 343027 333579 343030
rect 339401 343027 339467 343030
rect 244917 342954 244983 342957
rect 334709 342954 334775 342957
rect 244917 342952 334775 342954
rect 244917 342896 244922 342952
rect 244978 342896 334714 342952
rect 334770 342896 334775 342952
rect 244917 342894 334775 342896
rect 244917 342891 244983 342894
rect 334709 342891 334775 342894
rect 214598 342756 214604 342820
rect 214668 342818 214674 342820
rect 231117 342818 231183 342821
rect 214668 342816 231183 342818
rect 214668 342760 231122 342816
rect 231178 342760 231183 342816
rect 214668 342758 231183 342760
rect 214668 342756 214674 342758
rect 231117 342755 231183 342758
rect 231342 342756 231348 342820
rect 231412 342818 231418 342820
rect 295558 342818 295564 342820
rect 231412 342758 295564 342818
rect 231412 342756 231418 342758
rect 295558 342756 295564 342758
rect 295628 342756 295634 342820
rect 214281 342682 214347 342685
rect 283465 342682 283531 342685
rect 214281 342680 283531 342682
rect 214281 342624 214286 342680
rect 214342 342624 283470 342680
rect 283526 342624 283531 342680
rect 214281 342622 283531 342624
rect 214281 342619 214347 342622
rect 283465 342619 283531 342622
rect 214414 342484 214420 342548
rect 214484 342546 214490 342548
rect 224217 342546 224283 342549
rect 214484 342544 224283 342546
rect 214484 342488 224222 342544
rect 224278 342488 224283 342544
rect 214484 342486 224283 342488
rect 214484 342484 214490 342486
rect 224217 342483 224283 342486
rect 224718 342484 224724 342548
rect 224788 342546 224794 342548
rect 295374 342546 295380 342548
rect 224788 342486 295380 342546
rect 224788 342484 224794 342486
rect 295374 342484 295380 342486
rect 295444 342484 295450 342548
rect 214925 342410 214991 342413
rect 285949 342410 286015 342413
rect 214925 342408 286015 342410
rect 214925 342352 214930 342408
rect 214986 342352 285954 342408
rect 286010 342352 286015 342408
rect 214925 342350 286015 342352
rect 214925 342347 214991 342350
rect 285949 342347 286015 342350
rect 214833 342274 214899 342277
rect 294137 342274 294203 342277
rect 214833 342272 294203 342274
rect 214833 342216 214838 342272
rect 214894 342216 294142 342272
rect 294198 342216 294203 342272
rect 214833 342214 294203 342216
rect 214833 342211 214899 342214
rect 294137 342211 294203 342214
rect 206461 342138 206527 342141
rect 235993 342138 236059 342141
rect 206461 342136 236059 342138
rect 206461 342080 206466 342136
rect 206522 342080 235998 342136
rect 236054 342080 236059 342136
rect 206461 342078 236059 342080
rect 206461 342075 206527 342078
rect 235993 342075 236059 342078
rect 220302 341940 220308 342004
rect 220372 342002 220378 342004
rect 256693 342002 256759 342005
rect 220372 342000 256759 342002
rect 220372 341944 256698 342000
rect 256754 341944 256759 342000
rect 220372 341942 256759 341944
rect 220372 341940 220378 341942
rect 256693 341939 256759 341942
rect 147029 341866 147095 341869
rect 223297 341866 223363 341869
rect 147029 341864 223363 341866
rect 147029 341808 147034 341864
rect 147090 341808 223302 341864
rect 223358 341808 223363 341864
rect 147029 341806 223363 341808
rect 147029 341803 147095 341806
rect 223297 341803 223363 341806
rect 257153 341866 257219 341869
rect 288249 341866 288315 341869
rect 257153 341864 288315 341866
rect 257153 341808 257158 341864
rect 257214 341808 288254 341864
rect 288310 341808 288315 341864
rect 257153 341806 288315 341808
rect 257153 341803 257219 341806
rect 288249 341803 288315 341806
rect 164509 341730 164575 341733
rect 224953 341730 225019 341733
rect 164509 341728 225019 341730
rect 164509 341672 164514 341728
rect 164570 341672 224958 341728
rect 225014 341672 225019 341728
rect 164509 341670 225019 341672
rect 164509 341667 164575 341670
rect 224953 341667 225019 341670
rect 237005 341730 237071 341733
rect 240041 341730 240107 341733
rect 237005 341728 240107 341730
rect 237005 341672 237010 341728
rect 237066 341672 240046 341728
rect 240102 341672 240107 341728
rect 237005 341670 240107 341672
rect 237005 341667 237071 341670
rect 240041 341667 240107 341670
rect 269389 341730 269455 341733
rect 285397 341730 285463 341733
rect 269389 341728 285463 341730
rect 269389 341672 269394 341728
rect 269450 341672 285402 341728
rect 285458 341672 285463 341728
rect 269389 341670 285463 341672
rect 269389 341667 269455 341670
rect 285397 341667 285463 341670
rect 91093 341594 91159 341597
rect 216673 341594 216739 341597
rect 91093 341592 216739 341594
rect 91093 341536 91098 341592
rect 91154 341536 216678 341592
rect 216734 341536 216739 341592
rect 91093 341534 216739 341536
rect 91093 341531 91159 341534
rect 216673 341531 216739 341534
rect 224902 341532 224908 341596
rect 224972 341594 224978 341596
rect 279550 341594 279556 341596
rect 224972 341534 279556 341594
rect 224972 341532 224978 341534
rect 279550 341532 279556 341534
rect 279620 341532 279626 341596
rect 110321 341458 110387 341461
rect 220721 341458 220787 341461
rect 110321 341456 220787 341458
rect 110321 341400 110326 341456
rect 110382 341400 220726 341456
rect 220782 341400 220787 341456
rect 110321 341398 220787 341400
rect 110321 341395 110387 341398
rect 220721 341395 220787 341398
rect 239213 341458 239279 341461
rect 294229 341458 294295 341461
rect 239213 341456 294295 341458
rect 239213 341400 239218 341456
rect 239274 341400 294234 341456
rect 294290 341400 294295 341456
rect 239213 341398 294295 341400
rect 239213 341395 239279 341398
rect 294229 341395 294295 341398
rect 214649 341322 214715 341325
rect 270401 341322 270467 341325
rect 214649 341320 270467 341322
rect 214649 341264 214654 341320
rect 214710 341264 270406 341320
rect 270462 341264 270467 341320
rect 214649 341262 270467 341264
rect 214649 341259 214715 341262
rect 270401 341259 270467 341262
rect 222878 341124 222884 341188
rect 222948 341186 222954 341188
rect 280286 341186 280292 341188
rect 222948 341126 280292 341186
rect 222948 341124 222954 341126
rect 280286 341124 280292 341126
rect 280356 341124 280362 341188
rect 285673 341186 285739 341189
rect 286910 341186 286916 341188
rect 285673 341184 286916 341186
rect 285673 341128 285678 341184
rect 285734 341128 286916 341184
rect 285673 341126 286916 341128
rect 285673 341123 285739 341126
rect 286910 341124 286916 341126
rect 286980 341124 286986 341188
rect 217961 341050 218027 341053
rect 231117 341050 231183 341053
rect 217961 341048 231183 341050
rect 217961 340992 217966 341048
rect 218022 340992 231122 341048
rect 231178 340992 231183 341048
rect 217961 340990 231183 340992
rect 217961 340987 218027 340990
rect 231117 340987 231183 340990
rect 231526 340988 231532 341052
rect 231596 341050 231602 341052
rect 290590 341050 290596 341052
rect 231596 340990 290596 341050
rect 231596 340988 231602 340990
rect 290590 340988 290596 340990
rect 290660 340988 290666 341052
rect 211654 340852 211660 340916
rect 211724 340914 211730 340916
rect 296478 340914 296484 340916
rect 211724 340854 296484 340914
rect 211724 340852 211730 340854
rect 296478 340852 296484 340854
rect 296548 340852 296554 340916
rect 115565 340778 115631 340781
rect 216765 340778 216831 340781
rect 115565 340776 216831 340778
rect 115565 340720 115570 340776
rect 115626 340720 216770 340776
rect 216826 340720 216831 340776
rect 115565 340718 216831 340720
rect 115565 340715 115631 340718
rect 216765 340715 216831 340718
rect 155769 340642 155835 340645
rect 220721 340642 220787 340645
rect 155769 340640 220787 340642
rect 155769 340584 155774 340640
rect 155830 340584 220726 340640
rect 220782 340584 220787 340640
rect 155769 340582 220787 340584
rect 155769 340579 155835 340582
rect 220721 340579 220787 340582
rect 221222 340580 221228 340644
rect 221292 340642 221298 340644
rect 279918 340642 279924 340644
rect 221292 340582 279924 340642
rect 221292 340580 221298 340582
rect 279918 340580 279924 340582
rect 279988 340580 279994 340644
rect 190729 340506 190795 340509
rect 229921 340506 229987 340509
rect 190729 340504 229987 340506
rect 190729 340448 190734 340504
rect 190790 340448 229926 340504
rect 229982 340448 229987 340504
rect 190729 340446 229987 340448
rect 190729 340443 190795 340446
rect 229921 340443 229987 340446
rect 221038 340308 221044 340372
rect 221108 340370 221114 340372
rect 267590 340370 267596 340372
rect 221108 340310 267596 340370
rect 221108 340308 221114 340310
rect 267590 340308 267596 340310
rect 267660 340308 267666 340372
rect 268377 340370 268443 340373
rect 279734 340370 279740 340372
rect 268377 340368 279740 340370
rect 268377 340312 268382 340368
rect 268438 340312 279740 340368
rect 268377 340310 279740 340312
rect 268377 340307 268443 340310
rect 279734 340308 279740 340310
rect 279804 340308 279810 340372
rect 503621 340370 503687 340373
rect 499806 340368 503687 340370
rect 499806 340312 503626 340368
rect 503682 340312 503687 340368
rect 499806 340310 503687 340312
rect 215886 340172 215892 340236
rect 215956 340234 215962 340236
rect 224217 340234 224283 340237
rect 215956 340232 224283 340234
rect 215956 340176 224222 340232
rect 224278 340176 224283 340232
rect 215956 340174 224283 340176
rect 215956 340172 215962 340174
rect 224217 340171 224283 340174
rect 237833 340234 237899 340237
rect 237966 340234 237972 340236
rect 237833 340232 237972 340234
rect 237833 340176 237838 340232
rect 237894 340176 237972 340232
rect 237833 340174 237972 340176
rect 237833 340171 237899 340174
rect 237966 340172 237972 340174
rect 238036 340172 238042 340236
rect 238150 340172 238156 340236
rect 238220 340234 238226 340236
rect 280102 340234 280108 340236
rect 238220 340174 280108 340234
rect 238220 340172 238226 340174
rect 280102 340172 280108 340174
rect 280172 340172 280178 340236
rect 50337 340098 50403 340101
rect 241421 340098 241487 340101
rect 50337 340096 241487 340098
rect 50337 340040 50342 340096
rect 50398 340040 241426 340096
rect 241482 340040 241487 340096
rect 50337 340038 241487 340040
rect 50337 340035 50403 340038
rect 241421 340035 241487 340038
rect 241605 340098 241671 340101
rect 323761 340098 323827 340101
rect 241605 340096 323827 340098
rect 241605 340040 241610 340096
rect 241666 340040 323766 340096
rect 323822 340040 323827 340096
rect 241605 340038 323827 340040
rect 241605 340035 241671 340038
rect 323761 340035 323827 340038
rect 217777 339962 217843 339965
rect 268377 339962 268443 339965
rect 217777 339960 268443 339962
rect 217777 339904 217782 339960
rect 217838 339904 268382 339960
rect 268438 339904 268443 339960
rect 217777 339902 268443 339904
rect 217777 339899 217843 339902
rect 268377 339899 268443 339902
rect 104801 339826 104867 339829
rect 216673 339826 216739 339829
rect 104801 339824 216739 339826
rect 104801 339768 104806 339824
rect 104862 339768 216678 339824
rect 216734 339768 216739 339824
rect 104801 339766 216739 339768
rect 104801 339763 104867 339766
rect 216673 339763 216739 339766
rect 217593 339826 217659 339829
rect 280061 339826 280127 339829
rect 217593 339824 280127 339826
rect 217593 339768 217598 339824
rect 217654 339768 280066 339824
rect 280122 339768 280127 339824
rect 217593 339766 280127 339768
rect 217593 339763 217659 339766
rect 280061 339763 280127 339766
rect 499806 339728 499866 340310
rect 503621 340307 503687 340310
rect 217174 339628 217180 339692
rect 217244 339690 217250 339692
rect 222009 339690 222075 339693
rect 217244 339688 222075 339690
rect 217244 339632 222014 339688
rect 222070 339632 222075 339688
rect 217244 339630 222075 339632
rect 217244 339628 217250 339630
rect 222009 339627 222075 339630
rect 224217 339690 224283 339693
rect 296846 339690 296852 339692
rect 224217 339688 296852 339690
rect 224217 339632 224222 339688
rect 224278 339632 296852 339688
rect 224217 339630 296852 339632
rect 224217 339627 224283 339630
rect 296846 339628 296852 339630
rect 296916 339628 296922 339692
rect 98637 339554 98703 339557
rect 216857 339554 216923 339557
rect 98637 339552 216923 339554
rect 98637 339496 98642 339552
rect 98698 339496 216862 339552
rect 216918 339496 216923 339552
rect 98637 339494 216923 339496
rect 98637 339491 98703 339494
rect 216857 339491 216923 339494
rect 219934 339492 219940 339556
rect 220004 339554 220010 339556
rect 221917 339554 221983 339557
rect 220004 339552 221983 339554
rect 220004 339496 221922 339552
rect 221978 339496 221983 339552
rect 220004 339494 221983 339496
rect 220004 339492 220010 339494
rect 221917 339491 221983 339494
rect 230238 339492 230244 339556
rect 230308 339554 230314 339556
rect 238150 339554 238156 339556
rect 230308 339494 238156 339554
rect 230308 339492 230314 339494
rect 238150 339492 238156 339494
rect 238220 339492 238226 339556
rect 250989 339554 251055 339557
rect 255998 339554 256004 339556
rect 250989 339552 251098 339554
rect 250989 339496 250994 339552
rect 251050 339496 251098 339552
rect 250989 339491 251098 339496
rect 95877 339418 95943 339421
rect 97257 339418 97323 339421
rect 95877 339416 97323 339418
rect 95877 339360 95882 339416
rect 95938 339360 97262 339416
rect 97318 339360 97323 339416
rect 95877 339358 97323 339360
rect 95877 339355 95943 339358
rect 97257 339355 97323 339358
rect 239765 339418 239831 339421
rect 250897 339418 250963 339421
rect 239765 339416 250963 339418
rect 239765 339360 239770 339416
rect 239826 339360 250902 339416
rect 250958 339360 250963 339416
rect 239765 339358 250963 339360
rect 251038 339418 251098 339491
rect 253660 339494 256004 339554
rect 253660 339418 253720 339494
rect 255998 339492 256004 339494
rect 256068 339492 256074 339556
rect 274582 339554 274588 339556
rect 267598 339494 274588 339554
rect 267598 339418 267658 339494
rect 274582 339492 274588 339494
rect 274652 339492 274658 339556
rect 275737 339554 275803 339557
rect 331857 339554 331923 339557
rect 275737 339552 331923 339554
rect 275737 339496 275742 339552
rect 275798 339496 331862 339552
rect 331918 339496 331923 339552
rect 275737 339494 331923 339496
rect 275737 339491 275803 339494
rect 331857 339491 331923 339494
rect 274633 339418 274699 339421
rect 251038 339358 253720 339418
rect 253890 339358 267658 339418
rect 273210 339416 274699 339418
rect 273210 339360 274638 339416
rect 274694 339360 274699 339416
rect 273210 339358 274699 339360
rect 239765 339355 239831 339358
rect 250897 339355 250963 339358
rect 215109 339146 215175 339149
rect 239213 339146 239279 339149
rect 215109 339144 239279 339146
rect 215109 339088 215114 339144
rect 215170 339088 239218 339144
rect 239274 339088 239279 339144
rect 215109 339086 239279 339088
rect 215109 339083 215175 339086
rect 239213 339083 239279 339086
rect 218830 338948 218836 339012
rect 218900 339010 218906 339012
rect 253890 339010 253950 339358
rect 273210 339282 273270 339358
rect 274633 339355 274699 339358
rect 278405 339418 278471 339421
rect 278405 339416 278514 339418
rect 278405 339360 278410 339416
rect 278466 339360 278514 339416
rect 278405 339355 278514 339360
rect 278998 339356 279004 339420
rect 279068 339418 279074 339420
rect 279969 339418 280035 339421
rect 279068 339416 280035 339418
rect 279068 339360 279974 339416
rect 280030 339360 280035 339416
rect 279068 339358 280035 339360
rect 279068 339356 279074 339358
rect 279969 339355 280035 339358
rect 280153 339418 280219 339421
rect 283833 339418 283899 339421
rect 280153 339416 283899 339418
rect 280153 339360 280158 339416
rect 280214 339360 283838 339416
rect 283894 339360 283899 339416
rect 280153 339358 283899 339360
rect 280153 339355 280219 339358
rect 283833 339355 283899 339358
rect 263550 339222 273270 339282
rect 278454 339282 278514 339355
rect 278454 339222 287070 339282
rect 218900 338950 253950 339010
rect 218900 338948 218906 338950
rect 255998 338948 256004 339012
rect 256068 339010 256074 339012
rect 263550 339010 263610 339222
rect 280061 339146 280127 339149
rect 256068 338950 263610 339010
rect 273210 339144 280127 339146
rect 273210 339088 280066 339144
rect 280122 339088 280127 339144
rect 273210 339086 280127 339088
rect 287010 339146 287070 339222
rect 297541 339146 297607 339149
rect 287010 339144 297607 339146
rect 287010 339088 297546 339144
rect 297602 339088 297607 339144
rect 287010 339086 297607 339088
rect 256068 338948 256074 338950
rect 231117 338874 231183 338877
rect 273210 338874 273270 339086
rect 280061 339083 280127 339086
rect 297541 339083 297607 339086
rect 274582 338948 274588 339012
rect 274652 339010 274658 339012
rect 303838 339010 303844 339012
rect 274652 338950 303844 339010
rect 274652 338948 274658 338950
rect 303838 338948 303844 338950
rect 303908 338948 303914 339012
rect 231117 338872 251190 338874
rect 231117 338816 231122 338872
rect 231178 338816 251190 338872
rect 231117 338814 251190 338816
rect 231117 338811 231183 338814
rect 4102 338676 4108 338740
rect 4172 338738 4178 338740
rect 230974 338738 230980 338740
rect 4172 338678 230980 338738
rect 4172 338676 4178 338678
rect 230974 338676 230980 338678
rect 231044 338676 231050 338740
rect 239765 338738 239831 338741
rect 238710 338736 239831 338738
rect 238710 338680 239770 338736
rect 239826 338680 239831 338736
rect 238710 338678 239831 338680
rect 209313 338602 209379 338605
rect 238710 338602 238770 338678
rect 239765 338675 239831 338678
rect 209313 338600 238770 338602
rect 209313 338544 209318 338600
rect 209374 338544 238770 338600
rect 209313 338542 238770 338544
rect 251130 338602 251190 338814
rect 260790 338814 273270 338874
rect 260790 338602 260850 338814
rect 279918 338812 279924 338876
rect 279988 338874 279994 338876
rect 281901 338874 281967 338877
rect 279988 338872 281967 338874
rect 279988 338816 281906 338872
rect 281962 338816 281967 338872
rect 279988 338814 281967 338816
rect 279988 338812 279994 338814
rect 281901 338811 281967 338814
rect 283833 338874 283899 338877
rect 336641 338874 336707 338877
rect 283833 338872 336707 338874
rect 283833 338816 283838 338872
rect 283894 338816 336646 338872
rect 336702 338816 336707 338872
rect 283833 338814 336707 338816
rect 283833 338811 283899 338814
rect 336641 338811 336707 338814
rect 281257 338738 281323 338741
rect 358629 338738 358695 338741
rect 281257 338736 358695 338738
rect 281257 338680 281262 338736
rect 281318 338680 358634 338736
rect 358690 338680 358695 338736
rect 281257 338678 358695 338680
rect 281257 338675 281323 338678
rect 358629 338675 358695 338678
rect 251130 338542 260850 338602
rect 209313 338539 209379 338542
rect 267590 338540 267596 338604
rect 267660 338602 267666 338604
rect 291510 338602 291516 338604
rect 267660 338542 291516 338602
rect 267660 338540 267666 338542
rect 291510 338540 291516 338542
rect 291580 338540 291586 338604
rect 220486 338404 220492 338468
rect 220556 338466 220562 338468
rect 280061 338466 280127 338469
rect 220556 338464 280127 338466
rect 220556 338408 280066 338464
rect 280122 338408 280127 338464
rect 220556 338406 280127 338408
rect 220556 338404 220562 338406
rect 280061 338403 280127 338406
rect 281901 338466 281967 338469
rect 294638 338466 294644 338468
rect 281901 338464 294644 338466
rect 281901 338408 281906 338464
rect 281962 338408 294644 338464
rect 281901 338406 294644 338408
rect 281901 338403 281967 338406
rect 294638 338404 294644 338406
rect 294708 338404 294714 338468
rect 583520 338452 584960 338692
rect 216070 338268 216076 338332
rect 216140 338330 216146 338332
rect 280061 338330 280127 338333
rect 216140 338328 280127 338330
rect 216140 338272 280066 338328
rect 280122 338272 280127 338328
rect 216140 338270 280127 338272
rect 216140 338268 216146 338270
rect 280061 338267 280127 338270
rect 224166 338132 224172 338196
rect 224236 338194 224242 338196
rect 301814 338194 301820 338196
rect 224236 338134 301820 338194
rect 224236 338132 224242 338134
rect 301814 338132 301820 338134
rect 301884 338132 301890 338196
rect 279550 337996 279556 338060
rect 279620 338058 279626 338060
rect 280061 338058 280127 338061
rect 279620 338056 280127 338058
rect 279620 338000 280066 338056
rect 280122 338000 280127 338056
rect 279620 337998 280127 338000
rect 279620 337996 279626 337998
rect 280061 337995 280127 337998
rect 289997 338058 290063 338061
rect 290774 338058 290780 338060
rect 289997 338056 290780 338058
rect 289997 338000 290002 338056
rect 290058 338000 290780 338056
rect 289997 337998 290780 338000
rect 289997 337995 290063 337998
rect 290774 337996 290780 337998
rect 290844 337996 290850 338060
rect 279734 337860 279740 337924
rect 279804 337922 279810 337924
rect 280153 337922 280219 337925
rect 279804 337920 280219 337922
rect 279804 337864 280158 337920
rect 280214 337864 280219 337920
rect 279804 337862 280219 337864
rect 279804 337860 279810 337862
rect 280153 337859 280219 337862
rect 288617 337922 288683 337925
rect 295425 337922 295491 337925
rect 288617 337920 295491 337922
rect 288617 337864 288622 337920
rect 288678 337864 295430 337920
rect 295486 337864 295491 337920
rect 288617 337862 295491 337864
rect 288617 337859 288683 337862
rect 295425 337859 295491 337862
rect 220118 337724 220124 337788
rect 220188 337786 220194 337788
rect 290958 337786 290964 337788
rect 220188 337726 290964 337786
rect 220188 337724 220194 337726
rect 290958 337724 290964 337726
rect 291028 337724 291034 337788
rect 286869 337514 286935 337517
rect 304165 337514 304231 337517
rect 286869 337512 304231 337514
rect 286869 337456 286874 337512
rect 286930 337456 304170 337512
rect 304226 337456 304231 337512
rect 286869 337454 304231 337456
rect 286869 337451 286935 337454
rect 304165 337451 304231 337454
rect 285121 337378 285187 337381
rect 310421 337378 310487 337381
rect 285121 337376 310487 337378
rect 285121 337320 285126 337376
rect 285182 337320 310426 337376
rect 310482 337320 310487 337376
rect 285121 337318 310487 337320
rect 285121 337315 285187 337318
rect 310421 337315 310487 337318
rect 280061 336698 280127 336701
rect 285990 336698 285996 336700
rect 280061 336696 285996 336698
rect 280061 336640 280066 336696
rect 280122 336640 285996 336696
rect 280061 336638 285996 336640
rect 280061 336635 280127 336638
rect 285990 336636 285996 336638
rect 286060 336636 286066 336700
rect 280153 336290 280219 336293
rect 295793 336290 295859 336293
rect 280153 336288 295859 336290
rect 280153 336232 280158 336288
rect 280214 336232 295798 336288
rect 295854 336232 295859 336288
rect 280153 336230 295859 336232
rect 280153 336227 280219 336230
rect 295793 336227 295859 336230
rect 281349 336154 281415 336157
rect 299657 336154 299723 336157
rect 281349 336152 299723 336154
rect 281349 336096 281354 336152
rect 281410 336096 299662 336152
rect 299718 336096 299723 336152
rect 281349 336094 299723 336096
rect 281349 336091 281415 336094
rect 299657 336091 299723 336094
rect 281165 336018 281231 336021
rect 358537 336018 358603 336021
rect 281165 336016 358603 336018
rect 281165 335960 281170 336016
rect 281226 335960 358542 336016
rect 358598 335960 358603 336016
rect 281165 335958 358603 335960
rect 281165 335955 281231 335958
rect 358537 335955 358603 335958
rect 290365 334114 290431 334117
rect 290365 334112 360210 334114
rect 290365 334056 290370 334112
rect 290426 334056 360210 334112
rect 290365 334054 360210 334056
rect 290365 334051 290431 334054
rect 360150 334016 360210 334054
rect 503621 333842 503687 333845
rect 499806 333840 503687 333842
rect 499806 333784 503626 333840
rect 503682 333784 503687 333840
rect 499806 333782 503687 333784
rect 499806 333744 499866 333782
rect 503621 333779 503687 333782
rect 295425 333026 295491 333029
rect 295425 333024 360210 333026
rect 295425 332968 295430 333024
rect 295486 332968 360210 333024
rect 295425 332966 360210 332968
rect 295425 332963 295491 332966
rect 360150 332928 360210 332966
rect -960 332196 480 332436
rect 304165 331938 304231 331941
rect 304165 331936 360210 331938
rect 304165 331880 304170 331936
rect 304226 331880 360210 331936
rect 304165 331878 360210 331880
rect 304165 331875 304231 331878
rect 360150 331840 360210 331878
rect 310421 330850 310487 330853
rect 310421 330848 360210 330850
rect 310421 330792 310426 330848
rect 310482 330792 360210 330848
rect 310421 330790 360210 330792
rect 310421 330787 310487 330790
rect 360150 330752 360210 330790
rect 286685 329762 286751 329765
rect 286685 329760 360210 329762
rect 286685 329704 286690 329760
rect 286746 329704 360210 329760
rect 286685 329702 360210 329704
rect 286685 329699 286751 329702
rect 360150 329664 360210 329702
rect 292113 328674 292179 328677
rect 292113 328672 360210 328674
rect 292113 328616 292118 328672
rect 292174 328616 360210 328672
rect 292113 328614 360210 328616
rect 292113 328611 292179 328614
rect 360150 328576 360210 328614
rect 503621 328130 503687 328133
rect 499806 328128 503687 328130
rect 499806 328072 503626 328128
rect 503682 328072 503687 328128
rect 499806 328070 503687 328072
rect 499806 327760 499866 328070
rect 503621 328067 503687 328070
rect 336641 327586 336707 327589
rect 336641 327584 360210 327586
rect 336641 327528 336646 327584
rect 336702 327528 360210 327584
rect 336641 327526 360210 327528
rect 336641 327523 336707 327526
rect 360150 327488 360210 327526
rect 237741 327450 237807 327453
rect 237741 327448 239690 327450
rect 237741 327392 237746 327448
rect 237802 327392 239690 327448
rect 237741 327390 239690 327392
rect 237741 327387 237807 327390
rect 239630 327382 239690 327390
rect 239630 327322 240212 327382
rect 228725 326498 228791 326501
rect 237741 326498 237807 326501
rect 228725 326496 237807 326498
rect 228725 326440 228730 326496
rect 228786 326440 237746 326496
rect 237802 326440 237807 326496
rect 228725 326438 237807 326440
rect 228725 326435 228791 326438
rect 237741 326435 237807 326438
rect 297541 326498 297607 326501
rect 297541 326496 360210 326498
rect 297541 326440 297546 326496
rect 297602 326440 360210 326496
rect 297541 326438 360210 326440
rect 297541 326435 297607 326438
rect 360150 326400 360210 326438
rect 3550 326300 3556 326364
rect 3620 326362 3626 326364
rect 224309 326362 224375 326365
rect 3620 326360 224375 326362
rect 3620 326304 224314 326360
rect 224370 326304 224375 326360
rect 3620 326302 224375 326304
rect 3620 326300 3626 326302
rect 224309 326299 224375 326302
rect 231209 326362 231275 326365
rect 231209 326360 239690 326362
rect 231209 326304 231214 326360
rect 231270 326304 239690 326360
rect 231209 326302 239690 326304
rect 231209 326299 231275 326302
rect 239630 326294 239690 326302
rect 239630 326234 240212 326294
rect 358445 325546 358511 325549
rect 358445 325544 360210 325546
rect 358445 325488 358450 325544
rect 358506 325488 360210 325544
rect 358445 325486 360210 325488
rect 358445 325483 358511 325486
rect 360150 325312 360210 325486
rect 238017 325274 238083 325277
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 238017 325272 239690 325274
rect 238017 325216 238022 325272
rect 238078 325216 239690 325272
rect 238017 325214 239690 325216
rect 238017 325211 238083 325214
rect 239630 325206 239690 325214
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 239630 325146 240212 325206
rect 583520 325124 584960 325214
rect 295057 324322 295123 324325
rect 295057 324320 360210 324322
rect 295057 324264 295062 324320
rect 295118 324264 360210 324320
rect 295057 324262 360210 324264
rect 295057 324259 295123 324262
rect 360150 324224 360210 324262
rect 238109 324186 238175 324189
rect 238109 324184 239690 324186
rect 238109 324128 238114 324184
rect 238170 324128 239690 324184
rect 238109 324126 239690 324128
rect 238109 324123 238175 324126
rect 239630 324118 239690 324126
rect 239630 324058 240212 324118
rect 358629 323778 358695 323781
rect 358629 323776 360210 323778
rect 358629 323720 358634 323776
rect 358690 323720 360210 323776
rect 358629 323718 360210 323720
rect 358629 323715 358695 323718
rect 228817 323642 228883 323645
rect 237833 323642 237899 323645
rect 228817 323640 237899 323642
rect 228817 323584 228822 323640
rect 228878 323584 237838 323640
rect 237894 323584 237899 323640
rect 228817 323582 237899 323584
rect 228817 323579 228883 323582
rect 237833 323579 237899 323582
rect 360150 323136 360210 323718
rect 237097 323098 237163 323101
rect 237097 323096 239690 323098
rect 237097 323040 237102 323096
rect 237158 323040 239690 323096
rect 237097 323038 239690 323040
rect 237097 323035 237163 323038
rect 239630 323030 239690 323038
rect 239630 322970 240212 323030
rect 503621 322418 503687 322421
rect 499806 322416 503687 322418
rect 499806 322360 503626 322416
rect 503682 322360 503687 322416
rect 499806 322358 503687 322360
rect 285305 322146 285371 322149
rect 285305 322144 360210 322146
rect 285305 322088 285310 322144
rect 285366 322088 360210 322144
rect 285305 322086 360210 322088
rect 285305 322083 285371 322086
rect 360150 322048 360210 322086
rect 239397 322010 239463 322013
rect 239397 322008 239690 322010
rect 239397 321952 239402 322008
rect 239458 321952 239690 322008
rect 239397 321950 239690 321952
rect 239397 321947 239463 321950
rect 239630 321942 239690 321950
rect 239630 321882 240212 321942
rect 499806 321776 499866 322358
rect 503621 322355 503687 322358
rect 86217 321602 86283 321605
rect 86217 321600 113190 321602
rect 86217 321544 86222 321600
rect 86278 321544 113190 321600
rect 86217 321542 113190 321544
rect 86217 321539 86283 321542
rect 113130 321466 113190 321542
rect 113817 321466 113883 321469
rect 237925 321466 237991 321469
rect 113130 321464 237991 321466
rect 113130 321408 113822 321464
rect 113878 321408 237930 321464
rect 237986 321408 237991 321464
rect 113130 321406 237991 321408
rect 113817 321403 113883 321406
rect 237925 321403 237991 321406
rect 285397 321058 285463 321061
rect 285397 321056 360210 321058
rect 285397 321000 285402 321056
rect 285458 321000 360210 321056
rect 285397 320998 360210 321000
rect 285397 320995 285463 320998
rect 360150 320960 360210 320998
rect 230013 320922 230079 320925
rect 230013 320920 239690 320922
rect 230013 320864 230018 320920
rect 230074 320864 239690 320920
rect 230013 320862 239690 320864
rect 230013 320859 230079 320862
rect 239630 320854 239690 320862
rect 239630 320794 240212 320854
rect 300577 319970 300643 319973
rect 300577 319968 360210 319970
rect 300577 319912 300582 319968
rect 300638 319912 360210 319968
rect 300577 319910 360210 319912
rect 300577 319907 300643 319910
rect 360150 319872 360210 319910
rect 236729 319834 236795 319837
rect 236729 319832 239690 319834
rect 236729 319776 236734 319832
rect 236790 319776 239690 319832
rect 236729 319774 239690 319776
rect 236729 319771 236795 319774
rect 239630 319766 239690 319774
rect 239630 319706 240212 319766
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 288157 318882 288223 318885
rect 288157 318880 360210 318882
rect 288157 318824 288162 318880
rect 288218 318824 360210 318880
rect 288157 318822 360210 318824
rect 288157 318819 288223 318822
rect 360150 318784 360210 318822
rect 227529 318746 227595 318749
rect 227529 318744 239690 318746
rect 227529 318688 227534 318744
rect 227590 318688 239690 318744
rect 227529 318686 239690 318688
rect 227529 318683 227595 318686
rect 239630 318678 239690 318686
rect 239630 318618 240212 318678
rect 280889 317794 280955 317797
rect 280889 317792 360210 317794
rect 280889 317736 280894 317792
rect 280950 317736 360210 317792
rect 280889 317734 360210 317736
rect 280889 317731 280955 317734
rect 360150 317696 360210 317734
rect 238201 317658 238267 317661
rect 238201 317656 239690 317658
rect 238201 317600 238206 317656
rect 238262 317600 239690 317656
rect 238201 317598 239690 317600
rect 238201 317595 238267 317598
rect 239630 317590 239690 317598
rect 239630 317530 240212 317590
rect 232497 317386 232563 317389
rect 238017 317386 238083 317389
rect 232497 317384 238083 317386
rect 232497 317328 232502 317384
rect 232558 317328 238022 317384
rect 238078 317328 238083 317384
rect 232497 317326 238083 317328
rect 232497 317323 232563 317326
rect 238017 317323 238083 317326
rect 358537 317250 358603 317253
rect 358537 317248 360210 317250
rect 358537 317192 358542 317248
rect 358598 317192 360210 317248
rect 358537 317190 360210 317192
rect 358537 317187 358603 317190
rect 360150 316608 360210 317190
rect 239489 316570 239555 316573
rect 239489 316568 239690 316570
rect 239489 316512 239494 316568
rect 239550 316512 239690 316568
rect 239489 316510 239690 316512
rect 239489 316507 239555 316510
rect 239630 316502 239690 316510
rect 239630 316442 240212 316502
rect 522062 315890 522068 315892
rect 499806 315830 522068 315890
rect 499806 315792 499866 315830
rect 522062 315828 522068 315830
rect 522132 315828 522138 315892
rect 292297 315618 292363 315621
rect 292297 315616 360210 315618
rect 292297 315560 292302 315616
rect 292358 315560 360210 315616
rect 292297 315558 360210 315560
rect 292297 315555 292363 315558
rect 360150 315520 360210 315558
rect 238569 315482 238635 315485
rect 238569 315480 239690 315482
rect 238569 315424 238574 315480
rect 238630 315424 239690 315480
rect 238569 315422 239690 315424
rect 238569 315419 238635 315422
rect 239630 315414 239690 315422
rect 239630 315354 240212 315414
rect 351177 314530 351243 314533
rect 351177 314528 360210 314530
rect 351177 314472 351182 314528
rect 351238 314472 360210 314528
rect 351177 314470 360210 314472
rect 351177 314467 351243 314470
rect 360150 314432 360210 314470
rect 238293 314394 238359 314397
rect 238293 314392 239690 314394
rect 238293 314336 238298 314392
rect 238354 314336 239690 314392
rect 238293 314334 239690 314336
rect 238293 314331 238359 314334
rect 239630 314326 239690 314334
rect 239630 314266 240212 314326
rect 238569 313986 238635 313989
rect 239305 313986 239371 313989
rect 238569 313984 239371 313986
rect 238569 313928 238574 313984
rect 238630 313928 239310 313984
rect 239366 313928 239371 313984
rect 238569 313926 239371 313928
rect 238569 313923 238635 313926
rect 239305 313923 239371 313926
rect 288249 313442 288315 313445
rect 288249 313440 360210 313442
rect 288249 313384 288254 313440
rect 288310 313384 360210 313440
rect 288249 313382 360210 313384
rect 288249 313379 288315 313382
rect 360150 313344 360210 313382
rect 239630 313178 240212 313238
rect 230105 313170 230171 313173
rect 239630 313170 239690 313178
rect 230105 313168 239690 313170
rect 230105 313112 230110 313168
rect 230166 313112 239690 313168
rect 230105 313110 239690 313112
rect 230105 313107 230171 313110
rect 8109 312490 8175 312493
rect 178677 312490 178743 312493
rect 8109 312488 178743 312490
rect 8109 312432 8114 312488
rect 8170 312432 178682 312488
rect 178738 312432 178743 312488
rect 8109 312430 178743 312432
rect 8109 312427 8175 312430
rect 178677 312427 178743 312430
rect 299197 312354 299263 312357
rect 299197 312352 360210 312354
rect 299197 312296 299202 312352
rect 299258 312296 360210 312352
rect 299197 312294 360210 312296
rect 299197 312291 299263 312294
rect 360150 312256 360210 312294
rect 231301 312218 231367 312221
rect 231301 312216 239690 312218
rect 231301 312160 231306 312216
rect 231362 312160 239690 312216
rect 231301 312158 239690 312160
rect 231301 312155 231367 312158
rect 239630 312150 239690 312158
rect 239630 312090 240212 312150
rect 580390 312020 580396 312084
rect 580460 312082 580466 312084
rect 583520 312082 584960 312172
rect 580460 312022 584960 312082
rect 580460 312020 580466 312022
rect 583520 311932 584960 312022
rect 286777 311266 286843 311269
rect 286777 311264 360210 311266
rect 286777 311208 286782 311264
rect 286838 311208 360210 311264
rect 286777 311206 360210 311208
rect 286777 311203 286843 311206
rect 360150 311168 360210 311206
rect 228909 311130 228975 311133
rect 228909 311128 239690 311130
rect 228909 311072 228914 311128
rect 228970 311072 239690 311128
rect 228909 311070 239690 311072
rect 228909 311067 228975 311070
rect 239630 311062 239690 311070
rect 239630 311002 240212 311062
rect 350441 310178 350507 310181
rect 350441 310176 360210 310178
rect 350441 310120 350446 310176
rect 350502 310120 360210 310176
rect 350441 310118 360210 310120
rect 350441 310115 350507 310118
rect 360150 310080 360210 310118
rect 234102 309844 234108 309908
rect 234172 309906 234178 309908
rect 521878 309906 521884 309908
rect 234172 309846 240212 309906
rect 499806 309846 521884 309906
rect 234172 309844 234178 309846
rect 499806 309808 499866 309846
rect 521878 309844 521884 309846
rect 521948 309844 521954 309908
rect 280470 309362 280476 309364
rect 279956 309302 280476 309362
rect 280470 309300 280476 309302
rect 280540 309300 280546 309364
rect 345657 309090 345723 309093
rect 345657 309088 360210 309090
rect 345657 309032 345662 309088
rect 345718 309032 360210 309088
rect 345657 309030 360210 309032
rect 345657 309027 345723 309030
rect 360150 308992 360210 309030
rect 238477 308818 238543 308821
rect 280705 308818 280771 308821
rect 238477 308816 240212 308818
rect 238477 308760 238482 308816
rect 238538 308760 240212 308816
rect 238477 308758 240212 308760
rect 279956 308816 280771 308818
rect 279956 308760 280710 308816
rect 280766 308760 280771 308816
rect 279956 308758 280771 308760
rect 238477 308755 238543 308758
rect 280705 308755 280771 308758
rect 282913 308274 282979 308277
rect 279956 308272 282979 308274
rect 279956 308216 282918 308272
rect 282974 308216 282979 308272
rect 279956 308214 282979 308216
rect 282913 308211 282979 308214
rect 327809 308002 327875 308005
rect 327809 308000 360210 308002
rect 327809 307944 327814 308000
rect 327870 307944 360210 308000
rect 327809 307942 360210 307944
rect 327809 307939 327875 307942
rect 360150 307904 360210 307942
rect 230197 307730 230263 307733
rect 281809 307730 281875 307733
rect 230197 307728 240212 307730
rect 230197 307672 230202 307728
rect 230258 307672 240212 307728
rect 230197 307670 240212 307672
rect 279956 307728 281875 307730
rect 279956 307672 281814 307728
rect 281870 307672 281875 307728
rect 279956 307670 281875 307672
rect 230197 307667 230263 307670
rect 281809 307667 281875 307670
rect 280613 307186 280679 307189
rect 279956 307184 280679 307186
rect 279956 307128 280618 307184
rect 280674 307128 280679 307184
rect 279956 307126 280679 307128
rect 280613 307123 280679 307126
rect 280981 306914 281047 306917
rect 280981 306912 360210 306914
rect 280981 306856 280986 306912
rect 281042 306856 360210 306912
rect 280981 306854 360210 306856
rect 280981 306851 281047 306854
rect 360150 306816 360210 306854
rect 231393 306642 231459 306645
rect 283189 306642 283255 306645
rect 231393 306640 240212 306642
rect 231393 306584 231398 306640
rect 231454 306584 240212 306640
rect 231393 306582 240212 306584
rect 279956 306640 283255 306642
rect 279956 306584 283194 306640
rect 283250 306584 283255 306640
rect 279956 306582 283255 306584
rect 231393 306579 231459 306582
rect 283189 306579 283255 306582
rect 334801 306506 334867 306509
rect 337377 306506 337443 306509
rect 334801 306504 337443 306506
rect 334801 306448 334806 306504
rect 334862 306448 337382 306504
rect 337438 306448 337443 306504
rect 334801 306446 337443 306448
rect 334801 306443 334867 306446
rect 337377 306443 337443 306446
rect -960 306234 480 306324
rect 214782 306234 214788 306236
rect -960 306174 214788 306234
rect -960 306084 480 306174
rect 214782 306172 214788 306174
rect 214852 306172 214858 306236
rect 283557 306098 283623 306101
rect 279956 306096 283623 306098
rect 279956 306040 283562 306096
rect 283618 306040 283623 306096
rect 279956 306038 283623 306040
rect 283557 306035 283623 306038
rect 334709 305826 334775 305829
rect 334709 305824 360210 305826
rect 334709 305768 334714 305824
rect 334770 305768 360210 305824
rect 334709 305766 360210 305768
rect 334709 305763 334775 305766
rect 360150 305728 360210 305766
rect 236821 305554 236887 305557
rect 280429 305554 280495 305557
rect 236821 305552 240212 305554
rect 236821 305496 236826 305552
rect 236882 305496 240212 305552
rect 236821 305494 240212 305496
rect 279956 305552 280495 305554
rect 279956 305496 280434 305552
rect 280490 305496 280495 305552
rect 279956 305494 280495 305496
rect 236821 305491 236887 305494
rect 280429 305491 280495 305494
rect 283097 305010 283163 305013
rect 279956 305008 283163 305010
rect 279956 304952 283102 305008
rect 283158 304952 283163 305008
rect 279956 304950 283163 304952
rect 283097 304947 283163 304950
rect 292205 304738 292271 304741
rect 292205 304736 360210 304738
rect 292205 304680 292210 304736
rect 292266 304680 360210 304736
rect 292205 304678 360210 304680
rect 292205 304675 292271 304678
rect 360150 304640 360210 304678
rect 239581 304466 239647 304469
rect 280337 304466 280403 304469
rect 503621 304466 503687 304469
rect 239581 304464 240212 304466
rect 239581 304408 239586 304464
rect 239642 304408 240212 304464
rect 239581 304406 240212 304408
rect 279956 304464 280403 304466
rect 279956 304408 280342 304464
rect 280398 304408 280403 304464
rect 279956 304406 280403 304408
rect 239581 304403 239647 304406
rect 280337 304403 280403 304406
rect 499806 304464 503687 304466
rect 499806 304408 503626 304464
rect 503682 304408 503687 304464
rect 499806 304406 503687 304408
rect 280245 303922 280311 303925
rect 279956 303920 280311 303922
rect 279956 303864 280250 303920
rect 280306 303864 280311 303920
rect 279956 303862 280311 303864
rect 280245 303859 280311 303862
rect 499806 303824 499866 304406
rect 503621 304403 503687 304406
rect 323761 303514 323827 303517
rect 360150 303514 360210 303552
rect 323761 303512 360210 303514
rect 323761 303456 323766 303512
rect 323822 303456 360210 303512
rect 323761 303454 360210 303456
rect 323761 303451 323827 303454
rect 236545 303378 236611 303381
rect 284518 303378 284524 303380
rect 236545 303376 240212 303378
rect 236545 303320 236550 303376
rect 236606 303320 240212 303376
rect 236545 303318 240212 303320
rect 279956 303318 284524 303378
rect 236545 303315 236611 303318
rect 284518 303316 284524 303318
rect 284588 303316 284594 303380
rect 49325 303242 49391 303245
rect 62021 303242 62087 303245
rect 49325 303240 62087 303242
rect 49325 303184 49330 303240
rect 49386 303184 62026 303240
rect 62082 303184 62087 303240
rect 49325 303182 62087 303184
rect 49325 303179 49391 303182
rect 62021 303179 62087 303182
rect 49601 303106 49667 303109
rect 66161 303106 66227 303109
rect 49601 303104 66227 303106
rect 49601 303048 49606 303104
rect 49662 303048 66166 303104
rect 66222 303048 66227 303104
rect 49601 303046 66227 303048
rect 49601 303043 49667 303046
rect 66161 303043 66227 303046
rect 48037 302970 48103 302973
rect 68921 302970 68987 302973
rect 48037 302968 68987 302970
rect 48037 302912 48042 302968
rect 48098 302912 68926 302968
rect 68982 302912 68987 302968
rect 48037 302910 68987 302912
rect 48037 302907 48103 302910
rect 68921 302907 68987 302910
rect 75821 302970 75887 302973
rect 86217 302970 86283 302973
rect 75821 302968 86283 302970
rect 75821 302912 75826 302968
rect 75882 302912 86222 302968
rect 86278 302912 86283 302968
rect 75821 302910 86283 302912
rect 75821 302907 75887 302910
rect 86217 302907 86283 302910
rect 50521 302834 50587 302837
rect 71589 302834 71655 302837
rect 231117 302834 231183 302837
rect 280521 302834 280587 302837
rect 50521 302832 71655 302834
rect 50521 302776 50526 302832
rect 50582 302776 71594 302832
rect 71650 302776 71655 302832
rect 50521 302774 71655 302776
rect 50521 302771 50587 302774
rect 71589 302771 71655 302774
rect 74490 302832 231183 302834
rect 74490 302776 231122 302832
rect 231178 302776 231183 302832
rect 74490 302774 231183 302776
rect 279956 302832 280587 302834
rect 279956 302776 280526 302832
rect 280582 302776 280587 302832
rect 279956 302774 280587 302776
rect 48129 302426 48195 302429
rect 63493 302426 63559 302429
rect 48129 302424 63559 302426
rect 48129 302368 48134 302424
rect 48190 302368 63498 302424
rect 63554 302368 63559 302424
rect 48129 302366 63559 302368
rect 48129 302363 48195 302366
rect 63493 302363 63559 302366
rect 50429 302290 50495 302293
rect 74257 302290 74323 302293
rect 74490 302290 74550 302774
rect 231117 302771 231183 302774
rect 280521 302771 280587 302774
rect 312537 302834 312603 302837
rect 339125 302834 339191 302837
rect 312537 302832 339191 302834
rect 312537 302776 312542 302832
rect 312598 302776 339130 302832
rect 339186 302776 339191 302832
rect 312537 302774 339191 302776
rect 312537 302771 312603 302774
rect 339125 302771 339191 302774
rect 321093 302562 321159 302565
rect 321093 302560 360210 302562
rect 321093 302504 321098 302560
rect 321154 302504 360210 302560
rect 321093 302502 360210 302504
rect 321093 302499 321159 302502
rect 360150 302464 360210 302502
rect 50429 302288 74550 302290
rect 50429 302232 50434 302288
rect 50490 302232 74262 302288
rect 74318 302232 74550 302288
rect 50429 302230 74550 302232
rect 81065 302290 81131 302293
rect 96521 302290 96587 302293
rect 125685 302290 125751 302293
rect 81065 302288 93870 302290
rect 81065 302232 81070 302288
rect 81126 302232 93870 302288
rect 81065 302230 93870 302232
rect 50429 302227 50495 302230
rect 74257 302227 74323 302230
rect 81065 302227 81131 302230
rect 93810 301610 93870 302230
rect 96521 302288 125751 302290
rect 96521 302232 96526 302288
rect 96582 302232 125690 302288
rect 125746 302232 125751 302288
rect 96521 302230 125751 302232
rect 96521 302227 96587 302230
rect 125685 302227 125751 302230
rect 236637 302290 236703 302293
rect 283005 302290 283071 302293
rect 236637 302288 240212 302290
rect 236637 302232 236642 302288
rect 236698 302232 240212 302288
rect 236637 302230 240212 302232
rect 279956 302288 283071 302290
rect 279956 302232 283010 302288
rect 283066 302232 283071 302288
rect 279956 302230 283071 302232
rect 236637 302227 236703 302230
rect 283005 302227 283071 302230
rect 294454 301746 294460 301748
rect 279956 301686 294460 301746
rect 294454 301684 294460 301686
rect 294524 301684 294530 301748
rect 126881 301610 126947 301613
rect 93810 301608 126947 301610
rect 93810 301552 126886 301608
rect 126942 301552 126947 301608
rect 93810 301550 126947 301552
rect 126881 301547 126947 301550
rect 55070 301412 55076 301476
rect 55140 301474 55146 301476
rect 229829 301474 229895 301477
rect 55140 301472 229895 301474
rect 55140 301416 229834 301472
rect 229890 301416 229895 301472
rect 55140 301414 229895 301416
rect 55140 301412 55146 301414
rect 229829 301411 229895 301414
rect 280797 301474 280863 301477
rect 280797 301472 360210 301474
rect 280797 301416 280802 301472
rect 280858 301416 360210 301472
rect 280797 301414 360210 301416
rect 280797 301411 280863 301414
rect 360150 301376 360210 301414
rect 49509 301202 49575 301205
rect 61285 301202 61351 301205
rect 49509 301200 61351 301202
rect 49509 301144 49514 301200
rect 49570 301144 61290 301200
rect 61346 301144 61351 301200
rect 49509 301142 61351 301144
rect 49509 301139 49575 301142
rect 61285 301139 61351 301142
rect 231485 301202 231551 301205
rect 291377 301202 291443 301205
rect 231485 301200 240212 301202
rect 231485 301144 231490 301200
rect 231546 301144 240212 301200
rect 231485 301142 240212 301144
rect 279956 301200 291443 301202
rect 279956 301144 291382 301200
rect 291438 301144 291443 301200
rect 279956 301142 291443 301144
rect 231485 301139 231551 301142
rect 291377 301139 291443 301142
rect 47945 301066 48011 301069
rect 66069 301066 66135 301069
rect 47945 301064 66135 301066
rect 47945 301008 47950 301064
rect 48006 301008 66074 301064
rect 66130 301008 66135 301064
rect 47945 301006 66135 301008
rect 47945 301003 48011 301006
rect 66069 301003 66135 301006
rect 105905 301066 105971 301069
rect 133873 301066 133939 301069
rect 105905 301064 133939 301066
rect 105905 301008 105910 301064
rect 105966 301008 133878 301064
rect 133934 301008 133939 301064
rect 105905 301006 133939 301008
rect 105905 301003 105971 301006
rect 133873 301003 133939 301006
rect 49417 300930 49483 300933
rect 71221 300930 71287 300933
rect 49417 300928 71287 300930
rect 49417 300872 49422 300928
rect 49478 300872 71226 300928
rect 71282 300872 71287 300928
rect 49417 300870 71287 300872
rect 49417 300867 49483 300870
rect 71221 300867 71287 300870
rect 97717 300930 97783 300933
rect 132585 300930 132651 300933
rect 97717 300928 132651 300930
rect 97717 300872 97722 300928
rect 97778 300872 132590 300928
rect 132646 300872 132651 300928
rect 97717 300870 132651 300872
rect 97717 300867 97783 300870
rect 132585 300867 132651 300870
rect 126329 300794 126395 300797
rect 126881 300794 126947 300797
rect 228541 300794 228607 300797
rect 126329 300792 228607 300794
rect 126329 300736 126334 300792
rect 126390 300736 126886 300792
rect 126942 300736 228546 300792
rect 228602 300736 228607 300792
rect 126329 300734 228607 300736
rect 126329 300731 126395 300734
rect 126881 300731 126947 300734
rect 228541 300731 228607 300734
rect 332041 300794 332107 300797
rect 333513 300794 333579 300797
rect 332041 300792 333579 300794
rect 332041 300736 332046 300792
rect 332102 300736 333518 300792
rect 333574 300736 333579 300792
rect 332041 300734 333579 300736
rect 332041 300731 332107 300734
rect 333513 300731 333579 300734
rect 291142 300658 291148 300660
rect 279956 300598 291148 300658
rect 291142 300596 291148 300598
rect 291212 300596 291218 300660
rect 294965 300386 295031 300389
rect 294965 300384 360210 300386
rect 294965 300328 294970 300384
rect 295026 300328 360210 300384
rect 294965 300326 360210 300328
rect 294965 300323 295031 300326
rect 360150 300288 360210 300326
rect 97257 300114 97323 300117
rect 110321 300114 110387 300117
rect 97257 300112 110387 300114
rect 97257 300056 97262 300112
rect 97318 300056 110326 300112
rect 110382 300056 110387 300112
rect 97257 300054 110387 300056
rect 97257 300051 97323 300054
rect 110321 300051 110387 300054
rect 239673 300114 239739 300117
rect 292614 300114 292620 300116
rect 239673 300112 240212 300114
rect 239673 300056 239678 300112
rect 239734 300056 240212 300112
rect 239673 300054 240212 300056
rect 279956 300054 292620 300114
rect 239673 300051 239739 300054
rect 292614 300052 292620 300054
rect 292684 300052 292690 300116
rect 107239 299706 107305 299709
rect 131205 299706 131271 299709
rect 107239 299704 131271 299706
rect 107239 299648 107244 299704
rect 107300 299648 131210 299704
rect 131266 299648 131271 299704
rect 107239 299646 131271 299648
rect 107239 299643 107305 299646
rect 131205 299643 131271 299646
rect 108895 299570 108961 299573
rect 135253 299570 135319 299573
rect 295425 299570 295491 299573
rect 108895 299568 135319 299570
rect 108895 299512 108900 299568
rect 108956 299512 135258 299568
rect 135314 299512 135319 299568
rect 108895 299510 135319 299512
rect 279956 299568 295491 299570
rect 279956 299512 295430 299568
rect 295486 299512 295491 299568
rect 279956 299510 295491 299512
rect 108895 299507 108961 299510
rect 135253 299507 135319 299510
rect 295425 299507 295491 299510
rect 287830 299372 287836 299436
rect 287900 299434 287906 299436
rect 290181 299434 290247 299437
rect 287900 299432 290247 299434
rect 287900 299376 290186 299432
rect 290242 299376 290247 299432
rect 287900 299374 290247 299376
rect 287900 299372 287906 299374
rect 290181 299371 290247 299374
rect 300853 299434 300919 299437
rect 357249 299434 357315 299437
rect 300853 299432 357315 299434
rect 300853 299376 300858 299432
rect 300914 299376 357254 299432
rect 357310 299376 357315 299432
rect 300853 299374 357315 299376
rect 300853 299371 300919 299374
rect 357249 299371 357315 299374
rect 290733 299298 290799 299301
rect 290733 299296 360210 299298
rect 290733 299240 290738 299296
rect 290794 299240 360210 299296
rect 290733 299238 360210 299240
rect 290733 299235 290799 299238
rect 360150 299200 360210 299238
rect 226149 299026 226215 299029
rect 293953 299026 294019 299029
rect 226149 299024 240212 299026
rect 226149 298968 226154 299024
rect 226210 298968 240212 299024
rect 226149 298966 240212 298968
rect 279956 299024 294019 299026
rect 279956 298968 293958 299024
rect 294014 298968 294019 299024
rect 279956 298966 294019 298968
rect 226149 298963 226215 298966
rect 293953 298963 294019 298966
rect 358261 298754 358327 298757
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 358261 298752 360210 298754
rect 358261 298696 358266 298752
rect 358322 298696 360210 298752
rect 358261 298694 360210 298696
rect 358261 298691 358327 298694
rect 223062 298618 223068 298620
rect 109940 298558 223068 298618
rect 223062 298556 223068 298558
rect 223132 298556 223138 298620
rect 281901 298482 281967 298485
rect 279956 298480 281967 298482
rect 279956 298424 281906 298480
rect 281962 298424 281967 298480
rect 279956 298422 281967 298424
rect 281901 298419 281967 298422
rect 360150 298112 360210 298694
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 216622 298012 216628 298076
rect 216692 298074 216698 298076
rect 217961 298074 218027 298077
rect 216692 298072 218027 298074
rect 216692 298016 217966 298072
rect 218022 298016 218027 298072
rect 216692 298014 218027 298016
rect 216692 298012 216698 298014
rect 217961 298011 218027 298014
rect 238017 297938 238083 297941
rect 287278 297938 287284 297940
rect 238017 297936 240212 297938
rect 238017 297880 238022 297936
rect 238078 297880 240212 297936
rect 238017 297878 240212 297880
rect 279956 297878 287284 297938
rect 238017 297875 238083 297878
rect 287278 297876 287284 297878
rect 287348 297876 287354 297940
rect 503621 297938 503687 297941
rect 499806 297936 503687 297938
rect 499806 297880 503626 297936
rect 503682 297880 503687 297936
rect 499806 297878 503687 297880
rect 499806 297840 499866 297878
rect 503621 297875 503687 297878
rect 287094 297394 287100 297396
rect 279956 297334 287100 297394
rect 287094 297332 287100 297334
rect 287164 297332 287170 297396
rect 296253 297122 296319 297125
rect 296253 297120 360210 297122
rect 296253 297064 296258 297120
rect 296314 297064 360210 297120
rect 296253 297062 360210 297064
rect 296253 297059 296319 297062
rect 360150 297024 360210 297062
rect 217542 296986 217548 296988
rect 110462 296926 217548 296986
rect 110462 296918 110522 296926
rect 217542 296924 217548 296926
rect 217612 296924 217618 296988
rect 109940 296858 110522 296918
rect 237741 296850 237807 296853
rect 285622 296850 285628 296852
rect 237741 296848 240212 296850
rect 237741 296792 237746 296848
rect 237802 296792 240212 296848
rect 237741 296790 240212 296792
rect 279956 296790 285628 296850
rect 237741 296787 237807 296790
rect 285622 296788 285628 296790
rect 285692 296788 285698 296852
rect 287462 296306 287468 296308
rect 279956 296246 287468 296306
rect 287462 296244 287468 296246
rect 287532 296244 287538 296308
rect 305913 296034 305979 296037
rect 305913 296032 360210 296034
rect 305913 295976 305918 296032
rect 305974 295976 360210 296032
rect 305913 295974 360210 295976
rect 305913 295971 305979 295974
rect 360150 295936 360210 295974
rect 226241 295762 226307 295765
rect 285765 295762 285831 295765
rect 226241 295760 240212 295762
rect 226241 295704 226246 295760
rect 226302 295704 240212 295760
rect 226241 295702 240212 295704
rect 279956 295760 285831 295762
rect 279956 295704 285770 295760
rect 285826 295704 285831 295760
rect 279956 295702 285831 295704
rect 226241 295699 226307 295702
rect 285765 295699 285831 295702
rect 217358 295354 217364 295356
rect 110094 295294 217364 295354
rect 110094 295286 110154 295294
rect 217358 295292 217364 295294
rect 217428 295292 217434 295356
rect 283557 295354 283623 295357
rect 287145 295354 287211 295357
rect 283557 295352 287211 295354
rect 283557 295296 283562 295352
rect 283618 295296 287150 295352
rect 287206 295296 287211 295352
rect 283557 295294 287211 295296
rect 283557 295291 283623 295294
rect 287145 295291 287211 295294
rect 109940 295226 110154 295286
rect 287145 295218 287211 295221
rect 279956 295216 287211 295218
rect 279956 295160 287150 295216
rect 287206 295160 287211 295216
rect 279956 295158 287211 295160
rect 287145 295155 287211 295158
rect 300485 294946 300551 294949
rect 300485 294944 360210 294946
rect 300485 294888 300490 294944
rect 300546 294888 360210 294944
rect 300485 294886 360210 294888
rect 300485 294883 300551 294886
rect 360150 294848 360210 294886
rect 237833 294674 237899 294677
rect 284385 294674 284451 294677
rect 237833 294672 240212 294674
rect 237833 294616 237838 294672
rect 237894 294616 240212 294672
rect 237833 294614 240212 294616
rect 279956 294672 284451 294674
rect 279956 294616 284390 294672
rect 284446 294616 284451 294672
rect 279956 294614 284451 294616
rect 237833 294611 237899 294614
rect 284385 294611 284451 294614
rect 291285 294130 291351 294133
rect 279956 294128 291351 294130
rect 279956 294072 291290 294128
rect 291346 294072 291351 294128
rect 279956 294070 291351 294072
rect 291285 294067 291351 294070
rect 358353 293858 358419 293861
rect 358353 293856 360210 293858
rect 358353 293800 358358 293856
rect 358414 293800 360210 293856
rect 358353 293798 360210 293800
rect 358353 293795 358419 293798
rect 360150 293760 360210 293798
rect 220302 293722 220308 293724
rect 110462 293662 220308 293722
rect 110462 293654 110522 293662
rect 220302 293660 220308 293662
rect 220372 293660 220378 293724
rect 109940 293594 110522 293654
rect 224769 293586 224835 293589
rect 283005 293586 283071 293589
rect 224769 293584 240212 293586
rect 224769 293528 224774 293584
rect 224830 293528 240212 293584
rect 224769 293526 240212 293528
rect 279956 293584 283071 293586
rect 279956 293528 283010 293584
rect 283066 293528 283071 293584
rect 279956 293526 283071 293528
rect 224769 293523 224835 293526
rect 283005 293523 283071 293526
rect -960 293178 480 293268
rect 3366 293178 3372 293180
rect -960 293118 3372 293178
rect -960 293028 480 293118
rect 3366 293116 3372 293118
rect 3436 293116 3442 293180
rect 281809 293042 281875 293045
rect 279956 293040 281875 293042
rect 279956 292984 281814 293040
rect 281870 292984 281875 293040
rect 279956 292982 281875 292984
rect 281809 292979 281875 292982
rect 303245 292770 303311 292773
rect 303245 292768 360210 292770
rect 303245 292712 303250 292768
rect 303306 292712 360210 292768
rect 303245 292710 360210 292712
rect 303245 292707 303311 292710
rect 360150 292672 360210 292710
rect 331949 292634 332015 292637
rect 334801 292634 334867 292637
rect 331949 292632 334867 292634
rect 331949 292576 331954 292632
rect 332010 292576 334806 292632
rect 334862 292576 334867 292632
rect 331949 292574 334867 292576
rect 331949 292571 332015 292574
rect 334801 292571 334867 292574
rect 223389 292498 223455 292501
rect 281901 292498 281967 292501
rect 223389 292496 240212 292498
rect 223389 292440 223394 292496
rect 223450 292440 240212 292496
rect 223389 292438 240212 292440
rect 279956 292496 281967 292498
rect 279956 292440 281906 292496
rect 281962 292440 281967 292496
rect 279956 292438 281967 292440
rect 223389 292435 223455 292438
rect 281901 292435 281967 292438
rect 503621 292226 503687 292229
rect 499806 292224 503687 292226
rect 499806 292168 503626 292224
rect 503682 292168 503687 292224
rect 499806 292166 503687 292168
rect 227345 292090 227411 292093
rect 110462 292088 227411 292090
rect 110462 292032 227350 292088
rect 227406 292032 227411 292088
rect 110462 292030 227411 292032
rect 110462 292022 110522 292030
rect 227345 292027 227411 292030
rect 109940 291962 110522 292022
rect 283189 291954 283255 291957
rect 279956 291952 283255 291954
rect 279956 291896 283194 291952
rect 283250 291896 283255 291952
rect 279956 291894 283255 291896
rect 283189 291891 283255 291894
rect 499806 291856 499866 292166
rect 503621 292163 503687 292166
rect 110413 291818 110479 291821
rect 112437 291818 112503 291821
rect 110413 291816 112503 291818
rect 110413 291760 110418 291816
rect 110474 291760 112442 291816
rect 112498 291760 112503 291816
rect 110413 291758 112503 291760
rect 110413 291755 110479 291758
rect 112437 291755 112503 291758
rect 315481 291682 315547 291685
rect 315481 291680 360210 291682
rect 315481 291624 315486 291680
rect 315542 291624 360210 291680
rect 315481 291622 360210 291624
rect 315481 291619 315547 291622
rect 360150 291584 360210 291622
rect 229001 291410 229067 291413
rect 284518 291410 284524 291412
rect 229001 291408 240212 291410
rect 229001 291352 229006 291408
rect 229062 291352 240212 291408
rect 229001 291350 240212 291352
rect 279956 291350 284524 291410
rect 229001 291347 229067 291350
rect 284518 291348 284524 291350
rect 284588 291348 284594 291412
rect 329925 291138 329991 291141
rect 332041 291138 332107 291141
rect 329925 291136 332107 291138
rect 329925 291080 329930 291136
rect 329986 291080 332046 291136
rect 332102 291080 332107 291136
rect 329925 291078 332107 291080
rect 329925 291075 329991 291078
rect 332041 291075 332107 291078
rect 281901 290866 281967 290869
rect 279956 290864 281967 290866
rect 279956 290808 281906 290864
rect 281962 290808 281967 290864
rect 279956 290806 281967 290808
rect 281901 290803 281967 290806
rect 283649 290594 283715 290597
rect 283649 290592 360210 290594
rect 283649 290536 283654 290592
rect 283710 290536 360210 290592
rect 283649 290534 360210 290536
rect 283649 290531 283715 290534
rect 360150 290496 360210 290534
rect 220486 290458 220492 290460
rect 110462 290398 220492 290458
rect 110462 290390 110522 290398
rect 220486 290396 220492 290398
rect 220556 290396 220562 290460
rect 109940 290330 110522 290390
rect 223481 290322 223547 290325
rect 283097 290322 283163 290325
rect 223481 290320 240212 290322
rect 223481 290264 223486 290320
rect 223542 290264 240212 290320
rect 223481 290262 240212 290264
rect 279956 290320 283163 290322
rect 279956 290264 283102 290320
rect 283158 290264 283163 290320
rect 279956 290262 283163 290264
rect 223481 290259 223547 290262
rect 283097 290259 283163 290262
rect 225965 289778 226031 289781
rect 226190 289778 226196 289780
rect 225965 289776 226196 289778
rect 225965 289720 225970 289776
rect 226026 289720 226196 289776
rect 225965 289718 226196 289720
rect 225965 289715 226031 289718
rect 226190 289716 226196 289718
rect 226260 289716 226266 289780
rect 281901 289778 281967 289781
rect 279956 289776 281967 289778
rect 279956 289720 281906 289776
rect 281962 289720 281967 289776
rect 279956 289718 281967 289720
rect 281901 289715 281967 289718
rect 285213 289506 285279 289509
rect 285213 289504 360210 289506
rect 285213 289448 285218 289504
rect 285274 289448 360210 289504
rect 285213 289446 360210 289448
rect 285213 289443 285279 289446
rect 360150 289408 360210 289446
rect 238661 289234 238727 289237
rect 357198 289234 357204 289236
rect 238661 289232 240212 289234
rect 238661 289176 238666 289232
rect 238722 289176 240212 289232
rect 238661 289174 240212 289176
rect 279956 289174 357204 289234
rect 238661 289171 238727 289174
rect 357198 289172 357204 289174
rect 357268 289172 357274 289236
rect 226006 288826 226012 288828
rect 110462 288766 226012 288826
rect 110462 288758 110522 288766
rect 226006 288764 226012 288766
rect 226076 288764 226082 288828
rect 109940 288698 110522 288758
rect 354070 288690 354076 288692
rect 279956 288630 354076 288690
rect 354070 288628 354076 288630
rect 354140 288628 354146 288692
rect 322381 288418 322447 288421
rect 322381 288416 360210 288418
rect 322381 288360 322386 288416
rect 322442 288360 360210 288416
rect 322381 288358 360210 288360
rect 322381 288355 322447 288358
rect 360150 288320 360210 288358
rect 327809 288282 327875 288285
rect 329925 288282 329991 288285
rect 327809 288280 329991 288282
rect 327809 288224 327814 288280
rect 327870 288224 329930 288280
rect 329986 288224 329991 288280
rect 327809 288222 329991 288224
rect 327809 288219 327875 288222
rect 329925 288219 329991 288222
rect 232773 288146 232839 288149
rect 352966 288146 352972 288148
rect 232773 288144 240212 288146
rect 232773 288088 232778 288144
rect 232834 288088 240212 288144
rect 232773 288086 240212 288088
rect 279956 288086 352972 288146
rect 232773 288083 232839 288086
rect 352966 288084 352972 288086
rect 353036 288084 353042 288148
rect 357525 287874 357591 287877
rect 357525 287872 360210 287874
rect 357525 287816 357530 287872
rect 357586 287816 360210 287872
rect 357525 287814 360210 287816
rect 357525 287811 357591 287814
rect 355542 287602 355548 287604
rect 279956 287542 355548 287602
rect 355542 287540 355548 287542
rect 355612 287540 355618 287604
rect 360150 287232 360210 287814
rect 228214 287194 228220 287196
rect 110462 287134 228220 287194
rect 110462 287126 110522 287134
rect 228214 287132 228220 287134
rect 228284 287132 228290 287196
rect 109940 287066 110522 287126
rect 234470 286996 234476 287060
rect 234540 287058 234546 287060
rect 281993 287058 282059 287061
rect 234540 286998 240212 287058
rect 279956 287056 282059 287058
rect 279956 287000 281998 287056
rect 282054 287000 282059 287056
rect 279956 286998 282059 287000
rect 234540 286996 234546 286998
rect 281993 286995 282059 286998
rect 282545 286514 282611 286517
rect 503621 286514 503687 286517
rect 279956 286512 282611 286514
rect 279956 286456 282550 286512
rect 282606 286456 282611 286512
rect 279956 286454 282611 286456
rect 282545 286451 282611 286454
rect 499806 286512 503687 286514
rect 499806 286456 503626 286512
rect 503682 286456 503687 286512
rect 499806 286454 503687 286456
rect 299013 286242 299079 286245
rect 299013 286240 360210 286242
rect 299013 286184 299018 286240
rect 299074 286184 360210 286240
rect 299013 286182 360210 286184
rect 299013 286179 299079 286182
rect 360150 286144 360210 286182
rect 232589 285970 232655 285973
rect 355174 285970 355180 285972
rect 232589 285968 240212 285970
rect 232589 285912 232594 285968
rect 232650 285912 240212 285968
rect 232589 285910 240212 285912
rect 279956 285910 355180 285970
rect 232589 285907 232655 285910
rect 355174 285908 355180 285910
rect 355244 285908 355250 285972
rect 499806 285872 499866 286454
rect 503621 286451 503687 286454
rect 231526 285562 231532 285564
rect 110462 285502 231532 285562
rect 110462 285494 110522 285502
rect 231526 285500 231532 285502
rect 231596 285500 231602 285564
rect 109940 285434 110522 285494
rect 282269 285426 282335 285429
rect 279956 285424 282335 285426
rect 279956 285368 282274 285424
rect 282330 285368 282335 285424
rect 279956 285366 282335 285368
rect 282269 285363 282335 285366
rect 583520 285276 584960 285516
rect 284937 285154 285003 285157
rect 284937 285152 360210 285154
rect 284937 285096 284942 285152
rect 284998 285096 360210 285152
rect 284937 285094 360210 285096
rect 284937 285091 285003 285094
rect 360150 285056 360210 285094
rect 48078 284956 48084 285020
rect 48148 285018 48154 285020
rect 48148 284958 50140 285018
rect 48148 284956 48154 284958
rect 234286 284820 234292 284884
rect 234356 284882 234362 284884
rect 282085 284882 282151 284885
rect 234356 284822 240212 284882
rect 279956 284880 282151 284882
rect 279956 284824 282090 284880
rect 282146 284824 282151 284880
rect 279956 284822 282151 284824
rect 234356 284820 234362 284822
rect 282085 284819 282151 284822
rect 354254 284338 354260 284340
rect 279956 284278 354260 284338
rect 354254 284276 354260 284278
rect 354324 284276 354330 284340
rect 293493 284066 293559 284069
rect 293493 284064 360210 284066
rect 293493 284008 293498 284064
rect 293554 284008 360210 284064
rect 293493 284006 360210 284008
rect 293493 284003 293559 284006
rect 360150 283968 360210 284006
rect 227069 283930 227135 283933
rect 110462 283928 227135 283930
rect 110462 283872 227074 283928
rect 227130 283872 227135 283928
rect 110462 283870 227135 283872
rect 110462 283862 110522 283870
rect 227069 283867 227135 283870
rect 109940 283802 110522 283862
rect 235758 283732 235764 283796
rect 235828 283794 235834 283796
rect 282453 283794 282519 283797
rect 235828 283734 240212 283794
rect 279956 283792 282519 283794
rect 279956 283736 282458 283792
rect 282514 283736 282519 283792
rect 279956 283734 282519 283736
rect 235828 283732 235834 283734
rect 282453 283731 282519 283734
rect 356830 283250 356836 283252
rect 279956 283190 356836 283250
rect 356830 283188 356836 283190
rect 356900 283188 356906 283252
rect 318241 282842 318307 282845
rect 360150 282842 360210 282880
rect 318241 282840 360210 282842
rect 318241 282784 318246 282840
rect 318302 282784 360210 282840
rect 318241 282782 360210 282784
rect 318241 282779 318307 282782
rect 233693 282706 233759 282709
rect 282821 282706 282887 282709
rect 233693 282704 240212 282706
rect 233693 282648 233698 282704
rect 233754 282648 240212 282704
rect 233693 282646 240212 282648
rect 279956 282704 282887 282706
rect 279956 282648 282826 282704
rect 282882 282648 282887 282704
rect 279956 282646 282887 282648
rect 233693 282643 233759 282646
rect 282821 282643 282887 282646
rect 224902 282434 224908 282436
rect 219390 282374 224908 282434
rect 219390 282298 219450 282374
rect 224902 282372 224908 282374
rect 224972 282372 224978 282436
rect 110462 282238 219450 282298
rect 110462 282230 110522 282238
rect 224902 282236 224908 282300
rect 224972 282298 224978 282300
rect 226057 282298 226123 282301
rect 224972 282296 226123 282298
rect 224972 282240 226062 282296
rect 226118 282240 226123 282296
rect 224972 282238 226123 282240
rect 224972 282236 224978 282238
rect 226057 282235 226123 282238
rect 330477 282298 330543 282301
rect 331949 282298 332015 282301
rect 330477 282296 332015 282298
rect 330477 282240 330482 282296
rect 330538 282240 331954 282296
rect 332010 282240 332015 282296
rect 330477 282238 332015 282240
rect 330477 282235 330543 282238
rect 331949 282235 332015 282238
rect 357525 282298 357591 282301
rect 357525 282296 360210 282298
rect 357525 282240 357530 282296
rect 357586 282240 360210 282296
rect 357525 282238 360210 282240
rect 357525 282235 357591 282238
rect 109940 282170 110522 282230
rect 358118 282162 358124 282164
rect 279956 282102 358124 282162
rect 358118 282100 358124 282102
rect 358188 282100 358194 282164
rect 360150 281792 360210 282238
rect 233877 281618 233943 281621
rect 282177 281618 282243 281621
rect 233877 281616 240212 281618
rect 233877 281560 233882 281616
rect 233938 281560 240212 281616
rect 233877 281558 240212 281560
rect 279956 281616 282243 281618
rect 279956 281560 282182 281616
rect 282238 281560 282243 281616
rect 279956 281558 282243 281560
rect 233877 281555 233943 281558
rect 282177 281555 282243 281558
rect 349838 281074 349844 281076
rect 279956 281014 349844 281074
rect 349838 281012 349844 281014
rect 349908 281012 349914 281076
rect 319621 280802 319687 280805
rect 319621 280800 360210 280802
rect 319621 280744 319626 280800
rect 319682 280744 360210 280800
rect 319621 280742 360210 280744
rect 319621 280739 319687 280742
rect 360150 280704 360210 280742
rect 222878 280666 222884 280668
rect 110462 280606 222884 280666
rect 110462 280598 110522 280606
rect 222878 280604 222884 280606
rect 222948 280604 222954 280668
rect 354438 280666 354444 280668
rect 335310 280606 354444 280666
rect 109940 280538 110522 280598
rect 238385 280530 238451 280533
rect 335310 280530 335370 280606
rect 354438 280604 354444 280606
rect 354508 280604 354514 280668
rect 238385 280528 240212 280530
rect 238385 280472 238390 280528
rect 238446 280472 240212 280528
rect 238385 280470 240212 280472
rect 279956 280470 335370 280530
rect 238385 280467 238451 280470
rect -960 279972 480 280212
rect 282361 279986 282427 279989
rect 518934 279986 518940 279988
rect 279956 279984 282427 279986
rect 279956 279928 282366 279984
rect 282422 279928 282427 279984
rect 279956 279926 282427 279928
rect 282361 279923 282427 279926
rect 499806 279926 518940 279986
rect 499806 279888 499866 279926
rect 518934 279924 518940 279926
rect 519004 279924 519010 279988
rect 311433 279714 311499 279717
rect 311433 279712 360210 279714
rect 311433 279656 311438 279712
rect 311494 279656 360210 279712
rect 311433 279654 360210 279656
rect 311433 279651 311499 279654
rect 360150 279616 360210 279654
rect 233785 279442 233851 279445
rect 353886 279442 353892 279444
rect 233785 279440 240212 279442
rect 233785 279384 233790 279440
rect 233846 279384 240212 279440
rect 233785 279382 240212 279384
rect 279956 279382 353892 279442
rect 233785 279379 233851 279382
rect 353886 279380 353892 279382
rect 353956 279380 353962 279444
rect 227161 279034 227227 279037
rect 110462 279032 227227 279034
rect 110462 278976 227166 279032
rect 227222 278976 227227 279032
rect 110462 278974 227227 278976
rect 110462 278966 110522 278974
rect 227161 278971 227227 278974
rect 109940 278906 110522 278966
rect 282729 278898 282795 278901
rect 279956 278896 282795 278898
rect 279956 278840 282734 278896
rect 282790 278840 282795 278896
rect 279956 278838 282795 278840
rect 282729 278835 282795 278838
rect 308581 278626 308647 278629
rect 308581 278624 360210 278626
rect 308581 278568 308586 278624
rect 308642 278568 360210 278624
rect 308581 278566 360210 278568
rect 308581 278563 308647 278566
rect 360150 278528 360210 278566
rect 234153 278354 234219 278357
rect 338614 278354 338620 278356
rect 234153 278352 240212 278354
rect 234153 278296 234158 278352
rect 234214 278296 240212 278352
rect 234153 278294 240212 278296
rect 279956 278294 338620 278354
rect 234153 278291 234219 278294
rect 338614 278292 338620 278294
rect 338684 278292 338690 278356
rect 282637 277810 282703 277813
rect 279956 277808 282703 277810
rect 279956 277752 282642 277808
rect 282698 277752 282703 277808
rect 279956 277750 282703 277752
rect 282637 277747 282703 277750
rect 329097 277538 329163 277541
rect 329097 277536 360210 277538
rect 329097 277480 329102 277536
rect 329158 277480 360210 277536
rect 329097 277478 360210 277480
rect 329097 277475 329163 277478
rect 360150 277440 360210 277478
rect 226977 277402 227043 277405
rect 110462 277400 227043 277402
rect 110462 277344 226982 277400
rect 227038 277344 227043 277400
rect 110462 277342 227043 277344
rect 110462 277334 110522 277342
rect 226977 277339 227043 277342
rect 109940 277274 110522 277334
rect 234337 277266 234403 277269
rect 356646 277266 356652 277268
rect 234337 277264 240212 277266
rect 234337 277208 234342 277264
rect 234398 277208 240212 277264
rect 234337 277206 240212 277208
rect 279956 277206 356652 277266
rect 234337 277203 234403 277206
rect 356646 277204 356652 277206
rect 356716 277204 356722 277268
rect 357525 276858 357591 276861
rect 357525 276856 360210 276858
rect 357525 276800 357530 276856
rect 357586 276800 360210 276856
rect 357525 276798 360210 276800
rect 357525 276795 357591 276798
rect 351126 276722 351132 276724
rect 279956 276662 351132 276722
rect 351126 276660 351132 276662
rect 351196 276660 351202 276724
rect 360150 276352 360210 276798
rect 542854 276660 542860 276724
rect 542924 276722 542930 276724
rect 580390 276722 580396 276724
rect 542924 276662 580396 276722
rect 542924 276660 542930 276662
rect 580390 276660 580396 276662
rect 580460 276660 580466 276724
rect 235165 276178 235231 276181
rect 346894 276178 346900 276180
rect 235165 276176 240212 276178
rect 235165 276120 235170 276176
rect 235226 276120 240212 276176
rect 235165 276118 240212 276120
rect 279956 276118 346900 276178
rect 235165 276115 235231 276118
rect 346894 276116 346900 276118
rect 346964 276116 346970 276180
rect 220118 275770 220124 275772
rect 110462 275710 220124 275770
rect 110462 275702 110522 275710
rect 220118 275708 220124 275710
rect 220188 275708 220194 275772
rect 109940 275642 110522 275702
rect 349654 275634 349660 275636
rect 279956 275574 349660 275634
rect 349654 275572 349660 275574
rect 349724 275572 349730 275636
rect 112437 275362 112503 275365
rect 113909 275362 113975 275365
rect 112437 275360 113975 275362
rect 112437 275304 112442 275360
rect 112498 275304 113914 275360
rect 113970 275304 113975 275360
rect 112437 275302 113975 275304
rect 112437 275299 112503 275302
rect 113909 275299 113975 275302
rect 309869 275362 309935 275365
rect 309869 275360 360210 275362
rect 309869 275304 309874 275360
rect 309930 275304 360210 275360
rect 309869 275302 360210 275304
rect 309869 275299 309935 275302
rect 360150 275264 360210 275302
rect 233601 275090 233667 275093
rect 351310 275090 351316 275092
rect 233601 275088 240212 275090
rect 233601 275032 233606 275088
rect 233662 275032 240212 275088
rect 233601 275030 240212 275032
rect 279956 275030 351316 275090
rect 233601 275027 233667 275030
rect 351310 275028 351316 275030
rect 351380 275028 351386 275092
rect 329097 274682 329163 274685
rect 330477 274682 330543 274685
rect 329097 274680 330543 274682
rect 329097 274624 329102 274680
rect 329158 274624 330482 274680
rect 330538 274624 330543 274680
rect 329097 274622 330543 274624
rect 329097 274619 329163 274622
rect 330477 274619 330543 274622
rect 282310 274546 282316 274548
rect 279956 274486 282316 274546
rect 282310 274484 282316 274486
rect 282380 274484 282386 274548
rect 297449 274274 297515 274277
rect 503621 274274 503687 274277
rect 297449 274272 360210 274274
rect 297449 274216 297454 274272
rect 297510 274216 360210 274272
rect 297449 274214 360210 274216
rect 297449 274211 297515 274214
rect 360150 274176 360210 274214
rect 499806 274272 503687 274274
rect 499806 274216 503626 274272
rect 503682 274216 503687 274272
rect 499806 274214 503687 274216
rect 227478 274138 227484 274140
rect 110462 274078 227484 274138
rect 110462 274070 110522 274078
rect 227478 274076 227484 274078
rect 227548 274076 227554 274140
rect 109940 274010 110522 274070
rect 234061 274002 234127 274005
rect 352782 274002 352788 274004
rect 234061 274000 240212 274002
rect 234061 273944 234066 274000
rect 234122 273944 240212 274000
rect 234061 273942 240212 273944
rect 279956 273942 352788 274002
rect 234061 273939 234127 273942
rect 352782 273940 352788 273942
rect 352852 273940 352858 274004
rect 499806 273904 499866 274214
rect 503621 274211 503687 274214
rect 282678 273458 282684 273460
rect 279956 273398 282684 273458
rect 282678 273396 282684 273398
rect 282748 273396 282754 273460
rect 320909 273186 320975 273189
rect 320909 273184 360210 273186
rect 320909 273128 320914 273184
rect 320970 273128 360210 273184
rect 320909 273126 360210 273128
rect 320909 273123 320975 273126
rect 360150 273088 360210 273126
rect 325877 273050 325943 273053
rect 327809 273050 327875 273053
rect 325877 273048 327875 273050
rect 325877 272992 325882 273048
rect 325938 272992 327814 273048
rect 327870 272992 327875 273048
rect 325877 272990 327875 272992
rect 325877 272987 325943 272990
rect 327809 272987 327875 272990
rect 234245 272914 234311 272917
rect 357014 272914 357020 272916
rect 234245 272912 240212 272914
rect 234245 272856 234250 272912
rect 234306 272856 240212 272912
rect 234245 272854 240212 272856
rect 279956 272854 357020 272914
rect 234245 272851 234311 272854
rect 357014 272852 357020 272854
rect 357084 272852 357090 272916
rect 357525 272642 357591 272645
rect 357525 272640 360210 272642
rect 357525 272584 357530 272640
rect 357586 272584 360210 272640
rect 357525 272582 360210 272584
rect 357525 272579 357591 272582
rect 226926 272506 226932 272508
rect 110462 272446 226932 272506
rect 110462 272438 110522 272446
rect 226926 272444 226932 272446
rect 226996 272444 227002 272508
rect 109940 272378 110522 272438
rect 282126 272370 282132 272372
rect 279956 272310 282132 272370
rect 282126 272308 282132 272310
rect 282196 272308 282202 272372
rect 360150 272000 360210 272582
rect 580257 272234 580323 272237
rect 583520 272234 584960 272324
rect 580257 272232 584960 272234
rect 580257 272176 580262 272232
rect 580318 272176 584960 272232
rect 580257 272174 584960 272176
rect 580257 272171 580323 272174
rect 583520 272084 584960 272174
rect 237281 271826 237347 271829
rect 355358 271826 355364 271828
rect 237281 271824 240212 271826
rect 237281 271768 237286 271824
rect 237342 271768 240212 271824
rect 237281 271766 240212 271768
rect 279956 271766 355364 271826
rect 237281 271763 237347 271766
rect 355358 271764 355364 271766
rect 355428 271764 355434 271828
rect 357525 271418 357591 271421
rect 357525 271416 360210 271418
rect 357525 271360 357530 271416
rect 357586 271360 360210 271416
rect 357525 271358 360210 271360
rect 357525 271355 357591 271358
rect 357934 271282 357940 271284
rect 279956 271222 357940 271282
rect 357934 271220 357940 271222
rect 358004 271220 358010 271284
rect 360150 270912 360210 271358
rect 227110 270874 227116 270876
rect 110462 270814 227116 270874
rect 110462 270806 110522 270814
rect 227110 270812 227116 270814
rect 227180 270812 227186 270876
rect 109940 270746 110522 270806
rect 235073 270738 235139 270741
rect 282494 270738 282500 270740
rect 235073 270736 240212 270738
rect 235073 270680 235078 270736
rect 235134 270680 240212 270736
rect 235073 270678 240212 270680
rect 279956 270678 282500 270738
rect 235073 270675 235139 270678
rect 282494 270676 282500 270678
rect 282564 270676 282570 270740
rect 345606 270194 345612 270196
rect 279956 270134 345612 270194
rect 345606 270132 345612 270134
rect 345676 270132 345682 270196
rect 357525 270194 357591 270197
rect 357525 270192 360210 270194
rect 357525 270136 357530 270192
rect 357586 270136 360210 270192
rect 357525 270134 360210 270136
rect 357525 270131 357591 270134
rect 360150 269824 360210 270134
rect 235625 269650 235691 269653
rect 296989 269650 297055 269653
rect 235625 269648 240212 269650
rect 235625 269592 235630 269648
rect 235686 269592 240212 269648
rect 235625 269590 240212 269592
rect 279956 269648 297055 269650
rect 279956 269592 296994 269648
rect 297050 269592 297055 269648
rect 279956 269590 297055 269592
rect 235625 269587 235691 269590
rect 296989 269587 297055 269590
rect 227294 269242 227300 269244
rect 110462 269182 227300 269242
rect 110462 269174 110522 269182
rect 227294 269180 227300 269182
rect 227364 269180 227370 269244
rect 109940 269114 110522 269174
rect 282085 269106 282151 269109
rect 279956 269104 282151 269106
rect 279956 269048 282090 269104
rect 282146 269048 282151 269104
rect 279956 269046 282151 269048
rect 282085 269043 282151 269046
rect 301589 268834 301655 268837
rect 301589 268832 360210 268834
rect 301589 268776 301594 268832
rect 301650 268776 360210 268832
rect 301589 268774 360210 268776
rect 301589 268771 301655 268774
rect 360150 268736 360210 268774
rect 237189 268562 237255 268565
rect 280153 268562 280219 268565
rect 237189 268560 240212 268562
rect 237189 268504 237194 268560
rect 237250 268504 240212 268560
rect 237189 268502 240212 268504
rect 279956 268560 280219 268562
rect 279956 268504 280158 268560
rect 280214 268504 280219 268560
rect 279956 268502 280219 268504
rect 237189 268499 237255 268502
rect 280153 268499 280219 268502
rect 282821 268018 282887 268021
rect 518198 268018 518204 268020
rect 279956 268016 282887 268018
rect 279956 267960 282826 268016
rect 282882 267960 282887 268016
rect 279956 267958 282887 267960
rect 282821 267955 282887 267958
rect 499806 267958 518204 268018
rect 499806 267920 499866 267958
rect 518198 267956 518204 267958
rect 518268 267956 518274 268020
rect 292021 267746 292087 267749
rect 292021 267744 360210 267746
rect 292021 267688 292026 267744
rect 292082 267688 360210 267744
rect 292021 267686 360210 267688
rect 292021 267683 292087 267686
rect 360150 267648 360210 267686
rect 231342 267610 231348 267612
rect 110462 267550 231348 267610
rect 110462 267542 110522 267550
rect 231342 267548 231348 267550
rect 231412 267548 231418 267612
rect 109940 267482 110522 267542
rect 235717 267474 235783 267477
rect 294137 267474 294203 267477
rect 235717 267472 240212 267474
rect 235717 267416 235722 267472
rect 235778 267416 240212 267472
rect 235717 267414 240212 267416
rect 279956 267472 294203 267474
rect 279956 267416 294142 267472
rect 294198 267416 294203 267472
rect 279956 267414 294203 267416
rect 235717 267411 235783 267414
rect 294137 267411 294203 267414
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 285949 266930 286015 266933
rect 279956 266928 286015 266930
rect 279956 266872 285954 266928
rect 286010 266872 286015 266928
rect 279956 266870 286015 266872
rect 285949 266867 286015 266870
rect 294873 266658 294939 266661
rect 294873 266656 360210 266658
rect 294873 266600 294878 266656
rect 294934 266600 360210 266656
rect 294873 266598 360210 266600
rect 294873 266595 294939 266598
rect 360150 266560 360210 266598
rect 235533 266386 235599 266389
rect 283465 266386 283531 266389
rect 235533 266384 240212 266386
rect 235533 266328 235538 266384
rect 235594 266328 240212 266384
rect 235533 266326 240212 266328
rect 279956 266384 283531 266386
rect 279956 266328 283470 266384
rect 283526 266328 283531 266384
rect 279956 266326 283531 266328
rect 235533 266323 235599 266326
rect 283465 266323 283531 266326
rect 211654 265978 211660 265980
rect 110462 265918 211660 265978
rect 110462 265910 110522 265918
rect 211654 265916 211660 265918
rect 211724 265916 211730 265980
rect 109940 265850 110522 265910
rect 294229 265842 294295 265845
rect 279956 265840 294295 265842
rect 279956 265784 294234 265840
rect 294290 265784 294295 265840
rect 279956 265782 294295 265784
rect 294229 265779 294295 265782
rect 296161 265570 296227 265573
rect 296161 265568 360210 265570
rect 296161 265512 296166 265568
rect 296222 265512 360210 265568
rect 296161 265510 360210 265512
rect 296161 265507 296227 265510
rect 360150 265472 360210 265510
rect 235901 265298 235967 265301
rect 282821 265298 282887 265301
rect 235901 265296 240212 265298
rect 235901 265240 235906 265296
rect 235962 265240 240212 265296
rect 235901 265238 240212 265240
rect 279956 265296 282887 265298
rect 279956 265240 282826 265296
rect 282882 265240 282887 265296
rect 279956 265238 282887 265240
rect 235901 265235 235967 265238
rect 282821 265235 282887 265238
rect 113909 265026 113975 265029
rect 115197 265026 115263 265029
rect 113909 265024 115263 265026
rect 113909 264968 113914 265024
rect 113970 264968 115202 265024
rect 115258 264968 115263 265024
rect 113909 264966 115263 264968
rect 113909 264963 113975 264966
rect 115197 264963 115263 264966
rect 301129 264754 301195 264757
rect 279956 264752 301195 264754
rect 279956 264696 301134 264752
rect 301190 264696 301195 264752
rect 279956 264694 301195 264696
rect 301129 264691 301195 264694
rect 307201 264482 307267 264485
rect 307201 264480 360210 264482
rect 307201 264424 307206 264480
rect 307262 264424 360210 264480
rect 307201 264422 360210 264424
rect 307201 264419 307267 264422
rect 360150 264384 360210 264422
rect 215886 264346 215892 264348
rect 110462 264286 215892 264346
rect 110462 264278 110522 264286
rect 215886 264284 215892 264286
rect 215956 264284 215962 264348
rect 109940 264218 110522 264278
rect 235441 264210 235507 264213
rect 282821 264210 282887 264213
rect 235441 264208 240212 264210
rect 235441 264152 235446 264208
rect 235502 264152 240212 264208
rect 235441 264150 240212 264152
rect 279956 264208 282887 264210
rect 279956 264152 282826 264208
rect 282882 264152 282887 264208
rect 279956 264150 282887 264152
rect 235441 264147 235507 264150
rect 282821 264147 282887 264150
rect 295793 263666 295859 263669
rect 279956 263664 295859 263666
rect 279956 263608 295798 263664
rect 295854 263608 295859 263664
rect 279956 263606 295859 263608
rect 295793 263603 295859 263606
rect 320909 263666 320975 263669
rect 325141 263666 325207 263669
rect 320909 263664 325207 263666
rect 320909 263608 320914 263664
rect 320970 263608 325146 263664
rect 325202 263608 325207 263664
rect 320909 263606 325207 263608
rect 320909 263603 320975 263606
rect 325141 263603 325207 263606
rect 288065 263394 288131 263397
rect 288065 263392 360210 263394
rect 288065 263336 288070 263392
rect 288126 263336 360210 263392
rect 288065 263334 360210 263336
rect 288065 263331 288131 263334
rect 360150 263296 360210 263334
rect 235809 263122 235875 263125
rect 282821 263122 282887 263125
rect 235809 263120 240212 263122
rect 235809 263064 235814 263120
rect 235870 263064 240212 263120
rect 235809 263062 240212 263064
rect 279956 263120 282887 263122
rect 279956 263064 282826 263120
rect 282882 263064 282887 263120
rect 279956 263062 282887 263064
rect 235809 263059 235875 263062
rect 282821 263059 282887 263062
rect 216070 262714 216076 262716
rect 110462 262654 216076 262714
rect 110462 262646 110522 262654
rect 216070 262652 216076 262654
rect 216140 262652 216146 262716
rect 109940 262586 110522 262646
rect 282729 262578 282795 262581
rect 279956 262576 282795 262578
rect 279956 262520 282734 262576
rect 282790 262520 282795 262576
rect 279956 262518 282795 262520
rect 282729 262515 282795 262518
rect 293401 262306 293467 262309
rect 293401 262304 360210 262306
rect 293401 262248 293406 262304
rect 293462 262248 360210 262304
rect 293401 262246 360210 262248
rect 293401 262243 293467 262246
rect 360150 262208 360210 262246
rect 235257 262034 235323 262037
rect 282821 262034 282887 262037
rect 518014 262034 518020 262036
rect 235257 262032 240212 262034
rect 235257 261976 235262 262032
rect 235318 261976 240212 262032
rect 235257 261974 240212 261976
rect 279956 262032 282887 262034
rect 279956 261976 282826 262032
rect 282882 261976 282887 262032
rect 279956 261974 282887 261976
rect 235257 261971 235323 261974
rect 282821 261971 282887 261974
rect 499806 261974 518020 262034
rect 499806 261936 499866 261974
rect 518014 261972 518020 261974
rect 518084 261972 518090 262036
rect 357525 261626 357591 261629
rect 357525 261624 360210 261626
rect 357525 261568 357530 261624
rect 357586 261568 360210 261624
rect 357525 261566 360210 261568
rect 357525 261563 357591 261566
rect 302601 261490 302667 261493
rect 279956 261488 302667 261490
rect 279956 261432 302606 261488
rect 302662 261432 302667 261488
rect 279956 261430 302667 261432
rect 302601 261427 302667 261430
rect 360150 261120 360210 261566
rect 224401 261082 224467 261085
rect 110462 261080 224467 261082
rect 110462 261024 224406 261080
rect 224462 261024 224467 261080
rect 110462 261022 224467 261024
rect 110462 261014 110522 261022
rect 224401 261019 224467 261022
rect 109940 260954 110522 261014
rect 235349 260946 235415 260949
rect 283373 260946 283439 260949
rect 235349 260944 240212 260946
rect 235349 260888 235354 260944
rect 235410 260888 240212 260944
rect 235349 260886 240212 260888
rect 279956 260944 283439 260946
rect 279956 260888 283378 260944
rect 283434 260888 283439 260944
rect 279956 260886 283439 260888
rect 235349 260883 235415 260886
rect 283373 260883 283439 260886
rect 290089 260402 290155 260405
rect 279956 260400 290155 260402
rect 279956 260344 290094 260400
rect 290150 260344 290155 260400
rect 279956 260342 290155 260344
rect 290089 260339 290155 260342
rect 284886 260068 284892 260132
rect 284956 260130 284962 260132
rect 284956 260070 360210 260130
rect 284956 260068 284962 260070
rect 360150 260032 360210 260070
rect 234521 259858 234587 259861
rect 282821 259858 282887 259861
rect 234521 259856 240212 259858
rect 234521 259800 234526 259856
rect 234582 259800 240212 259856
rect 234521 259798 240212 259800
rect 279956 259856 282887 259858
rect 279956 259800 282826 259856
rect 282882 259800 282887 259856
rect 279956 259798 282887 259800
rect 234521 259795 234587 259798
rect 282821 259795 282887 259798
rect 224217 259450 224283 259453
rect 110462 259448 224283 259450
rect 110462 259392 224222 259448
rect 224278 259392 224283 259448
rect 110462 259390 224283 259392
rect 110462 259382 110522 259390
rect 224217 259387 224283 259390
rect 109940 259322 110522 259382
rect 282821 259314 282887 259317
rect 279956 259312 282887 259314
rect 279956 259256 282826 259312
rect 282882 259256 282887 259312
rect 279956 259254 282887 259256
rect 282821 259251 282887 259254
rect 305729 259042 305795 259045
rect 305729 259040 360210 259042
rect 305729 258984 305734 259040
rect 305790 258984 360210 259040
rect 305729 258982 360210 258984
rect 305729 258979 305795 258982
rect 360150 258944 360210 258982
rect 508446 258844 508452 258908
rect 508516 258906 508522 258908
rect 583520 258906 584960 258996
rect 508516 258846 584960 258906
rect 508516 258844 508522 258846
rect 233049 258770 233115 258773
rect 282637 258770 282703 258773
rect 233049 258768 240212 258770
rect 233049 258712 233054 258768
rect 233110 258712 240212 258768
rect 233049 258710 240212 258712
rect 279956 258768 282703 258770
rect 279956 258712 282642 258768
rect 282698 258712 282703 258768
rect 583520 258756 584960 258846
rect 279956 258710 282703 258712
rect 233049 258707 233115 258710
rect 282637 258707 282703 258710
rect 282729 258226 282795 258229
rect 279956 258224 282795 258226
rect 279956 258168 282734 258224
rect 282790 258168 282795 258224
rect 279956 258166 282795 258168
rect 282729 258163 282795 258166
rect 323669 257954 323735 257957
rect 323669 257952 360210 257954
rect 323669 257896 323674 257952
rect 323730 257896 360210 257952
rect 323669 257894 360210 257896
rect 323669 257891 323735 257894
rect 360150 257856 360210 257894
rect 224350 257818 224356 257820
rect 110462 257758 224356 257818
rect 110462 257750 110522 257758
rect 224350 257756 224356 257758
rect 224420 257756 224426 257820
rect 109940 257690 110522 257750
rect 232957 257682 233023 257685
rect 282821 257682 282887 257685
rect 232957 257680 240212 257682
rect 232957 257624 232962 257680
rect 233018 257624 240212 257680
rect 232957 257622 240212 257624
rect 279956 257680 282887 257682
rect 279956 257624 282826 257680
rect 282882 257624 282887 257680
rect 279956 257622 282887 257624
rect 232957 257619 233023 257622
rect 282821 257619 282887 257622
rect 282729 257138 282795 257141
rect 279956 257136 282795 257138
rect 279956 257080 282734 257136
rect 282790 257080 282795 257136
rect 279956 257078 282795 257080
rect 282729 257075 282795 257078
rect 314193 256866 314259 256869
rect 314193 256864 360210 256866
rect 314193 256808 314198 256864
rect 314254 256808 360210 256864
rect 314193 256806 360210 256808
rect 314193 256803 314259 256806
rect 360150 256768 360210 256806
rect 223614 256668 223620 256732
rect 223684 256730 223690 256732
rect 224677 256730 224743 256733
rect 503897 256730 503963 256733
rect 223684 256728 224743 256730
rect 223684 256672 224682 256728
rect 224738 256672 224743 256728
rect 223684 256670 224743 256672
rect 223684 256668 223690 256670
rect 224677 256667 224743 256670
rect 503670 256728 503963 256730
rect 503670 256672 503902 256728
rect 503958 256672 503963 256728
rect 503670 256670 503963 256672
rect 232865 256594 232931 256597
rect 282821 256594 282887 256597
rect 503670 256594 503730 256670
rect 503897 256667 503963 256670
rect 232865 256592 240212 256594
rect 232865 256536 232870 256592
rect 232926 256536 240212 256592
rect 232865 256534 240212 256536
rect 279956 256592 282887 256594
rect 279956 256536 282826 256592
rect 282882 256536 282887 256592
rect 279956 256534 282887 256536
rect 232865 256531 232931 256534
rect 282821 256531 282887 256534
rect 499806 256534 503730 256594
rect 221038 256186 221044 256188
rect 110462 256126 221044 256186
rect 110462 256118 110522 256126
rect 221038 256124 221044 256126
rect 221108 256124 221114 256188
rect 357525 256186 357591 256189
rect 357525 256184 360210 256186
rect 357525 256128 357530 256184
rect 357586 256128 360210 256184
rect 357525 256126 360210 256128
rect 357525 256123 357591 256126
rect 109940 256058 110522 256118
rect 282637 256050 282703 256053
rect 279956 256048 282703 256050
rect 279956 255992 282642 256048
rect 282698 255992 282703 256048
rect 279956 255990 282703 255992
rect 282637 255987 282703 255990
rect 360150 255680 360210 256126
rect 499806 255952 499866 256534
rect 232681 255506 232747 255509
rect 282729 255506 282795 255509
rect 232681 255504 240212 255506
rect 232681 255448 232686 255504
rect 232742 255448 240212 255504
rect 232681 255446 240212 255448
rect 279956 255504 282795 255506
rect 279956 255448 282734 255504
rect 282790 255448 282795 255504
rect 279956 255446 282795 255448
rect 232681 255443 232747 255446
rect 282729 255443 282795 255446
rect 220854 255308 220860 255372
rect 220924 255370 220930 255372
rect 222101 255370 222167 255373
rect 220924 255368 222167 255370
rect 220924 255312 222106 255368
rect 222162 255312 222167 255368
rect 220924 255310 222167 255312
rect 220924 255308 220930 255310
rect 222101 255307 222167 255310
rect 319621 255370 319687 255373
rect 320909 255370 320975 255373
rect 319621 255368 320975 255370
rect 319621 255312 319626 255368
rect 319682 255312 320914 255368
rect 320970 255312 320975 255368
rect 319621 255310 320975 255312
rect 319621 255307 319687 255310
rect 320909 255307 320975 255310
rect 48221 255098 48287 255101
rect 48221 255096 50140 255098
rect 48221 255040 48226 255096
rect 48282 255040 50140 255096
rect 48221 255038 50140 255040
rect 48221 255035 48287 255038
rect 304993 254962 305059 254965
rect 279956 254960 305059 254962
rect 279956 254904 304998 254960
rect 305054 254904 305059 254960
rect 279956 254902 305059 254904
rect 304993 254899 305059 254902
rect 357525 254962 357591 254965
rect 357525 254960 360210 254962
rect 357525 254904 357530 254960
rect 357586 254904 360210 254960
rect 357525 254902 360210 254904
rect 357525 254899 357591 254902
rect 360150 254592 360210 254902
rect 224534 254554 224540 254556
rect 109940 254494 224540 254554
rect 224534 254492 224540 254494
rect 224604 254492 224610 254556
rect 233969 254418 234035 254421
rect 282821 254418 282887 254421
rect 233969 254416 240212 254418
rect 233969 254360 233974 254416
rect 234030 254360 240212 254416
rect 233969 254358 240212 254360
rect 279956 254416 282887 254418
rect 279956 254360 282826 254416
rect 282882 254360 282887 254416
rect 279956 254358 282887 254360
rect 233969 254355 234035 254358
rect 282821 254355 282887 254358
rect -960 254146 480 254236
rect 48630 254146 48636 254148
rect -960 254086 48636 254146
rect -960 253996 480 254086
rect 48630 254084 48636 254086
rect 48700 254084 48706 254148
rect 223798 253948 223804 254012
rect 223868 254010 223874 254012
rect 224861 254010 224927 254013
rect 223868 254008 224927 254010
rect 223868 253952 224866 254008
rect 224922 253952 224927 254008
rect 223868 253950 224927 253952
rect 223868 253948 223874 253950
rect 224861 253947 224927 253950
rect 282821 253874 282887 253877
rect 279956 253872 282887 253874
rect 279956 253816 282826 253872
rect 282882 253816 282887 253872
rect 279956 253814 282887 253816
rect 282821 253811 282887 253814
rect 326981 253874 327047 253877
rect 329097 253874 329163 253877
rect 326981 253872 329163 253874
rect 326981 253816 326986 253872
rect 327042 253816 329102 253872
rect 329158 253816 329163 253872
rect 326981 253814 329163 253816
rect 326981 253811 327047 253814
rect 329097 253811 329163 253814
rect 304441 253602 304507 253605
rect 304441 253600 360210 253602
rect 304441 253544 304446 253600
rect 304502 253544 360210 253600
rect 304441 253542 360210 253544
rect 304441 253539 304507 253542
rect 360150 253504 360210 253542
rect 236361 253330 236427 253333
rect 282637 253330 282703 253333
rect 236361 253328 240212 253330
rect 236361 253272 236366 253328
rect 236422 253272 240212 253328
rect 236361 253270 240212 253272
rect 279956 253328 282703 253330
rect 279956 253272 282642 253328
rect 282698 253272 282703 253328
rect 279956 253270 282703 253272
rect 236361 253267 236427 253270
rect 282637 253267 282703 253270
rect 224718 252922 224724 252924
rect 110462 252862 224724 252922
rect 110462 252854 110522 252862
rect 224718 252860 224724 252862
rect 224788 252860 224794 252924
rect 109940 252794 110522 252854
rect 282729 252786 282795 252789
rect 279956 252784 282795 252786
rect 279956 252728 282734 252784
rect 282790 252728 282795 252784
rect 279956 252726 282795 252728
rect 282729 252723 282795 252726
rect 230054 252452 230060 252516
rect 230124 252514 230130 252516
rect 230289 252514 230355 252517
rect 230124 252512 230355 252514
rect 230124 252456 230294 252512
rect 230350 252456 230355 252512
rect 230124 252454 230355 252456
rect 230124 252452 230130 252454
rect 230289 252451 230355 252454
rect 303153 252514 303219 252517
rect 303153 252512 360210 252514
rect 303153 252456 303158 252512
rect 303214 252456 360210 252512
rect 303153 252454 360210 252456
rect 303153 252451 303219 252454
rect 360150 252416 360210 252454
rect 239765 252242 239831 252245
rect 282821 252242 282887 252245
rect 239765 252240 240212 252242
rect 239765 252184 239770 252240
rect 239826 252184 240212 252240
rect 239765 252182 240212 252184
rect 279956 252240 282887 252242
rect 279956 252184 282826 252240
rect 282882 252184 282887 252240
rect 279956 252182 282887 252184
rect 239765 252179 239831 252182
rect 282821 252179 282887 252182
rect 323669 252242 323735 252245
rect 326981 252242 327047 252245
rect 323669 252240 327047 252242
rect 323669 252184 323674 252240
rect 323730 252184 326986 252240
rect 327042 252184 327047 252240
rect 323669 252182 327047 252184
rect 323669 252179 323735 252182
rect 326981 252179 327047 252182
rect 282729 251698 282795 251701
rect 279956 251696 282795 251698
rect 279956 251640 282734 251696
rect 282790 251640 282795 251696
rect 279956 251638 282795 251640
rect 282729 251635 282795 251638
rect 300301 251426 300367 251429
rect 300301 251424 360210 251426
rect 300301 251368 300306 251424
rect 300362 251368 360210 251424
rect 300301 251366 360210 251368
rect 300301 251363 300367 251366
rect 360150 251328 360210 251366
rect 230238 251290 230244 251292
rect 110462 251230 230244 251290
rect 110462 251222 110522 251230
rect 230238 251228 230244 251230
rect 230308 251228 230314 251292
rect 109940 251162 110522 251222
rect 237005 251154 237071 251157
rect 282821 251154 282887 251157
rect 237005 251152 240212 251154
rect 237005 251096 237010 251152
rect 237066 251096 240212 251152
rect 237005 251094 240212 251096
rect 279956 251152 282887 251154
rect 279956 251096 282826 251152
rect 282882 251096 282887 251152
rect 279956 251094 282887 251096
rect 237005 251091 237071 251094
rect 282821 251091 282887 251094
rect 357525 250746 357591 250749
rect 357525 250744 360210 250746
rect 357525 250688 357530 250744
rect 357586 250688 360210 250744
rect 357525 250686 360210 250688
rect 357525 250683 357591 250686
rect 282729 250610 282795 250613
rect 279956 250608 282795 250610
rect 279956 250552 282734 250608
rect 282790 250552 282795 250608
rect 279956 250550 282795 250552
rect 282729 250547 282795 250550
rect 360150 250240 360210 250686
rect 502793 250610 502859 250613
rect 499806 250608 502859 250610
rect 499806 250552 502798 250608
rect 502854 250552 502859 250608
rect 499806 250550 502859 250552
rect 236913 250066 236979 250069
rect 282545 250066 282611 250069
rect 236913 250064 240212 250066
rect 236913 250008 236918 250064
rect 236974 250008 240212 250064
rect 236913 250006 240212 250008
rect 279956 250064 282611 250066
rect 279956 250008 282550 250064
rect 282606 250008 282611 250064
rect 279956 250006 282611 250008
rect 236913 250003 236979 250006
rect 282545 250003 282611 250006
rect 499806 249968 499866 250550
rect 502793 250547 502859 250550
rect 224166 249658 224172 249660
rect 110462 249598 224172 249658
rect 110462 249590 110522 249598
rect 224166 249596 224172 249598
rect 224236 249596 224242 249660
rect 109940 249530 110522 249590
rect 288566 249522 288572 249524
rect 279956 249462 288572 249522
rect 288566 249460 288572 249462
rect 288636 249460 288642 249524
rect 298921 249250 298987 249253
rect 298921 249248 360210 249250
rect 298921 249192 298926 249248
rect 298982 249192 360210 249248
rect 298921 249190 360210 249192
rect 298921 249187 298987 249190
rect 360150 249152 360210 249190
rect 282821 248978 282887 248981
rect 279956 248976 282887 248978
rect 279956 248920 282826 248976
rect 282882 248920 282887 248976
rect 279956 248918 282887 248920
rect 282821 248915 282887 248918
rect 282729 248434 282795 248437
rect 279956 248432 282795 248434
rect 279956 248376 282734 248432
rect 282790 248376 282795 248432
rect 279956 248374 282795 248376
rect 282729 248371 282795 248374
rect 286501 248162 286567 248165
rect 286501 248160 360210 248162
rect 286501 248104 286506 248160
rect 286562 248104 360210 248160
rect 286501 248102 360210 248104
rect 286501 248099 286567 248102
rect 360150 248064 360210 248102
rect 218973 248026 219039 248029
rect 110462 248024 219039 248026
rect 110462 247968 218978 248024
rect 219034 247968 219039 248024
rect 110462 247966 219039 247968
rect 110462 247958 110522 247966
rect 218973 247963 219039 247966
rect 109940 247898 110522 247958
rect 282637 247890 282703 247893
rect 279956 247888 282703 247890
rect 279956 247832 282642 247888
rect 282698 247832 282703 247888
rect 279956 247830 282703 247832
rect 282637 247827 282703 247830
rect 288525 247346 288591 247349
rect 279956 247344 288591 247346
rect 279956 247288 288530 247344
rect 288586 247288 288591 247344
rect 279956 247286 288591 247288
rect 288525 247283 288591 247286
rect 357525 246938 357591 246941
rect 360150 246938 360210 246976
rect 357525 246936 360210 246938
rect 357525 246880 357530 246936
rect 357586 246880 360210 246936
rect 357525 246878 360210 246880
rect 357525 246875 357591 246878
rect 238334 246740 238340 246804
rect 238404 246802 238410 246804
rect 282821 246802 282887 246805
rect 238404 246742 240212 246802
rect 279956 246800 282887 246802
rect 279956 246744 282826 246800
rect 282882 246744 282887 246800
rect 279956 246742 282887 246744
rect 238404 246740 238410 246742
rect 282821 246739 282887 246742
rect 218830 246394 218836 246396
rect 110462 246334 218836 246394
rect 110462 246326 110522 246334
rect 218830 246332 218836 246334
rect 218900 246332 218906 246396
rect 109940 246266 110522 246326
rect 289997 246258 290063 246261
rect 279956 246256 290063 246258
rect 279956 246200 290002 246256
rect 290058 246200 290063 246256
rect 279956 246198 290063 246200
rect 289997 246195 290063 246198
rect 301497 245986 301563 245989
rect 301497 245984 360210 245986
rect 301497 245928 301502 245984
rect 301558 245928 360210 245984
rect 301497 245926 360210 245928
rect 301497 245923 301563 245926
rect 360150 245888 360210 245926
rect 197854 245652 197860 245716
rect 197924 245714 197930 245716
rect 287646 245714 287652 245716
rect 197924 245654 240212 245714
rect 279956 245654 287652 245714
rect 197924 245652 197930 245654
rect 287646 245652 287652 245654
rect 287716 245652 287722 245716
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 290590 245170 290596 245172
rect 279956 245110 290596 245170
rect 290590 245108 290596 245110
rect 290660 245108 290666 245172
rect 357525 245170 357591 245173
rect 357525 245168 360210 245170
rect 357525 245112 357530 245168
rect 357586 245112 360210 245168
rect 357525 245110 360210 245112
rect 357525 245107 357591 245110
rect 360150 244800 360210 245110
rect 231158 244762 231164 244764
rect 110462 244702 231164 244762
rect 110462 244694 110522 244702
rect 231158 244700 231164 244702
rect 231228 244700 231234 244764
rect 109940 244634 110522 244694
rect 175917 244626 175983 244629
rect 283281 244626 283347 244629
rect 175917 244624 240212 244626
rect 175917 244568 175922 244624
rect 175978 244568 240212 244624
rect 175917 244566 240212 244568
rect 279956 244624 283347 244626
rect 279956 244568 283286 244624
rect 283342 244568 283347 244624
rect 279956 244566 283347 244568
rect 175917 244563 175983 244566
rect 283281 244563 283347 244566
rect 503805 244354 503871 244357
rect 503670 244352 503871 244354
rect 503670 244296 503810 244352
rect 503866 244296 503871 244352
rect 503670 244294 503871 244296
rect 503670 244218 503730 244294
rect 503805 244291 503871 244294
rect 499806 244158 503730 244218
rect 285990 244082 285996 244084
rect 279956 244022 285996 244082
rect 285990 244020 285996 244022
rect 286060 244020 286066 244084
rect 499806 243984 499866 244158
rect 357525 243946 357591 243949
rect 357525 243944 360210 243946
rect 357525 243888 357530 243944
rect 357586 243888 360210 243944
rect 357525 243886 360210 243888
rect 357525 243883 357591 243886
rect 360150 243712 360210 243886
rect 220353 243538 220419 243541
rect 280286 243538 280292 243540
rect 220353 243536 240212 243538
rect 220353 243480 220358 243536
rect 220414 243480 240212 243536
rect 220353 243478 240212 243480
rect 279956 243478 280292 243538
rect 220353 243475 220419 243478
rect 280286 243476 280292 243478
rect 280356 243476 280362 243540
rect 221222 243130 221228 243132
rect 110462 243070 221228 243130
rect 110462 243062 110522 243070
rect 221222 243068 221228 243070
rect 221292 243068 221298 243132
rect 109940 243002 110522 243062
rect 284753 242994 284819 242997
rect 279956 242992 284819 242994
rect 279956 242936 284758 242992
rect 284814 242936 284819 242992
rect 279956 242934 284819 242936
rect 284753 242931 284819 242934
rect 115197 242858 115263 242861
rect 116577 242858 116643 242861
rect 115197 242856 116643 242858
rect 115197 242800 115202 242856
rect 115258 242800 116582 242856
rect 116638 242800 116643 242856
rect 115197 242798 116643 242800
rect 115197 242795 115263 242798
rect 116577 242795 116643 242798
rect 318149 242722 318215 242725
rect 318149 242720 360210 242722
rect 318149 242664 318154 242720
rect 318210 242664 360210 242720
rect 318149 242662 360210 242664
rect 318149 242659 318215 242662
rect 360150 242624 360210 242662
rect 210550 242388 210556 242452
rect 210620 242450 210626 242452
rect 287053 242450 287119 242453
rect 210620 242390 240212 242450
rect 279956 242448 287119 242450
rect 279956 242392 287058 242448
rect 287114 242392 287119 242448
rect 279956 242390 287119 242392
rect 210620 242388 210626 242390
rect 287053 242387 287119 242390
rect 290774 241906 290780 241908
rect 279956 241846 290780 241906
rect 290774 241844 290780 241846
rect 290844 241844 290850 241908
rect 295977 241634 296043 241637
rect 295977 241632 360210 241634
rect 295977 241576 295982 241632
rect 296038 241576 360210 241632
rect 295977 241574 360210 241576
rect 295977 241571 296043 241574
rect 360150 241536 360210 241574
rect 218646 241498 218652 241500
rect 110462 241438 218652 241498
rect 110462 241430 110522 241438
rect 218646 241436 218652 241438
rect 218716 241436 218722 241500
rect 109940 241370 110522 241430
rect 233877 241362 233943 241365
rect 299422 241362 299428 241364
rect 233877 241360 240212 241362
rect 233877 241304 233882 241360
rect 233938 241304 240212 241360
rect 233877 241302 240212 241304
rect 279956 241302 299428 241362
rect 233877 241299 233943 241302
rect 299422 241300 299428 241302
rect 299492 241300 299498 241364
rect -960 241090 480 241180
rect 3550 241090 3556 241092
rect -960 241030 3556 241090
rect -960 240940 480 241030
rect 3550 241028 3556 241030
rect 3620 241028 3626 241092
rect 299606 240818 299612 240820
rect 279956 240758 299612 240818
rect 299606 240756 299612 240758
rect 299676 240756 299682 240820
rect 290457 240546 290523 240549
rect 290457 240544 360210 240546
rect 290457 240488 290462 240544
rect 290518 240488 360210 240544
rect 290457 240486 360210 240488
rect 290457 240483 290523 240486
rect 360150 240448 360210 240486
rect 227161 240274 227227 240277
rect 291326 240274 291332 240276
rect 227161 240272 240212 240274
rect 227161 240216 227166 240272
rect 227222 240216 240212 240272
rect 227161 240214 240212 240216
rect 279956 240214 291332 240274
rect 227161 240211 227227 240214
rect 291326 240212 291332 240214
rect 291396 240212 291402 240276
rect 77431 240138 77497 240141
rect 88701 240138 88767 240141
rect 77431 240136 88767 240138
rect 77431 240080 77436 240136
rect 77492 240080 88706 240136
rect 88762 240080 88767 240136
rect 77431 240078 88767 240080
rect 77431 240075 77497 240078
rect 88701 240075 88767 240078
rect 90679 240138 90745 240141
rect 93301 240138 93367 240141
rect 90679 240136 93367 240138
rect 90679 240080 90684 240136
rect 90740 240080 93306 240136
rect 93362 240080 93367 240136
rect 90679 240078 93367 240080
rect 90679 240075 90745 240078
rect 93301 240075 93367 240078
rect 93485 240138 93551 240141
rect 212073 240138 212139 240141
rect 93485 240136 212139 240138
rect 93485 240080 93490 240136
rect 93546 240080 212078 240136
rect 212134 240080 212139 240136
rect 93485 240078 212139 240080
rect 93485 240075 93551 240078
rect 212073 240075 212139 240078
rect 79409 240002 79475 240005
rect 212257 240002 212323 240005
rect 79409 240000 212323 240002
rect 79409 239944 79414 240000
rect 79470 239944 212262 240000
rect 212318 239944 212323 240000
rect 79409 239942 212323 239944
rect 79409 239939 79475 239942
rect 212257 239939 212323 239942
rect 92335 239866 92401 239869
rect 93301 239866 93367 239869
rect 217777 239866 217843 239869
rect 92335 239864 93226 239866
rect 92335 239808 92340 239864
rect 92396 239808 93226 239864
rect 92335 239806 93226 239808
rect 92335 239803 92401 239806
rect 93166 239730 93226 239806
rect 93301 239864 217843 239866
rect 93301 239808 93306 239864
rect 93362 239808 217782 239864
rect 217838 239808 217843 239864
rect 93301 239806 217843 239808
rect 93301 239803 93367 239806
rect 217777 239803 217843 239806
rect 217593 239730 217659 239733
rect 288382 239730 288388 239732
rect 93166 239728 217659 239730
rect 93166 239672 217598 239728
rect 217654 239672 217659 239728
rect 93166 239670 217659 239672
rect 279956 239670 288388 239730
rect 217593 239667 217659 239670
rect 288382 239668 288388 239670
rect 288452 239668 288458 239732
rect 357525 239730 357591 239733
rect 357525 239728 360210 239730
rect 357525 239672 357530 239728
rect 357586 239672 360210 239728
rect 357525 239670 360210 239672
rect 357525 239667 357591 239670
rect 88701 239594 88767 239597
rect 93485 239594 93551 239597
rect 88701 239592 93551 239594
rect 88701 239536 88706 239592
rect 88762 239536 93490 239592
rect 93546 239536 93551 239592
rect 88701 239534 93551 239536
rect 88701 239531 88767 239534
rect 93485 239531 93551 239534
rect 95969 239594 96035 239597
rect 214649 239594 214715 239597
rect 95969 239592 214715 239594
rect 95969 239536 95974 239592
rect 96030 239536 214654 239592
rect 214710 239536 214715 239592
rect 95969 239534 214715 239536
rect 95969 239531 96035 239534
rect 214649 239531 214715 239534
rect 94313 239458 94379 239461
rect 209037 239458 209103 239461
rect 94313 239456 209103 239458
rect 94313 239400 94318 239456
rect 94374 239400 209042 239456
rect 209098 239400 209103 239456
rect 94313 239398 209103 239400
rect 94313 239395 94379 239398
rect 209037 239395 209103 239398
rect 360150 239360 360210 239670
rect 107561 239322 107627 239325
rect 212441 239322 212507 239325
rect 107561 239320 212507 239322
rect 107561 239264 107566 239320
rect 107622 239264 212446 239320
rect 212502 239264 212507 239320
rect 107561 239262 212507 239264
rect 107561 239259 107627 239262
rect 212441 239259 212507 239262
rect 237782 239124 237788 239188
rect 237852 239186 237858 239188
rect 295558 239186 295564 239188
rect 237852 239126 240212 239186
rect 279956 239126 295564 239186
rect 237852 239124 237858 239126
rect 295558 239124 295564 239126
rect 295628 239124 295634 239188
rect 97625 238642 97691 238645
rect 215109 238642 215175 238645
rect 296662 238642 296668 238644
rect 97625 238640 215175 238642
rect 97625 238584 97630 238640
rect 97686 238584 215114 238640
rect 215170 238584 215175 238640
rect 97625 238582 215175 238584
rect 279956 238582 296668 238642
rect 97625 238579 97691 238582
rect 215109 238579 215175 238582
rect 296662 238580 296668 238582
rect 296732 238580 296738 238644
rect 66161 238506 66227 238509
rect 98637 238506 98703 238509
rect 66161 238504 98703 238506
rect 66161 238448 66166 238504
rect 66222 238448 98642 238504
rect 98698 238448 98703 238504
rect 66161 238446 98703 238448
rect 66161 238443 66227 238446
rect 98637 238443 98703 238446
rect 100661 238506 100727 238509
rect 108389 238506 108455 238509
rect 214281 238506 214347 238509
rect 100661 238504 108314 238506
rect 100661 238448 100666 238504
rect 100722 238448 108314 238504
rect 100661 238446 108314 238448
rect 100661 238443 100727 238446
rect 56225 238370 56291 238373
rect 88241 238370 88307 238373
rect 56225 238368 88307 238370
rect 56225 238312 56230 238368
rect 56286 238312 88246 238368
rect 88302 238312 88307 238368
rect 56225 238310 88307 238312
rect 56225 238307 56291 238310
rect 88241 238307 88307 238310
rect 99189 238370 99255 238373
rect 108113 238370 108179 238373
rect 99189 238368 108179 238370
rect 99189 238312 99194 238368
rect 99250 238312 108118 238368
rect 108174 238312 108179 238368
rect 99189 238310 108179 238312
rect 108254 238370 108314 238446
rect 108389 238504 214347 238506
rect 108389 238448 108394 238504
rect 108450 238448 214286 238504
rect 214342 238448 214347 238504
rect 108389 238446 214347 238448
rect 108389 238443 108455 238446
rect 214281 238443 214347 238446
rect 214925 238370 214991 238373
rect 108254 238368 214991 238370
rect 108254 238312 214930 238368
rect 214986 238312 214991 238368
rect 108254 238310 214991 238312
rect 99189 238307 99255 238310
rect 108113 238307 108179 238310
rect 214925 238307 214991 238310
rect 294689 238370 294755 238373
rect 502701 238370 502767 238373
rect 294689 238368 360210 238370
rect 294689 238312 294694 238368
rect 294750 238312 360210 238368
rect 294689 238310 360210 238312
rect 294689 238307 294755 238310
rect 360150 238272 360210 238310
rect 499806 238368 502767 238370
rect 499806 238312 502706 238368
rect 502762 238312 502767 238368
rect 499806 238310 502767 238312
rect 59261 238234 59327 238237
rect 88977 238234 89043 238237
rect 59261 238232 89043 238234
rect 59261 238176 59266 238232
rect 59322 238176 88982 238232
rect 89038 238176 89043 238232
rect 59261 238174 89043 238176
rect 59261 238171 59327 238174
rect 88977 238171 89043 238174
rect 102593 238234 102659 238237
rect 214741 238234 214807 238237
rect 102593 238232 214807 238234
rect 102593 238176 102598 238232
rect 102654 238176 214746 238232
rect 214802 238176 214807 238232
rect 102593 238174 214807 238176
rect 102593 238171 102659 238174
rect 214741 238171 214807 238174
rect 52913 238098 52979 238101
rect 81433 238098 81499 238101
rect 52913 238096 81499 238098
rect 52913 238040 52918 238096
rect 52974 238040 81438 238096
rect 81494 238040 81499 238096
rect 52913 238038 81499 238040
rect 52913 238035 52979 238038
rect 81433 238035 81499 238038
rect 82721 238098 82787 238101
rect 102133 238098 102199 238101
rect 82721 238096 102199 238098
rect 82721 238040 82726 238096
rect 82782 238040 102138 238096
rect 102194 238040 102199 238096
rect 82721 238038 102199 238040
rect 82721 238035 82787 238038
rect 102133 238035 102199 238038
rect 104249 238098 104315 238101
rect 214557 238098 214623 238101
rect 104249 238096 214623 238098
rect 104249 238040 104254 238096
rect 104310 238040 214562 238096
rect 214618 238040 214623 238096
rect 104249 238038 214623 238040
rect 104249 238035 104315 238038
rect 214557 238035 214623 238038
rect 237598 238036 237604 238100
rect 237668 238098 237674 238100
rect 296846 238098 296852 238100
rect 237668 238038 240212 238098
rect 279956 238038 296852 238098
rect 237668 238036 237674 238038
rect 296846 238036 296852 238038
rect 296916 238036 296922 238100
rect 499806 238000 499866 238310
rect 502701 238307 502767 238310
rect 57789 237962 57855 237965
rect 86861 237962 86927 237965
rect 57789 237960 86927 237962
rect 57789 237904 57794 237960
rect 57850 237904 86866 237960
rect 86922 237904 86927 237960
rect 57789 237902 86927 237904
rect 57789 237899 57855 237902
rect 86861 237899 86927 237902
rect 87689 237962 87755 237965
rect 104801 237962 104867 237965
rect 87689 237960 104867 237962
rect 87689 237904 87694 237960
rect 87750 237904 104806 237960
rect 104862 237904 104867 237960
rect 87689 237902 104867 237904
rect 87689 237899 87755 237902
rect 104801 237899 104867 237902
rect 105905 237962 105971 237965
rect 212349 237962 212415 237965
rect 105905 237960 212415 237962
rect 105905 237904 105910 237960
rect 105966 237904 212354 237960
rect 212410 237904 212415 237960
rect 105905 237902 212415 237904
rect 105905 237899 105971 237902
rect 212349 237899 212415 237902
rect 74441 237826 74507 237829
rect 99373 237826 99439 237829
rect 74441 237824 99439 237826
rect 74441 237768 74446 237824
rect 74502 237768 99378 237824
rect 99434 237768 99439 237824
rect 74441 237766 99439 237768
rect 74441 237763 74507 237766
rect 99373 237763 99439 237766
rect 108849 237826 108915 237829
rect 212165 237826 212231 237829
rect 108849 237824 212231 237826
rect 108849 237768 108854 237824
rect 108910 237768 212170 237824
rect 212226 237768 212231 237824
rect 108849 237766 212231 237768
rect 108849 237763 108915 237766
rect 212165 237763 212231 237766
rect 86033 237690 86099 237693
rect 106181 237690 106247 237693
rect 86033 237688 106247 237690
rect 86033 237632 86038 237688
rect 86094 237632 106186 237688
rect 106242 237632 106247 237688
rect 86033 237630 106247 237632
rect 86033 237627 86099 237630
rect 106181 237627 106247 237630
rect 89345 237554 89411 237557
rect 108297 237554 108363 237557
rect 282821 237554 282887 237557
rect 89345 237552 108363 237554
rect 89345 237496 89350 237552
rect 89406 237496 108302 237552
rect 108358 237496 108363 237552
rect 89345 237494 108363 237496
rect 279956 237552 282887 237554
rect 279956 237496 282826 237552
rect 282882 237496 282887 237552
rect 279956 237494 282887 237496
rect 89345 237491 89411 237494
rect 108297 237491 108363 237494
rect 282821 237491 282887 237494
rect 49325 237418 49391 237421
rect 53097 237418 53163 237421
rect 49325 237416 53163 237418
rect 49325 237360 49330 237416
rect 49386 237360 53102 237416
rect 53158 237360 53163 237416
rect 49325 237358 53163 237360
rect 49325 237355 49391 237358
rect 53097 237355 53163 237358
rect 61193 237418 61259 237421
rect 97901 237418 97967 237421
rect 61193 237416 97967 237418
rect 61193 237360 61198 237416
rect 61254 237360 97906 237416
rect 97962 237360 97967 237416
rect 61193 237358 97967 237360
rect 61193 237355 61259 237358
rect 97901 237355 97967 237358
rect 69473 237282 69539 237285
rect 223021 237282 223087 237285
rect 69473 237280 223087 237282
rect 69473 237224 69478 237280
rect 69534 237224 223026 237280
rect 223082 237224 223087 237280
rect 69473 237222 223087 237224
rect 69473 237219 69539 237222
rect 223021 237219 223087 237222
rect 307017 237282 307083 237285
rect 307017 237280 360210 237282
rect 307017 237224 307022 237280
rect 307078 237224 360210 237280
rect 307017 237222 360210 237224
rect 307017 237219 307083 237222
rect 360150 237184 360210 237222
rect 71129 237146 71195 237149
rect 222837 237146 222903 237149
rect 71129 237144 222903 237146
rect 71129 237088 71134 237144
rect 71190 237088 222842 237144
rect 222898 237088 222903 237144
rect 71129 237086 222903 237088
rect 71129 237083 71195 237086
rect 222837 237083 222903 237086
rect 62849 237010 62915 237013
rect 213177 237010 213243 237013
rect 62849 237008 213243 237010
rect 62849 236952 62854 237008
rect 62910 236952 213182 237008
rect 213238 236952 213243 237008
rect 62849 236950 213243 236952
rect 62849 236947 62915 236950
rect 213177 236947 213243 236950
rect 238150 236948 238156 237012
rect 238220 237010 238226 237012
rect 283557 237010 283623 237013
rect 238220 236950 240212 237010
rect 279956 237008 283623 237010
rect 279956 236952 283562 237008
rect 283618 236952 283623 237008
rect 279956 236950 283623 236952
rect 238220 236948 238226 236950
rect 283557 236947 283623 236950
rect 72785 236874 72851 236877
rect 220261 236874 220327 236877
rect 72785 236872 220327 236874
rect 72785 236816 72790 236872
rect 72846 236816 220266 236872
rect 220322 236816 220327 236872
rect 72785 236814 220327 236816
rect 72785 236811 72851 236814
rect 220261 236811 220327 236814
rect 81065 236738 81131 236741
rect 220077 236738 220143 236741
rect 81065 236736 220143 236738
rect 81065 236680 81070 236736
rect 81126 236680 220082 236736
rect 220138 236680 220143 236736
rect 81065 236678 220143 236680
rect 81065 236675 81131 236678
rect 220077 236675 220143 236678
rect 84101 236602 84167 236605
rect 211797 236602 211863 236605
rect 84101 236600 211863 236602
rect 84101 236544 84106 236600
rect 84162 236544 211802 236600
rect 211858 236544 211863 236600
rect 84101 236542 211863 236544
rect 84101 236539 84167 236542
rect 211797 236539 211863 236542
rect 284661 236466 284727 236469
rect 279956 236464 284727 236466
rect 279956 236408 284666 236464
rect 284722 236408 284727 236464
rect 279956 236406 284727 236408
rect 284661 236403 284727 236406
rect 289169 236194 289235 236197
rect 289169 236192 360210 236194
rect 289169 236136 289174 236192
rect 289230 236136 360210 236192
rect 289169 236134 360210 236136
rect 289169 236131 289235 236134
rect 360150 236096 360210 236134
rect 237373 236058 237439 236061
rect 237966 236058 237972 236060
rect 237373 236056 237972 236058
rect 237373 236000 237378 236056
rect 237434 236000 237972 236056
rect 237373 235998 237972 236000
rect 237373 235995 237439 235998
rect 237966 235996 237972 235998
rect 238036 235996 238042 236060
rect 59118 235860 59124 235924
rect 59188 235922 59194 235924
rect 281533 235922 281599 235925
rect 59188 235862 240212 235922
rect 279956 235920 281599 235922
rect 279956 235864 281538 235920
rect 281594 235864 281599 235920
rect 279956 235862 281599 235864
rect 59188 235860 59194 235862
rect 281533 235859 281599 235862
rect 64505 235786 64571 235789
rect 218789 235786 218855 235789
rect 64505 235784 218855 235786
rect 64505 235728 64510 235784
rect 64566 235728 218794 235784
rect 218850 235728 218855 235784
rect 64505 235726 218855 235728
rect 64505 235723 64571 235726
rect 218789 235723 218855 235726
rect 75821 235650 75887 235653
rect 211889 235650 211955 235653
rect 75821 235648 211955 235650
rect 75821 235592 75826 235648
rect 75882 235592 211894 235648
rect 211950 235592 211955 235648
rect 75821 235590 211955 235592
rect 75821 235587 75887 235590
rect 211889 235587 211955 235590
rect 357525 235514 357591 235517
rect 357525 235512 360210 235514
rect 357525 235456 357530 235512
rect 357586 235456 360210 235512
rect 357525 235454 360210 235456
rect 357525 235451 357591 235454
rect 56501 235378 56567 235381
rect 221457 235378 221523 235381
rect 291510 235378 291516 235380
rect 56501 235376 221523 235378
rect 56501 235320 56506 235376
rect 56562 235320 221462 235376
rect 221518 235320 221523 235376
rect 56501 235318 221523 235320
rect 279956 235318 291516 235378
rect 56501 235315 56567 235318
rect 221457 235315 221523 235318
rect 291510 235316 291516 235318
rect 291580 235316 291586 235380
rect 60406 235180 60412 235244
rect 60476 235242 60482 235244
rect 238334 235242 238340 235244
rect 60476 235182 238340 235242
rect 60476 235180 60482 235182
rect 238334 235180 238340 235182
rect 238404 235180 238410 235244
rect 360150 235008 360210 235454
rect 237966 234772 237972 234836
rect 238036 234834 238042 234836
rect 303654 234834 303660 234836
rect 238036 234774 240212 234834
rect 279956 234774 303660 234834
rect 238036 234772 238042 234774
rect 303654 234772 303660 234774
rect 303724 234772 303730 234836
rect 54569 234562 54635 234565
rect 221549 234562 221615 234565
rect 54569 234560 221615 234562
rect 54569 234504 54574 234560
rect 54630 234504 221554 234560
rect 221610 234504 221615 234560
rect 54569 234502 221615 234504
rect 54569 234499 54635 234502
rect 221549 234499 221615 234502
rect 295374 234290 295380 234292
rect 279956 234230 295380 234290
rect 295374 234228 295380 234230
rect 295444 234228 295450 234292
rect 293217 234018 293283 234021
rect 293217 234016 360210 234018
rect 293217 233960 293222 234016
rect 293278 233960 360210 234016
rect 293217 233958 360210 233960
rect 293217 233955 293283 233958
rect 360150 233920 360210 233958
rect 58566 233684 58572 233748
rect 58636 233746 58642 233748
rect 280286 233746 280292 233748
rect 58636 233686 240212 233746
rect 279956 233686 280292 233746
rect 58636 233684 58642 233686
rect 280286 233684 280292 233686
rect 280356 233684 280362 233748
rect 301814 233202 301820 233204
rect 279956 233142 301820 233202
rect 301814 233140 301820 233142
rect 301884 233140 301890 233204
rect 291929 232930 291995 232933
rect 502517 232930 502583 232933
rect 291929 232928 360210 232930
rect 291929 232872 291934 232928
rect 291990 232872 360210 232928
rect 291929 232870 360210 232872
rect 291929 232867 291995 232870
rect 360150 232832 360210 232870
rect 499806 232928 502583 232930
rect 499806 232872 502522 232928
rect 502578 232872 502583 232928
rect 499806 232870 502583 232872
rect 59261 232658 59327 232661
rect 306373 232658 306439 232661
rect 59261 232656 240212 232658
rect 59261 232600 59266 232656
rect 59322 232600 240212 232656
rect 59261 232598 240212 232600
rect 279956 232656 306439 232658
rect 279956 232600 306378 232656
rect 306434 232600 306439 232656
rect 279956 232598 306439 232600
rect 59261 232595 59327 232598
rect 306373 232595 306439 232598
rect 303838 232114 303844 232116
rect 279956 232054 303844 232114
rect 303838 232052 303844 232054
rect 303908 232052 303914 232116
rect 499806 232016 499866 232870
rect 502517 232867 502583 232870
rect 580349 232386 580415 232389
rect 583520 232386 584960 232476
rect 580349 232384 584960 232386
rect 580349 232328 580354 232384
rect 580410 232328 584960 232384
rect 580349 232326 584960 232328
rect 580349 232323 580415 232326
rect 583520 232236 584960 232326
rect 300209 231842 300275 231845
rect 300209 231840 360210 231842
rect 300209 231784 300214 231840
rect 300270 231784 360210 231840
rect 300209 231782 360210 231784
rect 300209 231779 300275 231782
rect 360150 231744 360210 231782
rect 237414 231508 237420 231572
rect 237484 231570 237490 231572
rect 285806 231570 285812 231572
rect 237484 231510 240212 231570
rect 279956 231510 285812 231570
rect 237484 231508 237490 231510
rect 285806 231508 285812 231510
rect 285876 231508 285882 231572
rect 357525 231298 357591 231301
rect 357525 231296 360210 231298
rect 357525 231240 357530 231296
rect 357586 231240 360210 231296
rect 357525 231238 360210 231240
rect 357525 231235 357591 231238
rect 60038 231100 60044 231164
rect 60108 231162 60114 231164
rect 237598 231162 237604 231164
rect 60108 231102 237604 231162
rect 60108 231100 60114 231102
rect 237598 231100 237604 231102
rect 237668 231100 237674 231164
rect 294638 231026 294644 231028
rect 279956 230966 294644 231026
rect 294638 230964 294644 230966
rect 294708 230964 294714 231028
rect 360150 230656 360210 231238
rect 58617 230482 58683 230485
rect 306414 230482 306420 230484
rect 58617 230480 240212 230482
rect 58617 230424 58622 230480
rect 58678 230424 240212 230480
rect 58617 230422 240212 230424
rect 279956 230422 306420 230482
rect 58617 230419 58683 230422
rect 306414 230420 306420 230422
rect 306484 230420 306490 230484
rect 322289 230482 322355 230485
rect 323669 230482 323735 230485
rect 322289 230480 323735 230482
rect 322289 230424 322294 230480
rect 322350 230424 323674 230480
rect 323730 230424 323735 230480
rect 322289 230422 323735 230424
rect 322289 230419 322355 230422
rect 323669 230419 323735 230422
rect 286225 229938 286291 229941
rect 279956 229936 286291 229938
rect 279956 229880 286230 229936
rect 286286 229880 286291 229936
rect 279956 229878 286291 229880
rect 286225 229875 286291 229878
rect 286317 229666 286383 229669
rect 286317 229664 360210 229666
rect 286317 229608 286322 229664
rect 286378 229608 360210 229664
rect 286317 229606 360210 229608
rect 286317 229603 286383 229606
rect 360150 229568 360210 229606
rect 238201 229394 238267 229397
rect 280245 229394 280311 229397
rect 238201 229392 240212 229394
rect 238201 229336 238206 229392
rect 238262 229336 240212 229392
rect 238201 229334 240212 229336
rect 279956 229392 280311 229394
rect 279956 229336 280250 229392
rect 280306 229336 280311 229392
rect 279956 229334 280311 229336
rect 238201 229331 238267 229334
rect 280245 229331 280311 229334
rect 282545 228850 282611 228853
rect 279956 228848 282611 228850
rect 279956 228792 282550 228848
rect 282606 228792 282611 228848
rect 279956 228790 282611 228792
rect 282545 228787 282611 228790
rect 302969 228578 303035 228581
rect 302969 228576 360210 228578
rect 302969 228520 302974 228576
rect 303030 228520 360210 228576
rect 302969 228518 360210 228520
rect 302969 228515 303035 228518
rect 360150 228480 360210 228518
rect 3366 228244 3372 228308
rect 3436 228306 3442 228308
rect 214782 228306 214788 228308
rect 3436 228246 214788 228306
rect 3436 228244 3442 228246
rect 214782 228244 214788 228246
rect 214852 228244 214858 228308
rect 238109 228306 238175 228309
rect 281533 228306 281599 228309
rect 238109 228304 240212 228306
rect 238109 228248 238114 228304
rect 238170 228248 240212 228304
rect 238109 228246 240212 228248
rect 279956 228304 281599 228306
rect 279956 228248 281538 228304
rect 281594 228248 281599 228304
rect 279956 228246 281599 228248
rect 238109 228243 238175 228246
rect 281533 228243 281599 228246
rect -960 227884 480 228124
rect 285029 227762 285095 227765
rect 279956 227760 285095 227762
rect 279956 227704 285034 227760
rect 285090 227704 285095 227760
rect 279956 227702 285095 227704
rect 285029 227699 285095 227702
rect 298737 227490 298803 227493
rect 298737 227488 360210 227490
rect 298737 227432 298742 227488
rect 298798 227432 360210 227488
rect 298737 227430 360210 227432
rect 298737 227427 298803 227430
rect 360150 227392 360210 227430
rect 238017 227218 238083 227221
rect 281625 227218 281691 227221
rect 238017 227216 240212 227218
rect 238017 227160 238022 227216
rect 238078 227160 240212 227216
rect 238017 227158 240212 227160
rect 279956 227216 281691 227218
rect 279956 227160 281630 227216
rect 281686 227160 281691 227216
rect 279956 227158 281691 227160
rect 238017 227155 238083 227158
rect 281625 227155 281691 227158
rect 58934 226884 58940 226948
rect 59004 226946 59010 226948
rect 237414 226946 237420 226948
rect 59004 226886 237420 226946
rect 59004 226884 59010 226886
rect 237414 226884 237420 226886
rect 237484 226884 237490 226948
rect 281993 226674 282059 226677
rect 279956 226672 282059 226674
rect 279956 226616 281998 226672
rect 282054 226616 282059 226672
rect 279956 226614 282059 226616
rect 281993 226611 282059 226614
rect 238569 226404 238635 226405
rect 238518 226402 238524 226404
rect 238478 226342 238524 226402
rect 238588 226400 238635 226404
rect 238630 226344 238635 226400
rect 238518 226340 238524 226342
rect 238588 226340 238635 226344
rect 238569 226339 238635 226340
rect 357525 226266 357591 226269
rect 360150 226266 360210 226304
rect 502609 226266 502675 226269
rect 357525 226264 360210 226266
rect 357525 226208 357530 226264
rect 357586 226208 360210 226264
rect 357525 226206 360210 226208
rect 499806 226264 502675 226266
rect 499806 226208 502614 226264
rect 502670 226208 502675 226264
rect 499806 226206 502675 226208
rect 357525 226203 357591 226206
rect 238293 226130 238359 226133
rect 280337 226130 280403 226133
rect 238293 226128 240212 226130
rect 238293 226072 238298 226128
rect 238354 226072 240212 226128
rect 238293 226070 240212 226072
rect 279956 226128 280403 226130
rect 279956 226072 280342 226128
rect 280398 226072 280403 226128
rect 279956 226070 280403 226072
rect 238293 226067 238359 226070
rect 280337 226067 280403 226070
rect 499806 226032 499866 226206
rect 502609 226203 502675 226206
rect 357709 225722 357775 225725
rect 357709 225720 360210 225722
rect 357709 225664 357714 225720
rect 357770 225664 360210 225720
rect 357709 225662 360210 225664
rect 357709 225659 357775 225662
rect 60222 225524 60228 225588
rect 60292 225586 60298 225588
rect 237782 225586 237788 225588
rect 60292 225526 237788 225586
rect 60292 225524 60298 225526
rect 237782 225524 237788 225526
rect 237852 225524 237858 225588
rect 285673 225586 285739 225589
rect 279956 225584 285739 225586
rect 279956 225528 285678 225584
rect 285734 225528 285739 225584
rect 279956 225526 285739 225528
rect 285673 225523 285739 225526
rect 360150 225216 360210 225662
rect 116577 225042 116643 225045
rect 118049 225042 118115 225045
rect 116577 225040 118115 225042
rect 116577 224984 116582 225040
rect 116638 224984 118054 225040
rect 118110 224984 118115 225040
rect 116577 224982 118115 224984
rect 116577 224979 116643 224982
rect 118049 224979 118115 224982
rect 216121 225042 216187 225045
rect 285949 225042 286015 225045
rect 216121 225040 240212 225042
rect 216121 224984 216126 225040
rect 216182 224984 240212 225040
rect 216121 224982 240212 224984
rect 279956 225040 286015 225042
rect 279956 224984 285954 225040
rect 286010 224984 286015 225040
rect 279956 224982 286015 224984
rect 216121 224979 216187 224982
rect 285949 224979 286015 224982
rect 282085 224498 282151 224501
rect 279956 224496 282151 224498
rect 279956 224440 282090 224496
rect 282146 224440 282151 224496
rect 279956 224438 282151 224440
rect 282085 224435 282151 224438
rect 357525 224498 357591 224501
rect 357525 224496 360210 224498
rect 357525 224440 357530 224496
rect 357586 224440 360210 224496
rect 357525 224438 360210 224440
rect 357525 224435 357591 224438
rect 360150 224128 360210 224438
rect 61377 223954 61443 223957
rect 286133 223954 286199 223957
rect 61377 223952 240212 223954
rect 61377 223896 61382 223952
rect 61438 223896 240212 223952
rect 61377 223894 240212 223896
rect 279956 223952 286199 223954
rect 279956 223896 286138 223952
rect 286194 223896 286199 223952
rect 279956 223894 286199 223896
rect 61377 223891 61443 223894
rect 286133 223891 286199 223894
rect 280153 223410 280219 223413
rect 279956 223408 280219 223410
rect 279956 223352 280158 223408
rect 280214 223352 280219 223408
rect 279956 223350 280219 223352
rect 280153 223347 280219 223350
rect 357525 223274 357591 223277
rect 357525 223272 360210 223274
rect 357525 223216 357530 223272
rect 357586 223216 360210 223272
rect 357525 223214 360210 223216
rect 357525 223211 357591 223214
rect 360150 223040 360210 223214
rect 61469 222866 61535 222869
rect 286041 222866 286107 222869
rect 61469 222864 240212 222866
rect 61469 222808 61474 222864
rect 61530 222808 240212 222864
rect 61469 222806 240212 222808
rect 279956 222864 286107 222866
rect 279956 222808 286046 222864
rect 286102 222808 286107 222864
rect 279956 222806 286107 222808
rect 61469 222803 61535 222806
rect 286041 222803 286107 222806
rect 118049 222322 118115 222325
rect 280521 222322 280587 222325
rect 118049 222320 120090 222322
rect 118049 222264 118054 222320
rect 118110 222264 120090 222320
rect 118049 222262 120090 222264
rect 279956 222320 280587 222322
rect 279956 222264 280526 222320
rect 280582 222264 280587 222320
rect 279956 222262 280587 222264
rect 118049 222259 118115 222262
rect 120030 222186 120090 222262
rect 280521 222259 280587 222262
rect 122097 222186 122163 222189
rect 120030 222184 122163 222186
rect 120030 222128 122102 222184
rect 122158 222128 122163 222184
rect 120030 222126 122163 222128
rect 122097 222123 122163 222126
rect 357525 222050 357591 222053
rect 357525 222048 360210 222050
rect 357525 221992 357530 222048
rect 357586 221992 360210 222048
rect 357525 221990 360210 221992
rect 357525 221987 357591 221990
rect 360150 221952 360210 221990
rect 60273 221778 60339 221781
rect 280613 221778 280679 221781
rect 60273 221776 240212 221778
rect 60273 221720 60278 221776
rect 60334 221720 240212 221776
rect 60273 221718 240212 221720
rect 279956 221776 280679 221778
rect 279956 221720 280618 221776
rect 280674 221720 280679 221776
rect 279956 221718 280679 221720
rect 60273 221715 60339 221718
rect 280613 221715 280679 221718
rect 357709 221506 357775 221509
rect 357709 221504 360210 221506
rect 357709 221448 357714 221504
rect 357770 221448 360210 221504
rect 357709 221446 360210 221448
rect 357709 221443 357775 221446
rect 285121 221234 285187 221237
rect 279956 221232 285187 221234
rect 279956 221176 285126 221232
rect 285182 221176 285187 221232
rect 279956 221174 285187 221176
rect 285121 221171 285187 221174
rect 360150 220864 360210 221446
rect 502425 220826 502491 220829
rect 499806 220824 502491 220826
rect 499806 220768 502430 220824
rect 502486 220768 502491 220824
rect 499806 220766 502491 220768
rect 59905 220690 59971 220693
rect 280429 220690 280495 220693
rect 59905 220688 240212 220690
rect 59905 220632 59910 220688
rect 59966 220632 240212 220688
rect 59905 220630 240212 220632
rect 279956 220688 280495 220690
rect 279956 220632 280434 220688
rect 280490 220632 280495 220688
rect 279956 220630 280495 220632
rect 59905 220627 59971 220630
rect 280429 220627 280495 220630
rect 59997 220146 60063 220149
rect 284753 220146 284819 220149
rect 59997 220144 219450 220146
rect 59997 220088 60002 220144
rect 60058 220088 219450 220144
rect 59997 220086 219450 220088
rect 279956 220144 284819 220146
rect 279956 220088 284758 220144
rect 284814 220088 284819 220144
rect 279956 220086 284819 220088
rect 59997 220083 60063 220086
rect 219390 219602 219450 220086
rect 284753 220083 284819 220086
rect 499806 220048 499866 220766
rect 502425 220763 502491 220766
rect 286409 219874 286475 219877
rect 286409 219872 360210 219874
rect 286409 219816 286414 219872
rect 286470 219816 360210 219872
rect 286409 219814 360210 219816
rect 286409 219811 286475 219814
rect 360150 219776 360210 219814
rect 230381 219602 230447 219605
rect 283557 219602 283623 219605
rect 219390 219600 240212 219602
rect 219390 219544 230386 219600
rect 230442 219544 240212 219600
rect 219390 219542 240212 219544
rect 279956 219600 283623 219602
rect 279956 219544 283562 219600
rect 283618 219544 283623 219600
rect 279956 219542 283623 219544
rect 230381 219539 230447 219542
rect 283557 219539 283623 219542
rect 67541 219330 67607 219333
rect 228357 219330 228423 219333
rect 67541 219328 228423 219330
rect 67541 219272 67546 219328
rect 67602 219272 228362 219328
rect 228418 219272 228423 219328
rect 67541 219270 228423 219272
rect 67541 219267 67607 219270
rect 228357 219267 228423 219270
rect 281809 219058 281875 219061
rect 279956 219056 281875 219058
rect 279956 219000 281814 219056
rect 281870 219000 281875 219056
rect 279956 218998 281875 219000
rect 281809 218995 281875 218998
rect 580441 219058 580507 219061
rect 583520 219058 584960 219148
rect 580441 219056 584960 219058
rect 580441 219000 580446 219056
rect 580502 219000 584960 219056
rect 580441 218998 584960 219000
rect 580441 218995 580507 218998
rect 583520 218908 584960 218998
rect 289445 218786 289511 218789
rect 289445 218784 360210 218786
rect 289445 218728 289450 218784
rect 289506 218728 360210 218784
rect 289445 218726 360210 218728
rect 289445 218723 289511 218726
rect 360150 218688 360210 218726
rect 3550 218588 3556 218652
rect 3620 218650 3626 218652
rect 213126 218650 213132 218652
rect 3620 218590 213132 218650
rect 3620 218588 3626 218590
rect 213126 218588 213132 218590
rect 213196 218588 213202 218652
rect 231577 218514 231643 218517
rect 280889 218514 280955 218517
rect 231577 218512 240212 218514
rect 231577 218456 231582 218512
rect 231638 218456 240212 218512
rect 231577 218454 240212 218456
rect 279956 218512 280955 218514
rect 279956 218456 280894 218512
rect 280950 218456 280955 218512
rect 279956 218454 280955 218456
rect 231577 218451 231643 218454
rect 280889 218451 280955 218454
rect 281717 217970 281783 217973
rect 279956 217968 281783 217970
rect 279956 217912 281722 217968
rect 281778 217912 281783 217968
rect 279956 217910 281783 217912
rect 281717 217907 281783 217910
rect 357525 217834 357591 217837
rect 357525 217832 360210 217834
rect 357525 217776 357530 217832
rect 357586 217776 360210 217832
rect 357525 217774 360210 217776
rect 357525 217771 357591 217774
rect 231577 217698 231643 217701
rect 219390 217696 231643 217698
rect 219390 217640 231582 217696
rect 231638 217640 231643 217696
rect 219390 217638 231643 217640
rect 60089 217290 60155 217293
rect 219390 217290 219450 217638
rect 231577 217635 231643 217638
rect 360150 217600 360210 217774
rect 231669 217426 231735 217429
rect 237465 217426 237531 217429
rect 281901 217426 281967 217429
rect 231669 217424 240212 217426
rect 231669 217368 231674 217424
rect 231730 217368 237470 217424
rect 237526 217368 240212 217424
rect 231669 217366 240212 217368
rect 279956 217424 281967 217426
rect 279956 217368 281906 217424
rect 281962 217368 281967 217424
rect 279956 217366 281967 217368
rect 231669 217363 231735 217366
rect 237465 217363 237531 217366
rect 281901 217363 281967 217366
rect 60089 217288 219450 217290
rect 60089 217232 60094 217288
rect 60150 217232 219450 217288
rect 60089 217230 219450 217232
rect 60089 217227 60155 217230
rect 282269 216882 282335 216885
rect 279956 216880 282335 216882
rect 279956 216824 282274 216880
rect 282330 216824 282335 216880
rect 279956 216822 282335 216824
rect 282269 216819 282335 216822
rect 357525 216610 357591 216613
rect 357525 216608 360210 216610
rect 357525 216552 357530 216608
rect 357586 216552 360210 216608
rect 357525 216550 360210 216552
rect 357525 216547 357591 216550
rect 360150 216512 360210 216550
rect 237373 216338 237439 216341
rect 238569 216338 238635 216341
rect 280705 216338 280771 216341
rect 237373 216336 240212 216338
rect 237373 216280 237378 216336
rect 237434 216280 238574 216336
rect 238630 216280 240212 216336
rect 237373 216278 240212 216280
rect 279956 216336 280771 216338
rect 279956 216280 280710 216336
rect 280766 216280 280771 216336
rect 279956 216278 280771 216280
rect 237373 216275 237439 216278
rect 238569 216275 238635 216278
rect 280705 216275 280771 216278
rect 282729 215794 282795 215797
rect 279956 215792 282795 215794
rect 279956 215736 282734 215792
rect 282790 215736 282795 215792
rect 279956 215734 282795 215736
rect 282729 215731 282795 215734
rect 287881 215522 287947 215525
rect 287881 215520 360210 215522
rect 287881 215464 287886 215520
rect 287942 215464 360210 215520
rect 287881 215462 360210 215464
rect 287881 215459 287947 215462
rect 360150 215424 360210 215462
rect 64137 215386 64203 215389
rect 237373 215386 237439 215389
rect 64137 215384 237439 215386
rect 64137 215328 64142 215384
rect 64198 215328 237378 215384
rect 237434 215328 237439 215384
rect 64137 215326 237439 215328
rect 64137 215323 64203 215326
rect 237373 215323 237439 215326
rect 238661 215250 238727 215253
rect 282177 215250 282243 215253
rect 238661 215248 240212 215250
rect 238661 215192 238666 215248
rect 238722 215192 240212 215248
rect 238661 215190 240212 215192
rect 279956 215248 282243 215250
rect 279956 215192 282182 215248
rect 282238 215192 282243 215248
rect 279956 215190 282243 215192
rect 238661 215187 238727 215190
rect 282177 215187 282243 215190
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 357525 214842 357591 214845
rect 357525 214840 360210 214842
rect 357525 214784 357530 214840
rect 357586 214784 360210 214840
rect 357525 214782 360210 214784
rect 357525 214779 357591 214782
rect 281758 214706 281764 214708
rect 279956 214646 281764 214706
rect 281758 214644 281764 214646
rect 281828 214644 281834 214708
rect 280797 214570 280863 214573
rect 281533 214570 281599 214573
rect 280797 214568 281599 214570
rect 280797 214512 280802 214568
rect 280858 214512 281538 214568
rect 281594 214512 281599 214568
rect 280797 214510 281599 214512
rect 280797 214507 280863 214510
rect 281533 214507 281599 214510
rect 360150 214336 360210 214782
rect 502333 214706 502399 214709
rect 499806 214704 502399 214706
rect 499806 214648 502338 214704
rect 502394 214648 502399 214704
rect 499806 214646 502399 214648
rect 35157 214162 35223 214165
rect 289905 214162 289971 214165
rect 35157 214160 240212 214162
rect 35157 214104 35162 214160
rect 35218 214104 240212 214160
rect 35157 214102 240212 214104
rect 279956 214160 289971 214162
rect 279956 214104 289910 214160
rect 289966 214104 289971 214160
rect 279956 214102 289971 214104
rect 35157 214099 35223 214102
rect 289905 214099 289971 214102
rect 499806 214064 499866 214646
rect 502333 214643 502399 214646
rect 284845 213618 284911 213621
rect 279956 213616 284911 213618
rect 279956 213560 284850 213616
rect 284906 213560 284911 213616
rect 279956 213558 284911 213560
rect 284845 213555 284911 213558
rect 300117 213346 300183 213349
rect 300117 213344 360210 213346
rect 300117 213288 300122 213344
rect 300178 213288 360210 213344
rect 300117 213286 360210 213288
rect 300117 213283 300183 213286
rect 360150 213248 360210 213286
rect 5257 213074 5323 213077
rect 283741 213074 283807 213077
rect 5257 213072 240212 213074
rect 5257 213016 5262 213072
rect 5318 213016 240212 213072
rect 5257 213014 240212 213016
rect 279956 213072 283807 213074
rect 279956 213016 283746 213072
rect 283802 213016 283807 213072
rect 279956 213014 283807 213016
rect 5257 213011 5323 213014
rect 283741 213011 283807 213014
rect 285857 212530 285923 212533
rect 279956 212528 285923 212530
rect 279956 212472 285862 212528
rect 285918 212472 285923 212528
rect 279956 212470 285923 212472
rect 285857 212467 285923 212470
rect 320541 212530 320607 212533
rect 322289 212530 322355 212533
rect 320541 212528 322355 212530
rect 320541 212472 320546 212528
rect 320602 212472 322294 212528
rect 322350 212472 322355 212528
rect 320541 212470 322355 212472
rect 320541 212467 320607 212470
rect 322289 212467 322355 212470
rect 357525 212394 357591 212397
rect 357525 212392 360210 212394
rect 357525 212336 357530 212392
rect 357586 212336 360210 212392
rect 357525 212334 360210 212336
rect 357525 212331 357591 212334
rect 360150 212160 360210 212334
rect 31017 211986 31083 211989
rect 286409 211986 286475 211989
rect 31017 211984 240212 211986
rect 31017 211928 31022 211984
rect 31078 211928 240212 211984
rect 31017 211926 240212 211928
rect 279956 211984 286475 211986
rect 279956 211928 286414 211984
rect 286470 211928 286475 211984
rect 279956 211926 286475 211928
rect 31017 211923 31083 211926
rect 286409 211923 286475 211926
rect 286317 211442 286383 211445
rect 279956 211440 286383 211442
rect 279956 211384 286322 211440
rect 286378 211384 286383 211440
rect 279956 211382 286383 211384
rect 286317 211379 286383 211382
rect 357525 211170 357591 211173
rect 357525 211168 360210 211170
rect 357525 211112 357530 211168
rect 357586 211112 360210 211168
rect 357525 211110 360210 211112
rect 357525 211107 357591 211110
rect 360150 211072 360210 211110
rect 6453 210898 6519 210901
rect 284937 210898 285003 210901
rect 6453 210896 240212 210898
rect 6453 210840 6458 210896
rect 6514 210840 240212 210896
rect 6453 210838 240212 210840
rect 279956 210896 285003 210898
rect 279956 210840 284942 210896
rect 284998 210840 285003 210896
rect 279956 210838 285003 210840
rect 6453 210835 6519 210838
rect 284937 210835 285003 210838
rect 292757 210354 292823 210357
rect 279956 210352 292823 210354
rect 279956 210296 292762 210352
rect 292818 210296 292823 210352
rect 279956 210294 292823 210296
rect 292757 210291 292823 210294
rect 286910 210020 286916 210084
rect 286980 210082 286986 210084
rect 286980 210022 360210 210082
rect 286980 210020 286986 210022
rect 360150 209984 360210 210022
rect 199377 209810 199443 209813
rect 283373 209810 283439 209813
rect 199377 209808 240212 209810
rect 199377 209752 199382 209808
rect 199438 209752 240212 209808
rect 199377 209750 240212 209752
rect 279956 209808 283439 209810
rect 279956 209752 283378 209808
rect 283434 209752 283439 209808
rect 279956 209750 283439 209752
rect 199377 209747 199443 209750
rect 283373 209747 283439 209750
rect 357525 209402 357591 209405
rect 357525 209400 360210 209402
rect 357525 209344 357530 209400
rect 357586 209344 360210 209400
rect 357525 209342 360210 209344
rect 357525 209339 357591 209342
rect 283465 209266 283531 209269
rect 279956 209264 283531 209266
rect 279956 209208 283470 209264
rect 283526 209208 283531 209264
rect 279956 209206 283531 209208
rect 283465 209203 283531 209206
rect 360150 208896 360210 209342
rect 159357 208722 159423 208725
rect 280838 208722 280844 208724
rect 159357 208720 240212 208722
rect 159357 208664 159362 208720
rect 159418 208664 240212 208720
rect 159357 208662 240212 208664
rect 279956 208662 280844 208722
rect 159357 208659 159423 208662
rect 280838 208660 280844 208662
rect 280908 208660 280914 208724
rect 318149 208586 318215 208589
rect 320541 208586 320607 208589
rect 318149 208584 320607 208586
rect 318149 208528 318154 208584
rect 318210 208528 320546 208584
rect 320602 208528 320607 208584
rect 318149 208526 320607 208528
rect 318149 208523 318215 208526
rect 320541 208523 320607 208526
rect 318333 208450 318399 208453
rect 319621 208450 319687 208453
rect 318333 208448 319687 208450
rect 318333 208392 318338 208448
rect 318394 208392 319626 208448
rect 319682 208392 319687 208448
rect 318333 208390 319687 208392
rect 318333 208387 318399 208390
rect 319621 208387 319687 208390
rect 501137 208314 501203 208317
rect 499806 208312 501203 208314
rect 499806 208256 501142 208312
rect 501198 208256 501203 208312
rect 499806 208254 501203 208256
rect 288709 208178 288775 208181
rect 279956 208176 288775 208178
rect 279956 208120 288714 208176
rect 288770 208120 288775 208176
rect 279956 208118 288775 208120
rect 288709 208115 288775 208118
rect 499806 208080 499866 208254
rect 501137 208251 501203 208254
rect 122097 208042 122163 208045
rect 124121 208042 124187 208045
rect 122097 208040 124187 208042
rect 122097 207984 122102 208040
rect 122158 207984 124126 208040
rect 124182 207984 124187 208040
rect 122097 207982 124187 207984
rect 122097 207979 122163 207982
rect 124121 207979 124187 207982
rect 357525 208042 357591 208045
rect 357525 208040 360210 208042
rect 357525 207984 357530 208040
rect 357586 207984 360210 208040
rect 357525 207982 360210 207984
rect 357525 207979 357591 207982
rect 360150 207808 360210 207982
rect 58750 207572 58756 207636
rect 58820 207634 58826 207636
rect 237966 207634 237972 207636
rect 58820 207574 237972 207634
rect 58820 207572 58826 207574
rect 237966 207572 237972 207574
rect 238036 207572 238042 207636
rect 288617 207634 288683 207637
rect 238710 207574 240212 207634
rect 279956 207632 288683 207634
rect 279956 207576 288622 207632
rect 288678 207576 288683 207632
rect 279956 207574 288683 207576
rect 211797 207498 211863 207501
rect 238710 207498 238770 207574
rect 288617 207571 288683 207574
rect 211797 207496 238770 207498
rect 211797 207440 211802 207496
rect 211858 207440 238770 207496
rect 211797 207438 238770 207440
rect 211797 207435 211863 207438
rect 288525 207090 288591 207093
rect 279956 207088 288591 207090
rect 279956 207032 288530 207088
rect 288586 207032 288591 207088
rect 279956 207030 288591 207032
rect 288525 207027 288591 207030
rect 357525 206818 357591 206821
rect 357525 206816 360210 206818
rect 357525 206760 357530 206816
rect 357586 206760 360210 206816
rect 357525 206758 360210 206760
rect 357525 206755 357591 206758
rect 360150 206720 360210 206758
rect 155217 206546 155283 206549
rect 287605 206546 287671 206549
rect 155217 206544 240212 206546
rect 155217 206488 155222 206544
rect 155278 206488 240212 206544
rect 155217 206486 240212 206488
rect 279956 206544 287671 206546
rect 279956 206488 287610 206544
rect 287666 206488 287671 206544
rect 279956 206486 287671 206488
rect 155217 206483 155283 206486
rect 287605 206483 287671 206486
rect 357525 206274 357591 206277
rect 357525 206272 360210 206274
rect 357525 206216 357530 206272
rect 357586 206216 360210 206272
rect 357525 206214 360210 206216
rect 357525 206211 357591 206214
rect 294137 206002 294203 206005
rect 279956 206000 294203 206002
rect 279956 205944 294142 206000
rect 294198 205944 294203 206000
rect 279956 205942 294203 205944
rect 294137 205939 294203 205942
rect 360150 205632 360210 206214
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 126421 205458 126487 205461
rect 286501 205458 286567 205461
rect 126421 205456 240212 205458
rect 126421 205400 126426 205456
rect 126482 205400 240212 205456
rect 126421 205398 240212 205400
rect 279956 205456 286567 205458
rect 279956 205400 286506 205456
rect 286562 205400 286567 205456
rect 279956 205398 286567 205400
rect 126421 205395 126487 205398
rect 286501 205395 286567 205398
rect 357525 205050 357591 205053
rect 357525 205048 360210 205050
rect 357525 204992 357530 205048
rect 357586 204992 360210 205048
rect 357525 204990 360210 204992
rect 357525 204987 357591 204990
rect 282126 204914 282132 204916
rect 279956 204854 282132 204914
rect 282126 204852 282132 204854
rect 282196 204852 282202 204916
rect 360150 204544 360210 204990
rect 126237 204370 126303 204373
rect 287513 204370 287579 204373
rect 126237 204368 240212 204370
rect 126237 204312 126242 204368
rect 126298 204312 240212 204368
rect 126237 204310 240212 204312
rect 279956 204368 287579 204370
rect 279956 204312 287518 204368
rect 287574 204312 287579 204368
rect 279956 204310 287579 204312
rect 126237 204307 126303 204310
rect 287513 204307 287579 204310
rect 124121 204098 124187 204101
rect 129089 204098 129155 204101
rect 124121 204096 129155 204098
rect 124121 204040 124126 204096
rect 124182 204040 129094 204096
rect 129150 204040 129155 204096
rect 124121 204038 129155 204040
rect 124121 204035 124187 204038
rect 129089 204035 129155 204038
rect 284661 203826 284727 203829
rect 279956 203824 284727 203826
rect 279956 203768 284666 203824
rect 284722 203768 284727 203824
rect 279956 203766 284727 203768
rect 284661 203763 284727 203766
rect 357525 203826 357591 203829
rect 357525 203824 360210 203826
rect 357525 203768 357530 203824
rect 357586 203768 360210 203824
rect 357525 203766 360210 203768
rect 357525 203763 357591 203766
rect 360150 203456 360210 203766
rect 126605 203282 126671 203285
rect 281625 203282 281691 203285
rect 126605 203280 240212 203282
rect 126605 203224 126610 203280
rect 126666 203224 240212 203280
rect 126605 203222 240212 203224
rect 279956 203280 281691 203282
rect 279956 203224 281630 203280
rect 281686 203224 281691 203280
rect 279956 203222 281691 203224
rect 126605 203219 126671 203222
rect 281625 203219 281691 203222
rect 287421 202738 287487 202741
rect 499665 202738 499731 202741
rect 279956 202736 287487 202738
rect 279956 202680 287426 202736
rect 287482 202680 287487 202736
rect 279956 202678 287487 202680
rect 287421 202675 287487 202678
rect 499622 202736 499731 202738
rect 499622 202680 499670 202736
rect 499726 202680 499731 202736
rect 499622 202675 499731 202680
rect 315389 202466 315455 202469
rect 315389 202464 360210 202466
rect 315389 202408 315394 202464
rect 315450 202408 360210 202464
rect 315389 202406 360210 202408
rect 315389 202403 315455 202406
rect 360150 202368 360210 202406
rect 57513 202194 57579 202197
rect 233877 202194 233943 202197
rect 287881 202194 287947 202197
rect 57513 202192 233943 202194
rect 57513 202136 57518 202192
rect 57574 202136 233882 202192
rect 233938 202136 233943 202192
rect 57513 202134 233943 202136
rect 57513 202131 57579 202134
rect 233877 202131 233943 202134
rect 238710 202134 240212 202194
rect 279956 202192 287947 202194
rect 279956 202136 287886 202192
rect 287942 202136 287947 202192
rect 279956 202134 287947 202136
rect 222837 202058 222903 202061
rect 238710 202058 238770 202134
rect 287881 202131 287947 202134
rect 499622 202096 499682 202675
rect 222837 202056 238770 202058
rect -960 201922 480 202012
rect 222837 202000 222842 202056
rect 222898 202000 238770 202056
rect 222837 201998 238770 202000
rect 222837 201995 222903 201998
rect 234654 201922 234660 201924
rect -960 201862 234660 201922
rect -960 201772 480 201862
rect 234654 201860 234660 201862
rect 234724 201860 234730 201924
rect 287329 201650 287395 201653
rect 279956 201648 287395 201650
rect 279956 201592 287334 201648
rect 287390 201592 287395 201648
rect 279956 201590 287395 201592
rect 287329 201587 287395 201590
rect 357525 201378 357591 201381
rect 357525 201376 360210 201378
rect 357525 201320 357530 201376
rect 357586 201320 360210 201376
rect 357525 201318 360210 201320
rect 357525 201315 357591 201318
rect 360150 201280 360210 201318
rect 209037 201106 209103 201109
rect 287053 201106 287119 201109
rect 209037 201104 240212 201106
rect 209037 201048 209042 201104
rect 209098 201048 240212 201104
rect 209037 201046 240212 201048
rect 279956 201104 287119 201106
rect 279956 201048 287058 201104
rect 287114 201048 287119 201104
rect 279956 201046 287119 201048
rect 209037 201043 209103 201046
rect 287053 201043 287119 201046
rect 357525 200834 357591 200837
rect 357525 200832 360210 200834
rect 357525 200776 357530 200832
rect 357586 200776 360210 200832
rect 357525 200774 360210 200776
rect 357525 200771 357591 200774
rect 287237 200562 287303 200565
rect 279956 200560 287303 200562
rect 279956 200504 287242 200560
rect 287298 200504 287303 200560
rect 279956 200502 287303 200504
rect 287237 200499 287303 200502
rect 360150 200192 360210 200774
rect 228357 200018 228423 200021
rect 285806 200018 285812 200020
rect 228357 200016 240212 200018
rect 228357 199960 228362 200016
rect 228418 199960 240212 200016
rect 228357 199958 240212 199960
rect 279956 199958 285812 200018
rect 228357 199955 228423 199958
rect 285806 199956 285812 199958
rect 285876 199956 285882 200020
rect 291469 199474 291535 199477
rect 279956 199472 291535 199474
rect 279956 199416 291474 199472
rect 291530 199416 291535 199472
rect 279956 199414 291535 199416
rect 291469 199411 291535 199414
rect 57421 199338 57487 199341
rect 227161 199338 227227 199341
rect 57421 199336 227227 199338
rect 57421 199280 57426 199336
rect 57482 199280 227166 199336
rect 227222 199280 227227 199336
rect 57421 199278 227227 199280
rect 57421 199275 57487 199278
rect 227161 199275 227227 199278
rect 304257 199202 304323 199205
rect 304257 199200 360210 199202
rect 304257 199144 304262 199200
rect 304318 199144 360210 199200
rect 304257 199142 360210 199144
rect 304257 199139 304323 199142
rect 360150 199104 360210 199142
rect 226977 198930 227043 198933
rect 281574 198930 281580 198932
rect 226977 198928 240212 198930
rect 226977 198872 226982 198928
rect 227038 198872 240212 198928
rect 226977 198870 240212 198872
rect 279956 198870 281580 198930
rect 226977 198867 227043 198870
rect 281574 198868 281580 198870
rect 281644 198868 281650 198932
rect 316769 198794 316835 198797
rect 318333 198794 318399 198797
rect 316769 198792 318399 198794
rect 316769 198736 316774 198792
rect 316830 198736 318338 198792
rect 318394 198736 318399 198792
rect 316769 198734 318399 198736
rect 316769 198731 316835 198734
rect 318333 198731 318399 198734
rect 282361 198386 282427 198389
rect 279956 198384 282427 198386
rect 279956 198328 282366 198384
rect 282422 198328 282427 198384
rect 279956 198326 282427 198328
rect 282361 198323 282427 198326
rect 57697 198114 57763 198117
rect 216121 198114 216187 198117
rect 57697 198112 216187 198114
rect 57697 198056 57702 198112
rect 57758 198056 216126 198112
rect 216182 198056 216187 198112
rect 57697 198054 216187 198056
rect 57697 198051 57763 198054
rect 216121 198051 216187 198054
rect 287697 198114 287763 198117
rect 287697 198112 360210 198114
rect 287697 198056 287702 198112
rect 287758 198056 360210 198112
rect 287697 198054 360210 198056
rect 287697 198051 287763 198054
rect 360150 198016 360210 198054
rect 60181 197978 60247 197981
rect 237465 197978 237531 197981
rect 60181 197976 237531 197978
rect 60181 197920 60186 197976
rect 60242 197920 237470 197976
rect 237526 197920 237531 197976
rect 60181 197918 237531 197920
rect 60181 197915 60247 197918
rect 237465 197915 237531 197918
rect 215937 197842 216003 197845
rect 281942 197842 281948 197844
rect 215937 197840 240212 197842
rect 215937 197784 215942 197840
rect 215998 197784 240212 197840
rect 215937 197782 240212 197784
rect 279956 197782 281948 197842
rect 215937 197779 216003 197782
rect 281942 197780 281948 197782
rect 282012 197780 282018 197844
rect 282545 197434 282611 197437
rect 282913 197434 282979 197437
rect 282545 197432 282979 197434
rect 282545 197376 282550 197432
rect 282606 197376 282918 197432
rect 282974 197376 282979 197432
rect 282545 197374 282979 197376
rect 282545 197371 282611 197374
rect 282913 197371 282979 197374
rect 280654 197298 280660 197300
rect 279956 197238 280660 197298
rect 280654 197236 280660 197238
rect 280724 197236 280730 197300
rect 291837 197026 291903 197029
rect 291837 197024 360210 197026
rect 291837 196968 291842 197024
rect 291898 196968 360210 197024
rect 291837 196966 360210 196968
rect 291837 196963 291903 196966
rect 360150 196928 360210 196966
rect 214557 196754 214623 196757
rect 284702 196754 284708 196756
rect 214557 196752 240212 196754
rect 214557 196696 214562 196752
rect 214618 196696 240212 196752
rect 214557 196694 240212 196696
rect 279956 196694 284708 196754
rect 214557 196691 214623 196694
rect 284702 196692 284708 196694
rect 284772 196692 284778 196756
rect 501229 196754 501295 196757
rect 499806 196752 501295 196754
rect 499806 196696 501234 196752
rect 501290 196696 501295 196752
rect 499806 196694 501295 196696
rect 58985 196618 59051 196621
rect 238201 196618 238267 196621
rect 58985 196616 238267 196618
rect 58985 196560 58990 196616
rect 59046 196560 238206 196616
rect 238262 196560 238267 196616
rect 58985 196558 238267 196560
rect 58985 196555 59051 196558
rect 238201 196555 238267 196558
rect 288893 196210 288959 196213
rect 279956 196208 288959 196210
rect 279956 196152 288898 196208
rect 288954 196152 288959 196208
rect 279956 196150 288959 196152
rect 288893 196147 288959 196150
rect 499806 196112 499866 196694
rect 501229 196691 501295 196694
rect 129089 196074 129155 196077
rect 130285 196074 130351 196077
rect 318149 196074 318215 196077
rect 129089 196072 130351 196074
rect 129089 196016 129094 196072
rect 129150 196016 130290 196072
rect 130346 196016 130351 196072
rect 129089 196014 130351 196016
rect 129089 196011 129155 196014
rect 130285 196011 130351 196014
rect 310470 196072 318215 196074
rect 310470 196016 318154 196072
rect 318210 196016 318215 196072
rect 310470 196014 318215 196016
rect 309041 195938 309107 195941
rect 310470 195938 310530 196014
rect 318149 196011 318215 196014
rect 309041 195936 310530 195938
rect 309041 195880 309046 195936
rect 309102 195880 310530 195936
rect 309041 195878 310530 195880
rect 357525 195938 357591 195941
rect 357525 195936 360210 195938
rect 357525 195880 357530 195936
rect 357586 195880 360210 195936
rect 357525 195878 360210 195880
rect 309041 195875 309107 195878
rect 357525 195875 357591 195878
rect 360150 195840 360210 195878
rect 188337 195666 188403 195669
rect 289077 195666 289143 195669
rect 188337 195664 240212 195666
rect 188337 195608 188342 195664
rect 188398 195608 240212 195664
rect 188337 195606 240212 195608
rect 279956 195664 289143 195666
rect 279956 195608 289082 195664
rect 289138 195608 289143 195664
rect 279956 195606 289143 195608
rect 188337 195603 188403 195606
rect 289077 195603 289143 195606
rect 60590 195196 60596 195260
rect 60660 195258 60666 195260
rect 238150 195258 238156 195260
rect 60660 195198 238156 195258
rect 60660 195196 60666 195198
rect 238150 195196 238156 195198
rect 238220 195196 238226 195260
rect 288801 195122 288867 195125
rect 279956 195120 288867 195122
rect 279956 195064 288806 195120
rect 288862 195064 288867 195120
rect 279956 195062 288867 195064
rect 288801 195059 288867 195062
rect 220077 194578 220143 194581
rect 288985 194578 289051 194581
rect 220077 194576 240212 194578
rect 220077 194520 220082 194576
rect 220138 194520 240212 194576
rect 220077 194518 240212 194520
rect 279956 194576 289051 194578
rect 279956 194520 288990 194576
rect 289046 194520 289051 194576
rect 279956 194518 289051 194520
rect 220077 194515 220143 194518
rect 288985 194515 289051 194518
rect 58893 194034 58959 194037
rect 238109 194034 238175 194037
rect 284886 194034 284892 194036
rect 58893 194032 238175 194034
rect 58893 193976 58898 194032
rect 58954 193976 238114 194032
rect 238170 193976 238175 194032
rect 58893 193974 238175 193976
rect 279956 193974 284892 194034
rect 58893 193971 58959 193974
rect 238109 193971 238175 193974
rect 284886 193972 284892 193974
rect 284956 193972 284962 194036
rect 18454 193836 18460 193900
rect 18524 193898 18530 193900
rect 237966 193898 237972 193900
rect 18524 193838 237972 193898
rect 18524 193836 18530 193838
rect 237966 193836 237972 193838
rect 238036 193836 238042 193900
rect 233877 193490 233943 193493
rect 283649 193490 283715 193493
rect 233877 193488 240212 193490
rect 233877 193432 233882 193488
rect 233938 193432 240212 193488
rect 233877 193430 240212 193432
rect 279956 193488 283715 193490
rect 279956 193432 283654 193488
rect 283710 193432 283715 193488
rect 279956 193430 283715 193432
rect 233877 193427 233943 193430
rect 283649 193427 283715 193430
rect 130285 193218 130351 193221
rect 131481 193218 131547 193221
rect 130285 193216 131547 193218
rect 130285 193160 130290 193216
rect 130346 193160 131486 193216
rect 131542 193160 131547 193216
rect 130285 193158 131547 193160
rect 130285 193155 130351 193158
rect 131481 193155 131547 193158
rect 280061 192946 280127 192949
rect 279956 192944 280127 192946
rect 279956 192888 280066 192944
rect 280122 192888 280127 192944
rect 279956 192886 280127 192888
rect 280061 192883 280127 192886
rect 59077 192674 59143 192677
rect 238017 192674 238083 192677
rect 59077 192672 238083 192674
rect 59077 192616 59082 192672
rect 59138 192616 238022 192672
rect 238078 192616 238083 192672
rect 59077 192614 238083 192616
rect 59077 192611 59143 192614
rect 238017 192611 238083 192614
rect 15694 192476 15700 192540
rect 15764 192538 15770 192540
rect 237414 192538 237420 192540
rect 15764 192478 237420 192538
rect 15764 192476 15770 192478
rect 237414 192476 237420 192478
rect 237484 192476 237490 192540
rect 580533 192538 580599 192541
rect 583520 192538 584960 192628
rect 580533 192536 584960 192538
rect 580533 192480 580538 192536
rect 580594 192480 584960 192536
rect 580533 192478 584960 192480
rect 580533 192475 580599 192478
rect 224217 192402 224283 192405
rect 282821 192402 282887 192405
rect 224217 192400 240212 192402
rect 224217 192344 224222 192400
rect 224278 192344 240212 192400
rect 224217 192342 240212 192344
rect 279956 192400 282887 192402
rect 279956 192344 282826 192400
rect 282882 192344 282887 192400
rect 583520 192388 584960 192478
rect 279956 192342 282887 192344
rect 224217 192339 224283 192342
rect 282821 192339 282887 192342
rect 283230 191858 283236 191860
rect 279956 191798 283236 191858
rect 283230 191796 283236 191798
rect 283300 191796 283306 191860
rect 309041 191858 309107 191861
rect 306330 191856 309107 191858
rect 306330 191800 309046 191856
rect 309102 191800 309107 191856
rect 306330 191798 309107 191800
rect 303521 191722 303587 191725
rect 306330 191722 306390 191798
rect 309041 191795 309107 191798
rect 303521 191720 306390 191722
rect 303521 191664 303526 191720
rect 303582 191664 306390 191720
rect 303521 191662 306390 191664
rect 303521 191659 303587 191662
rect 206277 191314 206343 191317
rect 281022 191314 281028 191316
rect 206277 191312 240212 191314
rect 206277 191256 206282 191312
rect 206338 191256 240212 191312
rect 206277 191254 240212 191256
rect 279956 191254 281028 191314
rect 206277 191251 206343 191254
rect 281022 191252 281028 191254
rect 281092 191252 281098 191316
rect 57881 191178 57947 191181
rect 220353 191178 220419 191181
rect 57881 191176 220419 191178
rect 57881 191120 57886 191176
rect 57942 191120 220358 191176
rect 220414 191120 220419 191176
rect 57881 191118 220419 191120
rect 57881 191115 57947 191118
rect 220353 191115 220419 191118
rect 26734 190980 26740 191044
rect 26804 191042 26810 191044
rect 238150 191042 238156 191044
rect 26804 190982 238156 191042
rect 26804 190980 26810 190982
rect 238150 190980 238156 190982
rect 238220 190980 238226 191044
rect 320817 190770 320883 190773
rect 279956 190768 320883 190770
rect 279956 190712 320822 190768
rect 320878 190712 320883 190768
rect 279956 190710 320883 190712
rect 320817 190707 320883 190710
rect 501045 190362 501111 190365
rect 499806 190360 501111 190362
rect 499806 190304 501050 190360
rect 501106 190304 501111 190360
rect 499806 190302 501111 190304
rect 146937 190226 147003 190229
rect 302918 190226 302924 190228
rect 146937 190224 240212 190226
rect 146937 190168 146942 190224
rect 146998 190168 240212 190224
rect 146937 190166 240212 190168
rect 279956 190166 302924 190226
rect 146937 190163 147003 190166
rect 302918 190164 302924 190166
rect 302988 190164 302994 190228
rect 499806 190128 499866 190302
rect 501045 190299 501111 190302
rect 57462 189620 57468 189684
rect 57532 189682 57538 189684
rect 210550 189682 210556 189684
rect 57532 189622 210556 189682
rect 57532 189620 57538 189622
rect 210550 189620 210556 189622
rect 210620 189620 210626 189684
rect 346894 189682 346900 189684
rect 279956 189622 346900 189682
rect 346894 189620 346900 189622
rect 346964 189620 346970 189684
rect 210417 189138 210483 189141
rect 345606 189138 345612 189140
rect 210417 189136 240212 189138
rect 210417 189080 210422 189136
rect 210478 189080 240212 189136
rect 210417 189078 240212 189080
rect 279956 189078 345612 189138
rect 210417 189075 210483 189078
rect 345606 189076 345612 189078
rect 345676 189076 345682 189140
rect -960 188866 480 188956
rect 3366 188866 3372 188868
rect -960 188806 3372 188866
rect -960 188716 480 188806
rect 3366 188804 3372 188806
rect 3436 188804 3442 188868
rect 327758 188594 327764 188596
rect 279956 188534 327764 188594
rect 327758 188532 327764 188534
rect 327828 188532 327834 188596
rect 315389 188458 315455 188461
rect 316769 188458 316835 188461
rect 315389 188456 316835 188458
rect 315389 188400 315394 188456
rect 315450 188400 316774 188456
rect 316830 188400 316835 188456
rect 315389 188398 316835 188400
rect 315389 188395 315455 188398
rect 316769 188395 316835 188398
rect 22686 188260 22692 188324
rect 22756 188322 22762 188324
rect 238334 188322 238340 188324
rect 22756 188262 238340 188322
rect 22756 188260 22762 188262
rect 238334 188260 238340 188262
rect 238404 188260 238410 188324
rect 140037 188050 140103 188053
rect 290774 188050 290780 188052
rect 140037 188048 240212 188050
rect 140037 187992 140042 188048
rect 140098 187992 240212 188048
rect 140037 187990 240212 187992
rect 279956 187990 290780 188050
rect 140037 187987 140103 187990
rect 290774 187988 290780 187990
rect 290844 187988 290850 188052
rect 238201 187914 238267 187917
rect 238661 187914 238727 187917
rect 219390 187912 238727 187914
rect 219390 187856 238206 187912
rect 238262 187856 238666 187912
rect 238722 187856 238727 187912
rect 219390 187854 238727 187856
rect 59169 187778 59235 187781
rect 219390 187778 219450 187854
rect 238201 187851 238267 187854
rect 238661 187851 238727 187854
rect 59169 187776 219450 187778
rect 59169 187720 59174 187776
rect 59230 187720 219450 187776
rect 59169 187718 219450 187720
rect 59169 187715 59235 187718
rect 237414 187716 237420 187780
rect 237484 187778 237490 187780
rect 238477 187778 238543 187781
rect 237484 187776 238543 187778
rect 237484 187720 238482 187776
rect 238538 187720 238543 187776
rect 237484 187718 238543 187720
rect 237484 187716 237490 187718
rect 238477 187715 238543 187718
rect 298737 187778 298803 187781
rect 303521 187778 303587 187781
rect 298737 187776 303587 187778
rect 298737 187720 298742 187776
rect 298798 187720 303526 187776
rect 303582 187720 303587 187776
rect 298737 187718 303587 187720
rect 298737 187715 298803 187718
rect 303521 187715 303587 187718
rect 313958 187506 313964 187508
rect 279956 187446 313964 187506
rect 313958 187444 313964 187446
rect 314028 187444 314034 187508
rect 55121 187370 55187 187373
rect 113817 187370 113883 187373
rect 55121 187368 113883 187370
rect 55121 187312 55126 187368
rect 55182 187312 113822 187368
rect 113878 187312 113883 187368
rect 55121 187310 113883 187312
rect 55121 187307 55187 187310
rect 113817 187307 113883 187310
rect 57789 187234 57855 187237
rect 175917 187234 175983 187237
rect 57789 187232 175983 187234
rect 57789 187176 57794 187232
rect 57850 187176 175922 187232
rect 175978 187176 175983 187232
rect 57789 187174 175983 187176
rect 57789 187171 57855 187174
rect 175917 187171 175983 187174
rect 92381 187098 92447 187101
rect 229737 187098 229803 187101
rect 92381 187096 229803 187098
rect 92381 187040 92386 187096
rect 92442 187040 229742 187096
rect 229798 187040 229803 187096
rect 92381 187038 229803 187040
rect 92381 187035 92447 187038
rect 229737 187035 229803 187038
rect 57646 186900 57652 186964
rect 57716 186962 57722 186964
rect 197854 186962 197860 186964
rect 57716 186902 197860 186962
rect 57716 186900 57722 186902
rect 197854 186900 197860 186902
rect 197924 186900 197930 186964
rect 197997 186962 198063 186965
rect 338614 186962 338620 186964
rect 197997 186960 240212 186962
rect 197997 186904 198002 186960
rect 198058 186904 240212 186960
rect 197997 186902 240212 186904
rect 279956 186902 338620 186962
rect 197997 186899 198063 186902
rect 338614 186900 338620 186902
rect 338684 186900 338690 186964
rect 300158 186418 300164 186420
rect 279956 186358 300164 186418
rect 300158 186356 300164 186358
rect 300228 186356 300234 186420
rect 45461 185874 45527 185877
rect 334566 185874 334572 185876
rect 45461 185872 240212 185874
rect 45461 185816 45466 185872
rect 45522 185816 240212 185872
rect 45461 185814 240212 185816
rect 279956 185814 334572 185874
rect 45461 185811 45527 185814
rect 334566 185812 334572 185814
rect 334636 185812 334642 185876
rect 58801 185738 58867 185741
rect 238293 185738 238359 185741
rect 58801 185736 238359 185738
rect 58801 185680 58806 185736
rect 58862 185680 238298 185736
rect 238354 185680 238359 185736
rect 58801 185678 238359 185680
rect 58801 185675 58867 185678
rect 238293 185675 238359 185678
rect 3366 185540 3372 185604
rect 3436 185602 3442 185604
rect 235390 185602 235396 185604
rect 3436 185542 235396 185602
rect 3436 185540 3442 185542
rect 235390 185540 235396 185542
rect 235460 185540 235466 185604
rect 57605 185466 57671 185469
rect 61469 185466 61535 185469
rect 57605 185464 61535 185466
rect 57605 185408 57610 185464
rect 57666 185408 61474 185464
rect 61530 185408 61535 185464
rect 57605 185406 61535 185408
rect 57605 185403 57671 185406
rect 61469 185403 61535 185406
rect 57329 185330 57395 185333
rect 64137 185330 64203 185333
rect 291878 185330 291884 185332
rect 57329 185328 64203 185330
rect 57329 185272 57334 185328
rect 57390 185272 64142 185328
rect 64198 185272 64203 185328
rect 57329 185270 64203 185272
rect 279956 185270 291884 185330
rect 57329 185267 57395 185270
rect 64137 185267 64203 185270
rect 291878 185268 291884 185270
rect 291948 185268 291954 185332
rect 48221 185058 48287 185061
rect 238017 185058 238083 185061
rect 48221 185056 238083 185058
rect 48221 185000 48226 185056
rect 48282 185000 238022 185056
rect 238078 185000 238083 185056
rect 48221 184998 238083 185000
rect 48221 184995 48287 184998
rect 238017 184995 238083 184998
rect 57145 184922 57211 184925
rect 61377 184922 61443 184925
rect 57145 184920 61443 184922
rect 57145 184864 57150 184920
rect 57206 184864 61382 184920
rect 61438 184864 61443 184920
rect 57145 184862 61443 184864
rect 57145 184859 57211 184862
rect 61377 184859 61443 184862
rect 131481 184922 131547 184925
rect 133137 184922 133203 184925
rect 503621 184922 503687 184925
rect 131481 184920 133203 184922
rect 131481 184864 131486 184920
rect 131542 184864 133142 184920
rect 133198 184864 133203 184920
rect 131481 184862 133203 184864
rect 131481 184859 131547 184862
rect 133137 184859 133203 184862
rect 499806 184920 503687 184922
rect 499806 184864 503626 184920
rect 503682 184864 503687 184920
rect 499806 184862 503687 184864
rect 41873 184786 41939 184789
rect 319294 184786 319300 184788
rect 41873 184784 240212 184786
rect 41873 184728 41878 184784
rect 41934 184728 240212 184784
rect 41873 184726 240212 184728
rect 279956 184726 319300 184786
rect 41873 184723 41939 184726
rect 319294 184724 319300 184726
rect 319364 184724 319370 184788
rect 3366 184452 3372 184516
rect 3436 184514 3442 184516
rect 134374 184514 134380 184516
rect 3436 184454 134380 184514
rect 3436 184452 3442 184454
rect 134374 184452 134380 184454
rect 134444 184452 134450 184516
rect 298870 184242 298876 184244
rect 279956 184182 298876 184242
rect 298870 184180 298876 184182
rect 298940 184180 298946 184244
rect 499806 184144 499866 184862
rect 503621 184859 503687 184862
rect 137277 183698 137343 183701
rect 342846 183698 342852 183700
rect 137277 183696 240212 183698
rect 137277 183640 137282 183696
rect 137338 183640 240212 183696
rect 137277 183638 240212 183640
rect 279956 183638 342852 183698
rect 137277 183635 137343 183638
rect 342846 183636 342852 183638
rect 342916 183636 342922 183700
rect 349654 183154 349660 183156
rect 279956 183094 349660 183154
rect 349654 183092 349660 183094
rect 349724 183092 349730 183156
rect 213177 182610 213243 182613
rect 335854 182610 335860 182612
rect 213177 182608 240212 182610
rect 213177 182552 213182 182608
rect 213238 182552 240212 182608
rect 213177 182550 240212 182552
rect 279956 182550 335860 182610
rect 213177 182547 213243 182550
rect 335854 182548 335860 182550
rect 335924 182548 335930 182612
rect 59670 182004 59676 182068
rect 59740 182066 59746 182068
rect 59905 182066 59971 182069
rect 294822 182066 294828 182068
rect 59740 182064 59971 182066
rect 59740 182008 59910 182064
rect 59966 182008 59971 182064
rect 59740 182006 59971 182008
rect 279956 182006 294828 182066
rect 59740 182004 59746 182006
rect 59905 182003 59971 182006
rect 294822 182004 294828 182006
rect 294892 182004 294898 182068
rect 60406 181732 60412 181796
rect 60476 181732 60482 181796
rect 355685 181794 355751 181797
rect 530577 181794 530643 181797
rect 355685 181792 530643 181794
rect 355685 181736 355690 181792
rect 355746 181736 530582 181792
rect 530638 181736 530643 181792
rect 355685 181734 530643 181736
rect 355685 181731 355751 181734
rect 530577 181731 530643 181734
rect 238109 181522 238175 181525
rect 307150 181522 307156 181524
rect 238109 181520 240212 181522
rect 238109 181464 238114 181520
rect 238170 181464 240212 181520
rect 238109 181462 240212 181464
rect 279956 181462 307156 181522
rect 238109 181459 238175 181462
rect 307150 181460 307156 181462
rect 307220 181460 307226 181524
rect 407614 181324 407620 181388
rect 407684 181386 407690 181388
rect 500953 181386 501019 181389
rect 407684 181384 501019 181386
rect 407684 181328 500958 181384
rect 501014 181328 501019 181384
rect 407684 181326 501019 181328
rect 407684 181324 407690 181326
rect 500953 181323 501019 181326
rect 214598 180978 214604 180980
rect 124844 180918 214604 180978
rect 214598 180916 214604 180918
rect 214668 180916 214674 180980
rect 353886 180978 353892 180980
rect 279956 180918 353892 180978
rect 353886 180916 353892 180918
rect 353956 180916 353962 180980
rect 359549 180570 359615 180573
rect 387977 180570 388043 180573
rect 359549 180568 388043 180570
rect 359549 180512 359554 180568
rect 359610 180512 387982 180568
rect 388038 180512 388043 180568
rect 359549 180510 388043 180512
rect 359549 180507 359615 180510
rect 387977 180507 388043 180510
rect 478045 180570 478111 180573
rect 525742 180570 525748 180572
rect 478045 180568 525748 180570
rect 478045 180512 478050 180568
rect 478106 180512 525748 180568
rect 478045 180510 525748 180512
rect 478045 180507 478111 180510
rect 525742 180508 525748 180510
rect 525812 180508 525818 180572
rect 151077 180434 151143 180437
rect 309726 180434 309732 180436
rect 151077 180432 240212 180434
rect 151077 180376 151082 180432
rect 151138 180376 240212 180432
rect 151077 180374 240212 180376
rect 279956 180374 309732 180434
rect 151077 180371 151143 180374
rect 309726 180372 309732 180374
rect 309796 180372 309802 180436
rect 336365 180434 336431 180437
rect 392025 180434 392091 180437
rect 336365 180432 392091 180434
rect 336365 180376 336370 180432
rect 336426 180376 392030 180432
rect 392086 180376 392091 180432
rect 336365 180374 392091 180376
rect 336365 180371 336431 180374
rect 392025 180371 392091 180374
rect 461853 180434 461919 180437
rect 535494 180434 535500 180436
rect 461853 180432 535500 180434
rect 461853 180376 461858 180432
rect 461914 180376 535500 180432
rect 461853 180374 535500 180376
rect 461853 180371 461919 180374
rect 535494 180372 535500 180374
rect 535564 180372 535570 180436
rect 347589 180298 347655 180301
rect 405181 180298 405247 180301
rect 347589 180296 405247 180298
rect 347589 180240 347594 180296
rect 347650 180240 405186 180296
rect 405242 180240 405247 180296
rect 347589 180238 405247 180240
rect 347589 180235 347655 180238
rect 405181 180235 405247 180238
rect 454769 180298 454835 180301
rect 529974 180298 529980 180300
rect 454769 180296 529980 180298
rect 454769 180240 454774 180296
rect 454830 180240 529980 180296
rect 454769 180238 529980 180240
rect 454769 180235 454835 180238
rect 529974 180236 529980 180238
rect 530044 180236 530050 180300
rect 359917 180162 359983 180165
rect 421373 180162 421439 180165
rect 359917 180160 421439 180162
rect 359917 180104 359922 180160
rect 359978 180104 421378 180160
rect 421434 180104 421439 180160
rect 359917 180102 421439 180104
rect 359917 180099 359983 180102
rect 421373 180099 421439 180102
rect 441613 180162 441679 180165
rect 517830 180162 517836 180164
rect 441613 180160 470610 180162
rect 441613 180104 441618 180160
rect 441674 180104 470610 180160
rect 441613 180102 470610 180104
rect 441613 180099 441679 180102
rect 470550 180026 470610 180102
rect 477174 180102 517836 180162
rect 477174 180026 477234 180102
rect 517830 180100 517836 180102
rect 517900 180100 517906 180164
rect 514886 180026 514892 180028
rect 470550 179966 477234 180026
rect 477358 179966 514892 180026
rect 57646 179828 57652 179892
rect 57716 179890 57722 179892
rect 351126 179890 351132 179892
rect 57716 179830 60076 179890
rect 279956 179830 351132 179890
rect 57716 179828 57722 179830
rect 351126 179828 351132 179830
rect 351196 179828 351202 179892
rect 407757 179890 407823 179893
rect 407757 179888 470610 179890
rect 407757 179832 407762 179888
rect 407818 179832 470610 179888
rect 407757 179830 470610 179832
rect 407757 179827 407823 179830
rect 470550 179618 470610 179830
rect 473997 179754 474063 179757
rect 477358 179754 477418 179966
rect 514886 179964 514892 179966
rect 514956 179964 514962 180028
rect 499757 179890 499823 179893
rect 473997 179752 477418 179754
rect 473997 179696 474002 179752
rect 474058 179696 477418 179752
rect 473997 179694 477418 179696
rect 480210 179888 499823 179890
rect 480210 179832 499762 179888
rect 499818 179832 499823 179888
rect 480210 179830 499823 179832
rect 473997 179691 474063 179694
rect 480210 179618 480270 179830
rect 499757 179827 499823 179830
rect 470550 179558 480270 179618
rect 57881 179484 57947 179485
rect 57830 179420 57836 179484
rect 57900 179482 57947 179484
rect 57900 179480 57992 179482
rect 57942 179424 57992 179480
rect 57900 179422 57992 179424
rect 57900 179420 57947 179422
rect 57881 179419 57947 179420
rect 141417 179346 141483 179349
rect 341885 179346 341951 179349
rect 410241 179346 410307 179349
rect 141417 179344 240212 179346
rect 124814 179210 124874 179316
rect 141417 179288 141422 179344
rect 141478 179288 240212 179344
rect 141417 179286 240212 179288
rect 279956 179286 283298 179346
rect 141417 179283 141483 179286
rect 214414 179210 214420 179212
rect 124814 179150 214420 179210
rect 214414 179148 214420 179150
rect 214484 179148 214490 179212
rect 283238 179077 283298 179286
rect 341885 179344 410307 179346
rect 341885 179288 341890 179344
rect 341946 179288 410246 179344
rect 410302 179288 410307 179344
rect 341885 179286 410307 179288
rect 341885 179283 341951 179286
rect 410241 179283 410307 179286
rect 415301 179346 415367 179349
rect 504030 179346 504036 179348
rect 415301 179344 504036 179346
rect 415301 179288 415306 179344
rect 415362 179288 504036 179344
rect 415301 179286 504036 179288
rect 415301 179283 415367 179286
rect 504030 179284 504036 179286
rect 504100 179284 504106 179348
rect 334750 179148 334756 179212
rect 334820 179210 334826 179212
rect 583520 179210 584960 179300
rect 334820 179150 584960 179210
rect 334820 179148 334826 179150
rect 283238 179072 283347 179077
rect 283238 179016 283286 179072
rect 283342 179016 283347 179072
rect 283238 179014 283347 179016
rect 283281 179011 283347 179014
rect 338941 179074 339007 179077
rect 411253 179074 411319 179077
rect 338941 179072 411319 179074
rect 338941 179016 338946 179072
rect 339002 179016 411258 179072
rect 411314 179016 411319 179072
rect 338941 179014 411319 179016
rect 338941 179011 339007 179014
rect 411253 179011 411319 179014
rect 462865 179074 462931 179077
rect 510654 179074 510660 179076
rect 462865 179072 510660 179074
rect 462865 179016 462870 179072
rect 462926 179016 510660 179072
rect 462865 179014 510660 179016
rect 462865 179011 462931 179014
rect 510654 179012 510660 179014
rect 510724 179012 510730 179076
rect 583520 179060 584960 179150
rect 349889 178938 349955 178941
rect 414289 178938 414355 178941
rect 349889 178936 414355 178938
rect 349889 178880 349894 178936
rect 349950 178880 414294 178936
rect 414350 178880 414355 178936
rect 349889 178878 414355 178880
rect 349889 178875 349955 178878
rect 414289 178875 414355 178878
rect 457805 178938 457871 178941
rect 503662 178938 503668 178940
rect 457805 178936 503668 178938
rect 457805 178880 457810 178936
rect 457866 178880 503668 178936
rect 457805 178878 503668 178880
rect 457805 178875 457871 178878
rect 503662 178876 503668 178878
rect 503732 178876 503738 178940
rect 296110 178802 296116 178804
rect 279956 178742 296116 178802
rect 296110 178740 296116 178742
rect 296180 178740 296186 178804
rect 456793 178802 456859 178805
rect 503110 178802 503116 178804
rect 456793 178800 503116 178802
rect 456793 178744 456798 178800
rect 456854 178744 503116 178800
rect 456793 178742 503116 178744
rect 456793 178739 456859 178742
rect 503110 178740 503116 178742
rect 503180 178740 503186 178804
rect 283281 178666 283347 178669
rect 355174 178666 355180 178668
rect 283281 178664 355180 178666
rect 283281 178608 283286 178664
rect 283342 178608 355180 178664
rect 283281 178606 355180 178608
rect 283281 178603 283347 178606
rect 355174 178604 355180 178606
rect 355244 178604 355250 178668
rect 130377 178258 130443 178261
rect 327574 178258 327580 178260
rect 130377 178256 240212 178258
rect 130377 178200 130382 178256
rect 130438 178200 240212 178256
rect 130377 178198 240212 178200
rect 279956 178198 327580 178258
rect 130377 178195 130443 178198
rect 327574 178196 327580 178198
rect 327644 178196 327650 178260
rect 57789 177986 57855 177989
rect 358169 177986 358235 177989
rect 372797 177986 372863 177989
rect 57789 177984 60076 177986
rect 57789 177928 57794 177984
rect 57850 177928 60076 177984
rect 57789 177926 60076 177928
rect 358169 177984 372863 177986
rect 358169 177928 358174 177984
rect 358230 177928 372802 177984
rect 372858 177928 372863 177984
rect 358169 177926 372863 177928
rect 57789 177923 57855 177926
rect 358169 177923 358235 177926
rect 372797 177923 372863 177926
rect 490189 177986 490255 177989
rect 522982 177986 522988 177988
rect 490189 177984 522988 177986
rect 490189 177928 490194 177984
rect 490250 177928 522988 177984
rect 490189 177926 522988 177928
rect 490189 177923 490255 177926
rect 522982 177924 522988 177926
rect 523052 177924 523058 177988
rect 336089 177850 336155 177853
rect 371785 177850 371851 177853
rect 336089 177848 371851 177850
rect 336089 177792 336094 177848
rect 336150 177792 371790 177848
rect 371846 177792 371851 177848
rect 336089 177790 371851 177792
rect 336089 177787 336155 177790
rect 371785 177787 371851 177790
rect 471973 177850 472039 177853
rect 512126 177850 512132 177852
rect 471973 177848 512132 177850
rect 471973 177792 471978 177848
rect 472034 177792 512132 177848
rect 471973 177790 512132 177792
rect 471973 177787 472039 177790
rect 512126 177788 512132 177790
rect 512196 177788 512202 177852
rect 217174 177714 217180 177716
rect 124844 177654 217180 177714
rect 217174 177652 217180 177654
rect 217244 177652 217250 177716
rect 302734 177714 302740 177716
rect 279956 177654 302740 177714
rect 302734 177652 302740 177654
rect 302804 177652 302810 177716
rect 355501 177714 355567 177717
rect 374821 177714 374887 177717
rect 355501 177712 374887 177714
rect 355501 177656 355506 177712
rect 355562 177656 374826 177712
rect 374882 177656 374887 177712
rect 355501 177654 374887 177656
rect 355501 177651 355567 177654
rect 374821 177651 374887 177654
rect 487153 177714 487219 177717
rect 521694 177714 521700 177716
rect 487153 177712 521700 177714
rect 487153 177656 487158 177712
rect 487214 177656 521700 177712
rect 487153 177654 521700 177656
rect 487153 177651 487219 177654
rect 521694 177652 521700 177654
rect 521764 177652 521770 177716
rect 349797 177578 349863 177581
rect 413277 177578 413343 177581
rect 349797 177576 413343 177578
rect 349797 177520 349802 177576
rect 349858 177520 413282 177576
rect 413338 177520 413343 177576
rect 349797 177518 413343 177520
rect 349797 177515 349863 177518
rect 413277 177515 413343 177518
rect 481081 177578 481147 177581
rect 515070 177578 515076 177580
rect 481081 177576 515076 177578
rect 481081 177520 481086 177576
rect 481142 177520 515076 177576
rect 481081 177518 515076 177520
rect 481081 177515 481147 177518
rect 515070 177516 515076 177518
rect 515140 177516 515146 177580
rect 493225 177442 493291 177445
rect 525926 177442 525932 177444
rect 493225 177440 525932 177442
rect 493225 177384 493230 177440
rect 493286 177384 525932 177440
rect 493225 177382 525932 177384
rect 493225 177379 493291 177382
rect 525926 177380 525932 177382
rect 525996 177380 526002 177444
rect 438577 177306 438643 177309
rect 499798 177306 499804 177308
rect 438577 177304 499804 177306
rect 438577 177248 438582 177304
rect 438638 177248 499804 177304
rect 438577 177246 499804 177248
rect 438577 177243 438643 177246
rect 499798 177244 499804 177246
rect 499868 177244 499874 177308
rect 186957 177170 187023 177173
rect 294638 177170 294644 177172
rect 186957 177168 240212 177170
rect 186957 177112 186962 177168
rect 187018 177112 240212 177168
rect 186957 177110 240212 177112
rect 279956 177110 294644 177170
rect 186957 177107 187023 177110
rect 294638 177108 294644 177110
rect 294708 177108 294714 177172
rect 133137 176762 133203 176765
rect 134517 176762 134583 176765
rect 133137 176760 134583 176762
rect 133137 176704 133142 176760
rect 133198 176704 134522 176760
rect 134578 176704 134583 176760
rect 133137 176702 134583 176704
rect 133137 176699 133203 176702
rect 134517 176699 134583 176702
rect 299974 176626 299980 176628
rect 279956 176566 299980 176626
rect 299974 176564 299980 176566
rect 300044 176564 300050 176628
rect 341609 176626 341675 176629
rect 391013 176626 391079 176629
rect 341609 176624 391079 176626
rect 341609 176568 341614 176624
rect 341670 176568 391018 176624
rect 391074 176568 391079 176624
rect 341609 176566 391079 176568
rect 341609 176563 341675 176566
rect 391013 176563 391079 176566
rect 420361 176626 420427 176629
rect 510470 176626 510476 176628
rect 420361 176624 510476 176626
rect 420361 176568 420366 176624
rect 420422 176568 510476 176624
rect 420361 176566 510476 176568
rect 420361 176563 420427 176566
rect 510470 176564 510476 176566
rect 510540 176564 510546 176628
rect 57513 176490 57579 176493
rect 57646 176490 57652 176492
rect 57513 176488 57652 176490
rect 57513 176432 57518 176488
rect 57574 176432 57652 176488
rect 57513 176430 57652 176432
rect 57513 176427 57579 176430
rect 57646 176428 57652 176430
rect 57716 176428 57722 176492
rect 437565 176490 437631 176493
rect 527214 176490 527220 176492
rect 437565 176488 527220 176490
rect 437565 176432 437570 176488
rect 437626 176432 527220 176488
rect 437565 176430 527220 176432
rect 437565 176427 437631 176430
rect 527214 176428 527220 176430
rect 527284 176428 527290 176492
rect 433517 176354 433583 176357
rect 508998 176354 509004 176356
rect 433517 176352 509004 176354
rect 433517 176296 433522 176352
rect 433578 176296 509004 176352
rect 433517 176294 509004 176296
rect 433517 176291 433583 176294
rect 508998 176292 509004 176294
rect 509068 176292 509074 176356
rect 216622 176218 216628 176220
rect 124814 176158 216628 176218
rect -960 175796 480 176036
rect 57830 176020 57836 176084
rect 57900 176082 57906 176084
rect 57900 176022 60076 176082
rect 124814 176052 124874 176158
rect 216622 176156 216628 176158
rect 216692 176156 216698 176220
rect 435541 176218 435607 176221
rect 510838 176218 510844 176220
rect 435541 176216 510844 176218
rect 435541 176160 435546 176216
rect 435602 176160 510844 176216
rect 435541 176158 510844 176160
rect 435541 176155 435607 176158
rect 510838 176156 510844 176158
rect 510908 176156 510914 176220
rect 142797 176082 142863 176085
rect 289486 176082 289492 176084
rect 142797 176080 240212 176082
rect 142797 176024 142802 176080
rect 142858 176024 240212 176080
rect 142797 176022 240212 176024
rect 279956 176022 289492 176082
rect 57900 176020 57906 176022
rect 142797 176019 142863 176022
rect 289486 176020 289492 176022
rect 289556 176020 289562 176084
rect 424409 176082 424475 176085
rect 499614 176082 499620 176084
rect 424409 176080 499620 176082
rect 424409 176024 424414 176080
rect 424470 176024 499620 176080
rect 424409 176022 499620 176024
rect 424409 176019 424475 176022
rect 499614 176020 499620 176022
rect 499684 176020 499690 176084
rect 356646 175538 356652 175540
rect 279956 175478 356652 175538
rect 356646 175476 356652 175478
rect 356716 175476 356722 175540
rect 315389 175402 315455 175405
rect 313230 175400 315455 175402
rect 313230 175344 315394 175400
rect 315450 175344 315455 175400
rect 313230 175342 315455 175344
rect 57421 175266 57487 175269
rect 57830 175266 57836 175268
rect 57421 175264 57836 175266
rect 57421 175208 57426 175264
rect 57482 175208 57836 175264
rect 57421 175206 57836 175208
rect 57421 175203 57487 175206
rect 57830 175204 57836 175206
rect 57900 175204 57906 175268
rect 310513 175266 310579 175269
rect 313230 175266 313290 175342
rect 315389 175339 315455 175342
rect 310513 175264 313290 175266
rect 310513 175208 310518 175264
rect 310574 175208 313290 175264
rect 310513 175206 313290 175208
rect 418337 175266 418403 175269
rect 506790 175266 506796 175268
rect 418337 175264 506796 175266
rect 418337 175208 418342 175264
rect 418398 175208 506796 175264
rect 418337 175206 506796 175208
rect 310513 175203 310579 175206
rect 418337 175203 418403 175206
rect 506790 175204 506796 175206
rect 506860 175204 506866 175268
rect 422385 175130 422451 175133
rect 500166 175130 500172 175132
rect 422385 175128 500172 175130
rect 422385 175072 422390 175128
rect 422446 175072 500172 175128
rect 422385 175070 500172 175072
rect 422385 175067 422451 175070
rect 500166 175068 500172 175070
rect 500236 175068 500242 175132
rect 57881 174994 57947 174997
rect 58617 174994 58683 174997
rect 57881 174992 58683 174994
rect 57881 174936 57886 174992
rect 57942 174936 58622 174992
rect 58678 174936 58683 174992
rect 57881 174934 58683 174936
rect 57881 174931 57947 174934
rect 58617 174931 58683 174934
rect 138657 174994 138723 174997
rect 288934 174994 288940 174996
rect 138657 174992 240212 174994
rect 138657 174936 138662 174992
rect 138718 174936 240212 174992
rect 138657 174934 240212 174936
rect 279956 174934 288940 174994
rect 138657 174931 138723 174934
rect 288934 174932 288940 174934
rect 289004 174932 289010 174996
rect 425421 174994 425487 174997
rect 501638 174994 501644 174996
rect 425421 174992 501644 174994
rect 425421 174936 425426 174992
rect 425482 174936 501644 174992
rect 425421 174934 501644 174936
rect 425421 174931 425487 174934
rect 501638 174932 501644 174934
rect 501708 174932 501714 174996
rect 428457 174858 428523 174861
rect 503846 174858 503852 174860
rect 428457 174856 503852 174858
rect 428457 174800 428462 174856
rect 428518 174800 503852 174856
rect 428457 174798 503852 174800
rect 428457 174795 428523 174798
rect 503846 174796 503852 174798
rect 503916 174796 503922 174860
rect 432505 174722 432571 174725
rect 507894 174722 507900 174724
rect 432505 174720 507900 174722
rect 432505 174664 432510 174720
rect 432566 174664 507900 174720
rect 432505 174662 507900 174664
rect 432505 174659 432571 174662
rect 507894 174660 507900 174662
rect 507964 174660 507970 174724
rect 289486 174524 289492 174588
rect 289556 174586 289562 174588
rect 357934 174586 357940 174588
rect 289556 174526 357940 174586
rect 289556 174524 289562 174526
rect 357934 174524 357940 174526
rect 358004 174524 358010 174588
rect 431493 174586 431559 174589
rect 506606 174586 506612 174588
rect 431493 174584 506612 174586
rect 431493 174528 431498 174584
rect 431554 174528 506612 174584
rect 431493 174526 506612 174528
rect 431493 174523 431559 174526
rect 506606 174524 506612 174526
rect 506676 174524 506682 174588
rect 226190 174450 226196 174452
rect 124844 174390 226196 174450
rect 226190 174388 226196 174390
rect 226260 174388 226266 174452
rect 305494 174450 305500 174452
rect 279956 174390 305500 174450
rect 305494 174388 305500 174390
rect 305564 174388 305570 174452
rect 439589 174450 439655 174453
rect 514702 174450 514708 174452
rect 439589 174448 514708 174450
rect 439589 174392 439594 174448
rect 439650 174392 514708 174448
rect 439589 174390 514708 174392
rect 439589 174387 439655 174390
rect 514702 174388 514708 174390
rect 514772 174388 514778 174452
rect 57462 174116 57468 174180
rect 57532 174178 57538 174180
rect 57532 174118 60076 174178
rect 57532 174116 57538 174118
rect 238017 173906 238083 173909
rect 238661 173906 238727 173909
rect 295926 173906 295932 173908
rect 238017 173904 240212 173906
rect 238017 173848 238022 173904
rect 238078 173848 238666 173904
rect 238722 173848 240212 173904
rect 238017 173846 240212 173848
rect 279956 173846 295932 173906
rect 238017 173843 238083 173846
rect 238661 173843 238727 173846
rect 295926 173844 295932 173846
rect 295996 173844 296002 173908
rect 304206 173362 304212 173364
rect 279956 173302 304212 173362
rect 304206 173300 304212 173302
rect 304276 173300 304282 173364
rect 48221 173226 48287 173229
rect 57237 173226 57303 173229
rect 48221 173224 57303 173226
rect 48221 173168 48226 173224
rect 48282 173168 57242 173224
rect 57298 173168 57303 173224
rect 48221 173166 57303 173168
rect 48221 173163 48287 173166
rect 57237 173163 57303 173166
rect 355869 173226 355935 173229
rect 365713 173226 365779 173229
rect 355869 173224 365779 173226
rect 355869 173168 355874 173224
rect 355930 173168 365718 173224
rect 365774 173168 365779 173224
rect 355869 173166 365779 173168
rect 355869 173163 355935 173166
rect 365713 173163 365779 173166
rect 219934 172818 219940 172820
rect 124844 172758 219940 172818
rect 219934 172756 219940 172758
rect 220004 172756 220010 172820
rect 235901 172818 235967 172821
rect 322054 172818 322060 172820
rect 235901 172816 240212 172818
rect 235901 172760 235906 172816
rect 235962 172760 240212 172816
rect 235901 172758 240212 172760
rect 279956 172758 322060 172818
rect 235901 172755 235967 172758
rect 322054 172756 322060 172758
rect 322124 172756 322130 172820
rect 358721 172546 358787 172549
rect 407113 172546 407179 172549
rect 358721 172544 407179 172546
rect 358721 172488 358726 172544
rect 358782 172488 407118 172544
rect 407174 172488 407179 172544
rect 358721 172486 407179 172488
rect 358721 172483 358787 172486
rect 407113 172483 407179 172486
rect 57278 172348 57284 172412
rect 57348 172410 57354 172412
rect 57881 172410 57947 172413
rect 57348 172408 57947 172410
rect 57348 172352 57886 172408
rect 57942 172352 57947 172408
rect 57348 172350 57947 172352
rect 57348 172348 57354 172350
rect 57881 172347 57947 172350
rect 57646 172212 57652 172276
rect 57716 172274 57722 172276
rect 323526 172274 323532 172276
rect 57716 172214 60076 172274
rect 279956 172214 323532 172274
rect 57716 172212 57722 172214
rect 323526 172212 323532 172214
rect 323596 172212 323602 172276
rect 231158 171668 231164 171732
rect 231228 171730 231234 171732
rect 311014 171730 311020 171732
rect 231228 171670 240212 171730
rect 279956 171670 311020 171730
rect 231228 171668 231234 171670
rect 311014 171668 311020 171670
rect 311084 171668 311090 171732
rect 360009 171730 360075 171733
rect 402973 171730 403039 171733
rect 360009 171728 403039 171730
rect 360009 171672 360014 171728
rect 360070 171672 402978 171728
rect 403034 171672 403039 171728
rect 360009 171670 403039 171672
rect 360009 171667 360075 171670
rect 402973 171667 403039 171670
rect 220854 171186 220860 171188
rect 124844 171126 220860 171186
rect 220854 171124 220860 171126
rect 220924 171124 220930 171188
rect 291694 171186 291700 171188
rect 279956 171126 291700 171186
rect 291694 171124 291700 171126
rect 291764 171124 291770 171188
rect 228214 170580 228220 170644
rect 228284 170642 228290 170644
rect 282821 170642 282887 170645
rect 228284 170582 240212 170642
rect 279956 170640 282887 170642
rect 279956 170584 282826 170640
rect 282882 170584 282887 170640
rect 279956 170582 282887 170584
rect 228284 170580 228290 170582
rect 282821 170579 282887 170582
rect 57830 170308 57836 170372
rect 57900 170370 57906 170372
rect 57900 170310 60076 170370
rect 57900 170308 57906 170310
rect 291561 170098 291627 170101
rect 279956 170096 291627 170098
rect 279956 170040 291566 170096
rect 291622 170040 291627 170096
rect 279956 170038 291627 170040
rect 291561 170035 291627 170038
rect 282126 169764 282132 169828
rect 282196 169826 282202 169828
rect 283281 169826 283347 169829
rect 282196 169824 283347 169826
rect 282196 169768 283286 169824
rect 283342 169768 283347 169824
rect 282196 169766 283347 169768
rect 282196 169764 282202 169766
rect 283281 169763 283347 169766
rect 308397 169826 308463 169829
rect 310421 169826 310487 169829
rect 308397 169824 310487 169826
rect 308397 169768 308402 169824
rect 308458 169768 310426 169824
rect 310482 169768 310487 169824
rect 308397 169766 310487 169768
rect 308397 169763 308463 169766
rect 310421 169763 310487 169766
rect 223798 169690 223804 169692
rect 124814 169630 223804 169690
rect 124814 169524 124874 169630
rect 223798 169628 223804 169630
rect 223868 169628 223874 169692
rect 134374 169492 134380 169556
rect 134444 169554 134450 169556
rect 290590 169554 290596 169556
rect 134444 169494 240212 169554
rect 279956 169494 290596 169554
rect 134444 169492 134450 169494
rect 290590 169492 290596 169494
rect 290660 169492 290666 169556
rect 360326 169084 360332 169148
rect 360396 169146 360402 169148
rect 394969 169146 395035 169149
rect 360396 169144 395035 169146
rect 360396 169088 394974 169144
rect 395030 169088 395035 169144
rect 360396 169086 395035 169088
rect 360396 169084 360402 169086
rect 394969 169083 395035 169086
rect 291326 169010 291332 169012
rect 279956 168950 291332 169010
rect 291326 168948 291332 168950
rect 291396 168948 291402 169012
rect 364977 169010 365043 169013
rect 529197 169010 529263 169013
rect 364977 169008 529263 169010
rect 364977 168952 364982 169008
rect 365038 168952 529202 169008
rect 529258 168952 529263 169008
rect 364977 168950 529263 168952
rect 364977 168947 365043 168950
rect 529197 168947 529263 168950
rect 59854 168676 59860 168740
rect 59924 168738 59930 168740
rect 60273 168738 60339 168741
rect 59924 168736 60339 168738
rect 59924 168680 60278 168736
rect 60334 168680 60339 168736
rect 59924 168678 60339 168680
rect 59924 168676 59930 168678
rect 60273 168675 60339 168678
rect 60222 168404 60228 168468
rect 60292 168404 60298 168468
rect 235390 168404 235396 168468
rect 235460 168466 235466 168468
rect 282821 168466 282887 168469
rect 235460 168406 240212 168466
rect 279956 168464 282887 168466
rect 279956 168408 282826 168464
rect 282882 168408 282887 168464
rect 279956 168406 282887 168408
rect 235460 168404 235466 168406
rect 282821 168403 282887 168406
rect 223614 167922 223620 167924
rect 124844 167862 223620 167922
rect 223614 167860 223620 167862
rect 223684 167860 223690 167924
rect 282637 167922 282703 167925
rect 279956 167920 282703 167922
rect 279956 167864 282642 167920
rect 282698 167864 282703 167920
rect 279956 167862 282703 167864
rect 282637 167859 282703 167862
rect 304349 167650 304415 167653
rect 369853 167650 369919 167653
rect 304349 167648 369919 167650
rect 304349 167592 304354 167648
rect 304410 167592 369858 167648
rect 369914 167592 369919 167648
rect 304349 167590 369919 167592
rect 304349 167587 304415 167590
rect 369853 167587 369919 167590
rect 213126 167316 213132 167380
rect 213196 167378 213202 167380
rect 282453 167378 282519 167381
rect 213196 167318 240212 167378
rect 279956 167376 282519 167378
rect 279956 167320 282458 167376
rect 282514 167320 282519 167376
rect 279956 167318 282519 167320
rect 213196 167316 213202 167318
rect 282453 167315 282519 167318
rect 58566 167044 58572 167108
rect 58636 167106 58642 167108
rect 59261 167106 59327 167109
rect 58636 167104 59327 167106
rect 58636 167048 59266 167104
rect 59322 167048 59327 167104
rect 58636 167046 59327 167048
rect 58636 167044 58642 167046
rect 59261 167043 59327 167046
rect 134517 167106 134583 167109
rect 136541 167106 136607 167109
rect 134517 167104 136607 167106
rect 134517 167048 134522 167104
rect 134578 167048 136546 167104
rect 136602 167048 136607 167104
rect 134517 167046 136607 167048
rect 134517 167043 134583 167046
rect 136541 167043 136607 167046
rect 282821 166834 282887 166837
rect 279956 166832 282887 166834
rect 279956 166776 282826 166832
rect 282882 166776 282887 166832
rect 279956 166774 282887 166776
rect 282821 166771 282887 166774
rect 60038 166500 60044 166564
rect 60108 166500 60114 166564
rect 214782 166364 214788 166428
rect 214852 166426 214858 166428
rect 214852 166366 238770 166426
rect 214852 166364 214858 166366
rect 229870 166290 229876 166292
rect 124844 166230 229876 166290
rect 229870 166228 229876 166230
rect 229940 166228 229946 166292
rect 238710 166290 238770 166366
rect 283046 166290 283052 166292
rect 238710 166230 240212 166290
rect 279956 166230 283052 166290
rect 283046 166228 283052 166230
rect 283116 166228 283122 166292
rect 363597 166290 363663 166293
rect 524321 166290 524387 166293
rect 363597 166288 524387 166290
rect 363597 166232 363602 166288
rect 363658 166232 524326 166288
rect 524382 166232 524387 166288
rect 363597 166230 524387 166232
rect 363597 166227 363663 166230
rect 524321 166227 524387 166230
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 284334 165746 284340 165748
rect 279956 165686 284340 165746
rect 284334 165684 284340 165686
rect 284404 165684 284410 165748
rect 583520 165732 584960 165822
rect 230974 165140 230980 165204
rect 231044 165202 231050 165204
rect 282821 165202 282887 165205
rect 231044 165142 240212 165202
rect 279956 165200 282887 165202
rect 279956 165144 282826 165200
rect 282882 165144 282887 165200
rect 279956 165142 282887 165144
rect 231044 165140 231050 165142
rect 282821 165139 282887 165142
rect 60590 164596 60596 164660
rect 60660 164596 60666 164660
rect 222694 164658 222700 164660
rect 124844 164598 222700 164658
rect 222694 164596 222700 164598
rect 222764 164596 222770 164660
rect 282862 164658 282868 164660
rect 279956 164598 282868 164658
rect 282862 164596 282868 164598
rect 282932 164596 282938 164660
rect 224309 164114 224375 164117
rect 298134 164114 298140 164116
rect 224309 164112 240212 164114
rect 224309 164056 224314 164112
rect 224370 164056 240212 164112
rect 224309 164054 240212 164056
rect 279956 164054 298140 164114
rect 224309 164051 224375 164054
rect 298134 164052 298140 164054
rect 298204 164052 298210 164116
rect 282821 163570 282887 163573
rect 279956 163568 282887 163570
rect 279956 163512 282826 163568
rect 282882 163512 282887 163568
rect 279956 163510 282887 163512
rect 282821 163507 282887 163510
rect 224902 163162 224908 163164
rect 124814 163102 224908 163162
rect 124814 162996 124874 163102
rect 224902 163100 224908 163102
rect 224972 163100 224978 163164
rect -960 162890 480 162980
rect 137134 162964 137140 163028
rect 137204 163026 137210 163028
rect 282637 163026 282703 163029
rect 137204 162966 240212 163026
rect 279956 163024 282703 163026
rect 279956 162968 282642 163024
rect 282698 162968 282703 163024
rect 279956 162966 282703 162968
rect 137204 162964 137210 162966
rect 282637 162963 282703 162966
rect 3417 162890 3483 162893
rect 308397 162890 308463 162893
rect -960 162888 3483 162890
rect -960 162832 3422 162888
rect 3478 162832 3483 162888
rect -960 162830 3483 162832
rect -960 162740 480 162830
rect 3417 162827 3483 162830
rect 306330 162888 308463 162890
rect 306330 162832 308402 162888
rect 308458 162832 308463 162888
rect 306330 162830 308463 162832
rect 58893 162754 58959 162757
rect 59118 162754 59124 162756
rect 58893 162752 59124 162754
rect 58893 162696 58898 162752
rect 58954 162696 59124 162752
rect 58893 162694 59124 162696
rect 58893 162691 58959 162694
rect 59118 162692 59124 162694
rect 59188 162692 59194 162756
rect 59302 162692 59308 162756
rect 59372 162754 59378 162756
rect 303981 162754 304047 162757
rect 306330 162754 306390 162830
rect 308397 162827 308463 162830
rect 59372 162694 60076 162754
rect 303981 162752 306390 162754
rect 303981 162696 303986 162752
rect 304042 162696 306390 162752
rect 303981 162694 306390 162696
rect 59372 162692 59378 162694
rect 303981 162691 304047 162694
rect 282821 162482 282887 162485
rect 279956 162480 282887 162482
rect 279956 162424 282826 162480
rect 282882 162424 282887 162480
rect 279956 162422 282887 162424
rect 282821 162419 282887 162422
rect 293350 162012 293356 162076
rect 293420 162074 293426 162076
rect 580206 162074 580212 162076
rect 293420 162014 580212 162074
rect 293420 162012 293426 162014
rect 580206 162012 580212 162014
rect 580276 162012 580282 162076
rect 238334 161876 238340 161940
rect 238404 161938 238410 161940
rect 282637 161938 282703 161941
rect 238404 161878 240212 161938
rect 279956 161936 282703 161938
rect 279956 161880 282642 161936
rect 282698 161880 282703 161936
rect 279956 161878 282703 161880
rect 238404 161876 238410 161878
rect 282637 161875 282703 161878
rect 230054 161394 230060 161396
rect 124844 161334 230060 161394
rect 230054 161332 230060 161334
rect 230124 161332 230130 161396
rect 282821 161394 282887 161397
rect 279956 161392 282887 161394
rect 279956 161336 282826 161392
rect 282882 161336 282887 161392
rect 279956 161334 282887 161336
rect 282821 161331 282887 161334
rect 58750 160788 58756 160852
rect 58820 160850 58826 160852
rect 58820 160790 60076 160850
rect 58820 160788 58826 160790
rect 237966 160788 237972 160852
rect 238036 160850 238042 160852
rect 303981 160850 304047 160853
rect 238036 160790 240212 160850
rect 279956 160848 304047 160850
rect 279956 160792 303986 160848
rect 304042 160792 304047 160848
rect 279956 160790 304047 160792
rect 238036 160788 238042 160790
rect 303981 160787 304047 160790
rect 291837 160714 291903 160717
rect 580441 160714 580507 160717
rect 291837 160712 580507 160714
rect 291837 160656 291842 160712
rect 291898 160656 580446 160712
rect 580502 160656 580507 160712
rect 291837 160654 580507 160656
rect 291837 160651 291903 160654
rect 580441 160651 580507 160654
rect 298737 160306 298803 160309
rect 279956 160304 298803 160306
rect 279956 160248 298742 160304
rect 298798 160248 298803 160304
rect 279956 160246 298803 160248
rect 298737 160243 298803 160246
rect 58750 160108 58756 160172
rect 58820 160170 58826 160172
rect 58985 160170 59051 160173
rect 58820 160168 59051 160170
rect 58820 160112 58990 160168
rect 59046 160112 59051 160168
rect 58820 160110 59051 160112
rect 58820 160108 58826 160110
rect 58985 160107 59051 160110
rect 136633 160170 136699 160173
rect 143441 160170 143507 160173
rect 136633 160168 143507 160170
rect 136633 160112 136638 160168
rect 136694 160112 143446 160168
rect 143502 160112 143507 160168
rect 136633 160110 143507 160112
rect 136633 160107 136699 160110
rect 143441 160107 143507 160110
rect 235574 159762 235580 159764
rect 124844 159702 235580 159762
rect 235574 159700 235580 159702
rect 235644 159700 235650 159764
rect 238150 159700 238156 159764
rect 238220 159762 238226 159764
rect 500217 159762 500283 159765
rect 238220 159702 240212 159762
rect 279956 159760 500283 159762
rect 279956 159704 500222 159760
rect 500278 159704 500283 159760
rect 279956 159702 500283 159704
rect 238220 159700 238226 159702
rect 500217 159699 500283 159702
rect 508078 159218 508084 159220
rect 279956 159158 508084 159218
rect 508078 159156 508084 159158
rect 508148 159156 508154 159220
rect 57646 158884 57652 158948
rect 57716 158946 57722 158948
rect 57716 158886 60076 158946
rect 57716 158884 57722 158886
rect 57697 158810 57763 158813
rect 57830 158810 57836 158812
rect 57697 158808 57836 158810
rect 57697 158752 57702 158808
rect 57758 158752 57836 158808
rect 57697 158750 57836 158752
rect 57697 158747 57763 158750
rect 57830 158748 57836 158750
rect 57900 158748 57906 158812
rect 238477 158674 238543 158677
rect 547873 158674 547939 158677
rect 238477 158672 240212 158674
rect 238477 158616 238482 158672
rect 238538 158616 240212 158672
rect 238477 158614 240212 158616
rect 279956 158672 547939 158674
rect 279956 158616 547878 158672
rect 547934 158616 547939 158672
rect 279956 158614 547939 158616
rect 238477 158611 238543 158614
rect 547873 158611 547939 158614
rect 235758 158130 235764 158132
rect 124844 158070 235764 158130
rect 235758 158068 235764 158070
rect 235828 158068 235834 158132
rect 558126 158130 558132 158132
rect 279956 158070 558132 158130
rect 558126 158068 558132 158070
rect 558196 158068 558202 158132
rect 178677 157586 178743 157589
rect 555366 157586 555372 157588
rect 178677 157584 240212 157586
rect 178677 157528 178682 157584
rect 178738 157528 240212 157584
rect 178677 157526 240212 157528
rect 279956 157526 555372 157586
rect 178677 157523 178743 157526
rect 555366 157524 555372 157526
rect 555436 157524 555442 157588
rect 58566 156980 58572 157044
rect 58636 157042 58642 157044
rect 551134 157042 551140 157044
rect 58636 156982 60076 157042
rect 279956 156982 551140 157042
rect 58636 156980 58642 156982
rect 551134 156980 551140 156982
rect 551204 156980 551210 157044
rect 58382 156572 58388 156636
rect 58452 156634 58458 156636
rect 58801 156634 58867 156637
rect 58452 156632 58867 156634
rect 58452 156576 58806 156632
rect 58862 156576 58867 156632
rect 58452 156574 58867 156576
rect 58452 156572 58458 156574
rect 58801 156571 58867 156574
rect 235206 156572 235212 156636
rect 235276 156634 235282 156636
rect 235717 156634 235783 156637
rect 235276 156632 235783 156634
rect 235276 156576 235722 156632
rect 235778 156576 235783 156632
rect 235276 156574 235783 156576
rect 235276 156572 235282 156574
rect 235717 156571 235783 156574
rect 235390 156498 235396 156500
rect 124844 156438 235396 156498
rect 235390 156436 235396 156438
rect 235460 156436 235466 156500
rect 238385 156498 238451 156501
rect 548374 156498 548380 156500
rect 238385 156496 240212 156498
rect 238385 156440 238390 156496
rect 238446 156440 240212 156496
rect 238385 156438 240212 156440
rect 279956 156438 548380 156498
rect 238385 156435 238451 156438
rect 548374 156436 548380 156438
rect 548444 156436 548450 156500
rect 58566 155892 58572 155956
rect 58636 155954 58642 155956
rect 59077 155954 59143 155957
rect 58636 155952 59143 155954
rect 58636 155896 59082 155952
rect 59138 155896 59143 155952
rect 58636 155894 59143 155896
rect 58636 155892 58642 155894
rect 59077 155891 59143 155894
rect 143441 155954 143507 155957
rect 147673 155954 147739 155957
rect 143441 155952 147739 155954
rect 143441 155896 143446 155952
rect 143502 155896 147678 155952
rect 147734 155896 147739 155952
rect 143441 155894 147739 155896
rect 143441 155891 143507 155894
rect 147673 155891 147739 155894
rect 234654 155892 234660 155956
rect 234724 155954 234730 155956
rect 235809 155954 235875 155957
rect 547086 155954 547092 155956
rect 234724 155952 235875 155954
rect 234724 155896 235814 155952
rect 235870 155896 235875 155952
rect 234724 155894 235875 155896
rect 279956 155894 547092 155954
rect 234724 155892 234730 155894
rect 235809 155891 235875 155894
rect 547086 155892 547092 155894
rect 547156 155892 547162 155956
rect 237373 155410 237439 155413
rect 544326 155410 544332 155412
rect 237373 155408 240212 155410
rect 237373 155352 237378 155408
rect 237434 155352 240212 155408
rect 237373 155350 240212 155352
rect 279956 155350 544332 155410
rect 237373 155347 237439 155350
rect 544326 155348 544332 155350
rect 544396 155348 544402 155412
rect 58934 155076 58940 155140
rect 59004 155138 59010 155140
rect 59004 155078 60076 155138
rect 59004 155076 59010 155078
rect 235206 154866 235212 154868
rect 124844 154806 235212 154866
rect 235206 154804 235212 154806
rect 235276 154804 235282 154868
rect 293350 154866 293356 154868
rect 279956 154806 293356 154866
rect 293350 154804 293356 154806
rect 293420 154804 293426 154868
rect 57462 154396 57468 154460
rect 57532 154458 57538 154460
rect 57605 154458 57671 154461
rect 57532 154456 57671 154458
rect 57532 154400 57610 154456
rect 57666 154400 57671 154456
rect 57532 154398 57671 154400
rect 57532 154396 57538 154398
rect 57605 154395 57671 154398
rect 237373 154322 237439 154325
rect 542854 154322 542860 154324
rect 237373 154320 240212 154322
rect 237373 154264 237378 154320
rect 237434 154264 240212 154320
rect 237373 154262 240212 154264
rect 279956 154262 542860 154322
rect 237373 154259 237439 154262
rect 542854 154260 542860 154262
rect 542924 154260 542930 154324
rect 508446 153778 508452 153780
rect 279956 153718 508452 153778
rect 508446 153716 508452 153718
rect 508516 153716 508522 153780
rect 147673 153370 147739 153373
rect 147673 153368 238770 153370
rect 147673 153312 147678 153368
rect 147734 153312 238770 153368
rect 147673 153310 238770 153312
rect 147673 153307 147739 153310
rect 57278 153172 57284 153236
rect 57348 153234 57354 153236
rect 235349 153234 235415 153237
rect 57348 153174 60076 153234
rect 124844 153232 235415 153234
rect 124844 153176 235354 153232
rect 235410 153176 235415 153232
rect 124844 153174 235415 153176
rect 238710 153234 238770 153310
rect 291837 153234 291903 153237
rect 238710 153174 240212 153234
rect 279956 153232 291903 153234
rect 279956 153176 291842 153232
rect 291898 153176 291903 153232
rect 279956 153174 291903 153176
rect 57348 153172 57354 153174
rect 235349 153171 235415 153174
rect 291837 153171 291903 153174
rect 334750 152690 334756 152692
rect 279956 152630 334756 152690
rect 334750 152628 334756 152630
rect 334820 152628 334826 152692
rect 580165 152690 580231 152693
rect 583520 152690 584960 152780
rect 580165 152688 584960 152690
rect 580165 152632 580170 152688
rect 580226 152632 584960 152688
rect 580165 152630 584960 152632
rect 580165 152627 580231 152630
rect 583520 152540 584960 152630
rect 237281 152146 237347 152149
rect 306414 152146 306420 152148
rect 237281 152144 240212 152146
rect 237281 152088 237286 152144
rect 237342 152088 240212 152144
rect 237281 152086 240212 152088
rect 279956 152086 306420 152146
rect 237281 152083 237347 152086
rect 306414 152084 306420 152086
rect 306484 152084 306490 152148
rect 238150 151602 238156 151604
rect 124844 151542 238156 151602
rect 238150 151540 238156 151542
rect 238220 151540 238226 151604
rect 313774 151602 313780 151604
rect 279956 151542 313780 151602
rect 313774 151540 313780 151542
rect 313844 151540 313850 151604
rect 58750 151268 58756 151332
rect 58820 151330 58826 151332
rect 58820 151270 60076 151330
rect 58820 151268 58826 151270
rect 339125 151194 339191 151197
rect 375833 151194 375899 151197
rect 339125 151192 375899 151194
rect 339125 151136 339130 151192
rect 339186 151136 375838 151192
rect 375894 151136 375899 151192
rect 339125 151134 375899 151136
rect 339125 151131 339191 151134
rect 375833 151131 375899 151134
rect 231761 151058 231827 151061
rect 231761 151056 240212 151058
rect 231761 151000 231766 151056
rect 231822 151000 240212 151056
rect 231761 150998 240212 151000
rect 279956 150998 296730 151058
rect 231761 150995 231827 150998
rect 296670 150922 296730 150998
rect 306414 150996 306420 151060
rect 306484 151058 306490 151060
rect 580206 151058 580212 151060
rect 306484 150998 580212 151058
rect 306484 150996 306490 150998
rect 580206 150996 580212 150998
rect 580276 150996 580282 151060
rect 306966 150922 306972 150924
rect 296670 150862 306972 150922
rect 306966 150860 306972 150862
rect 307036 150860 307042 150924
rect 298686 150514 298692 150516
rect 279956 150454 298692 150514
rect 298686 150452 298692 150454
rect 298756 150452 298762 150516
rect 233141 150106 233207 150109
rect 233141 150104 239690 150106
rect 233141 150048 233146 150104
rect 233202 150048 239690 150104
rect 233141 150046 239690 150048
rect 233141 150043 233207 150046
rect 239630 150038 239690 150046
rect 239630 149978 240212 150038
rect 237966 149970 237972 149972
rect -960 149834 480 149924
rect 124844 149910 237972 149970
rect 237966 149908 237972 149910
rect 238036 149908 238042 149972
rect 54334 149834 54340 149836
rect -960 149774 54340 149834
rect -960 149684 480 149774
rect 54334 149772 54340 149774
rect 54404 149772 54410 149836
rect 59118 149364 59124 149428
rect 59188 149426 59194 149428
rect 59188 149366 60076 149426
rect 59188 149364 59194 149366
rect 227621 149018 227687 149021
rect 227621 149016 239690 149018
rect 227621 148960 227626 149016
rect 227682 148960 239690 149016
rect 227621 148958 239690 148960
rect 227621 148955 227687 148958
rect 239630 148950 239690 148958
rect 239630 148890 240212 148950
rect 323577 148610 323643 148613
rect 383009 148610 383075 148613
rect 323577 148608 383075 148610
rect 323577 148552 323582 148608
rect 323638 148552 383014 148608
rect 383070 148552 383075 148608
rect 323577 148550 383075 148552
rect 323577 148547 323643 148550
rect 383009 148547 383075 148550
rect 318057 148474 318123 148477
rect 379421 148474 379487 148477
rect 318057 148472 379487 148474
rect 318057 148416 318062 148472
rect 318118 148416 379426 148472
rect 379482 148416 379487 148472
rect 318057 148414 379487 148416
rect 318057 148411 318123 148414
rect 379421 148411 379487 148414
rect 127566 148338 127572 148340
rect 124844 148278 127572 148338
rect 127566 148276 127572 148278
rect 127636 148276 127642 148340
rect 316677 148338 316743 148341
rect 378225 148338 378291 148341
rect 316677 148336 378291 148338
rect 316677 148280 316682 148336
rect 316738 148280 378230 148336
rect 378286 148280 378291 148336
rect 316677 148278 378291 148280
rect 316677 148275 316743 148278
rect 378225 148275 378291 148278
rect 239857 147862 239923 147865
rect 239857 147860 240212 147862
rect 239857 147804 239862 147860
rect 239918 147804 240212 147860
rect 239857 147802 240212 147804
rect 239857 147799 239923 147802
rect 352557 147658 352623 147661
rect 353937 147658 354003 147661
rect 352557 147656 364350 147658
rect 352557 147600 352562 147656
rect 352618 147600 353942 147656
rect 353998 147600 364350 147656
rect 352557 147598 364350 147600
rect 352557 147595 352623 147598
rect 353937 147595 354003 147598
rect 58566 147460 58572 147524
rect 58636 147522 58642 147524
rect 58636 147462 60076 147522
rect 58636 147460 58642 147462
rect 297357 147386 297423 147389
rect 355961 147386 356027 147389
rect 297357 147384 356027 147386
rect 297357 147328 297362 147384
rect 297418 147328 355966 147384
rect 356022 147328 356027 147384
rect 297357 147326 356027 147328
rect 297357 147323 297423 147326
rect 355961 147323 356027 147326
rect 364290 147250 364350 147598
rect 400949 147250 401015 147253
rect 364290 147248 401015 147250
rect 364290 147192 400954 147248
rect 401010 147192 401015 147248
rect 364290 147190 401015 147192
rect 400949 147187 401015 147190
rect 350073 147114 350139 147117
rect 357525 147114 357591 147117
rect 367461 147114 367527 147117
rect 350073 147112 367527 147114
rect 350073 147056 350078 147112
rect 350134 147056 357530 147112
rect 357586 147056 367466 147112
rect 367522 147056 367527 147112
rect 350073 147054 367527 147056
rect 350073 147051 350139 147054
rect 357525 147051 357591 147054
rect 367461 147051 367527 147054
rect 295609 146978 295675 146981
rect 295977 146978 296043 146981
rect 358721 146978 358787 146981
rect 295609 146976 358787 146978
rect 295609 146920 295614 146976
rect 295670 146920 295982 146976
rect 296038 146920 358726 146976
rect 358782 146920 358787 146976
rect 295609 146918 358787 146920
rect 295609 146915 295675 146918
rect 295977 146915 296043 146918
rect 358721 146915 358787 146918
rect 239857 146774 239923 146777
rect 239857 146772 240212 146774
rect 239857 146716 239862 146772
rect 239918 146716 240212 146772
rect 239857 146714 240212 146716
rect 239857 146711 239923 146714
rect 127750 146706 127756 146708
rect 124844 146646 127756 146706
rect 127750 146644 127756 146646
rect 127820 146644 127826 146708
rect 355317 146706 355383 146709
rect 399753 146706 399819 146709
rect 355317 146704 399819 146706
rect 355317 146648 355322 146704
rect 355378 146648 399758 146704
rect 399814 146648 399819 146704
rect 355317 146646 399819 146648
rect 355317 146643 355383 146646
rect 399753 146643 399819 146646
rect 352741 146570 352807 146573
rect 357341 146570 357407 146573
rect 402145 146570 402211 146573
rect 352741 146568 402211 146570
rect 352741 146512 352746 146568
rect 352802 146512 357346 146568
rect 357402 146512 402150 146568
rect 402206 146512 402211 146568
rect 352741 146510 402211 146512
rect 352741 146507 352807 146510
rect 357341 146507 357407 146510
rect 402145 146507 402211 146510
rect 352925 146434 352991 146437
rect 402973 146434 403039 146437
rect 352925 146432 403039 146434
rect 352925 146376 352930 146432
rect 352986 146376 402978 146432
rect 403034 146376 403039 146432
rect 352925 146374 403039 146376
rect 352925 146371 352991 146374
rect 402973 146371 403039 146374
rect 239806 145624 239812 145688
rect 239876 145686 239882 145688
rect 239876 145626 240212 145686
rect 239876 145624 239882 145626
rect 58382 145556 58388 145620
rect 58452 145618 58458 145620
rect 58452 145558 60076 145618
rect 58452 145556 58458 145558
rect 127934 145074 127940 145076
rect 124844 145014 127940 145074
rect 127934 145012 127940 145014
rect 128004 145012 128010 145076
rect 57145 144802 57211 144805
rect 57646 144802 57652 144804
rect 57145 144800 57652 144802
rect 57145 144744 57150 144800
rect 57206 144744 57652 144800
rect 57145 144742 57652 144744
rect 57145 144739 57211 144742
rect 57646 144740 57652 144742
rect 57716 144740 57722 144804
rect 407205 144802 407271 144805
rect 407614 144802 407620 144804
rect 393270 144800 407620 144802
rect 393270 144744 407210 144800
rect 407266 144744 407620 144800
rect 393270 144742 407620 144744
rect 239622 144536 239628 144600
rect 239692 144598 239698 144600
rect 239692 144538 240212 144598
rect 239692 144536 239698 144538
rect 358537 144530 358603 144533
rect 393270 144530 393330 144742
rect 407205 144739 407271 144742
rect 407614 144740 407620 144742
rect 407684 144740 407690 144804
rect 358537 144528 393330 144530
rect 358537 144472 358542 144528
rect 358598 144472 393330 144528
rect 358537 144470 393330 144472
rect 358537 144467 358603 144470
rect 355501 144394 355567 144397
rect 396165 144394 396231 144397
rect 355501 144392 396231 144394
rect 355501 144336 355506 144392
rect 355562 144336 396170 144392
rect 396226 144336 396231 144392
rect 355501 144334 396231 144336
rect 355501 144331 355567 144334
rect 396165 144331 396231 144334
rect 57830 143652 57836 143716
rect 57900 143714 57906 143716
rect 57900 143654 60076 143714
rect 57900 143652 57906 143654
rect 239806 143448 239812 143512
rect 239876 143510 239882 143512
rect 239876 143450 240212 143510
rect 239876 143448 239882 143450
rect 57789 143442 57855 143445
rect 59997 143442 60063 143445
rect 128118 143442 128124 143444
rect 57789 143440 60063 143442
rect 57789 143384 57794 143440
rect 57850 143384 60002 143440
rect 60058 143384 60063 143440
rect 57789 143382 60063 143384
rect 124844 143382 128124 143442
rect 57789 143379 57855 143382
rect 59997 143379 60063 143382
rect 128118 143380 128124 143382
rect 128188 143380 128194 143444
rect 302918 142700 302924 142764
rect 302988 142762 302994 142764
rect 302988 142702 357450 142762
rect 302988 142700 302994 142702
rect 239622 142360 239628 142424
rect 239692 142422 239698 142424
rect 239692 142362 240212 142422
rect 239692 142360 239698 142362
rect 357390 142082 357450 142702
rect 357390 142022 360210 142082
rect 57646 141748 57652 141812
rect 57716 141810 57722 141812
rect 127709 141810 127775 141813
rect 57716 141750 60076 141810
rect 124844 141808 127775 141810
rect 124844 141752 127714 141808
rect 127770 141752 127775 141808
rect 124844 141750 127775 141752
rect 57716 141748 57722 141750
rect 127709 141747 127775 141750
rect 238518 141340 238524 141404
rect 238588 141402 238594 141404
rect 238588 141342 239690 141402
rect 238588 141340 238594 141342
rect 239630 141334 239690 141342
rect 327758 141340 327764 141404
rect 327828 141402 327834 141404
rect 357382 141402 357388 141404
rect 327828 141342 357388 141402
rect 327828 141340 327834 141342
rect 357382 141340 357388 141342
rect 357452 141340 357458 141404
rect 360150 141372 360210 142022
rect 239630 141274 240212 141334
rect 235717 140314 235783 140317
rect 235717 140312 239690 140314
rect 235717 140256 235722 140312
rect 235778 140256 239690 140312
rect 235717 140254 239690 140256
rect 235717 140251 235783 140254
rect 239630 140246 239690 140254
rect 346894 140252 346900 140316
rect 346964 140314 346970 140316
rect 346964 140254 360180 140314
rect 346964 140252 346970 140254
rect 239630 140186 240212 140246
rect 127617 140178 127683 140181
rect 124844 140176 127683 140178
rect 124844 140120 127622 140176
rect 127678 140120 127683 140176
rect 124844 140118 127683 140120
rect 127617 140115 127683 140118
rect 290774 139980 290780 140044
rect 290844 140042 290850 140044
rect 357566 140042 357572 140044
rect 290844 139982 357572 140042
rect 290844 139980 290850 139982
rect 357566 139980 357572 139982
rect 357636 139980 357642 140044
rect 57462 139844 57468 139908
rect 57532 139906 57538 139908
rect 57532 139846 60076 139906
rect 57532 139844 57538 139846
rect 580206 139300 580212 139364
rect 580276 139362 580282 139364
rect 583520 139362 584960 139452
rect 580276 139302 584960 139362
rect 580276 139300 580282 139302
rect 345606 139164 345612 139228
rect 345676 139226 345682 139228
rect 407205 139226 407271 139229
rect 345676 139166 360180 139226
rect 404892 139224 407271 139226
rect 404892 139168 407210 139224
rect 407266 139168 407271 139224
rect 583520 139212 584960 139302
rect 404892 139166 407271 139168
rect 345676 139164 345682 139166
rect 407205 139163 407271 139166
rect 239630 139098 240212 139158
rect 238477 139090 238543 139093
rect 239630 139090 239690 139098
rect 238477 139088 239690 139090
rect 238477 139032 238482 139088
rect 238538 139032 239690 139088
rect 238477 139030 239690 139032
rect 238477 139027 238543 139030
rect 59854 138484 59860 138548
rect 59924 138546 59930 138548
rect 127893 138546 127959 138549
rect 59924 138486 60106 138546
rect 124844 138544 127959 138546
rect 124844 138488 127898 138544
rect 127954 138488 127959 138544
rect 124844 138486 127959 138488
rect 59924 138484 59930 138486
rect 60046 137972 60106 138486
rect 127893 138483 127959 138486
rect 357382 138076 357388 138140
rect 357452 138138 357458 138140
rect 357452 138078 360180 138138
rect 357452 138076 357458 138078
rect 239814 138010 240212 138070
rect 238385 138002 238451 138005
rect 239814 138002 239874 138010
rect 238385 138000 239874 138002
rect 238385 137944 238390 138000
rect 238446 137944 239874 138000
rect 238385 137942 239874 137944
rect 238385 137939 238451 137942
rect 338614 137260 338620 137324
rect 338684 137322 338690 137324
rect 357382 137322 357388 137324
rect 338684 137262 357388 137322
rect 338684 137260 338690 137262
rect 357382 137260 357388 137262
rect 357452 137260 357458 137324
rect 357566 136988 357572 137052
rect 357636 137050 357642 137052
rect 357636 136990 360180 137050
rect 357636 136988 357642 136990
rect 239630 136922 240212 136982
rect 235257 136914 235323 136917
rect 124844 136912 235323 136914
rect -960 136778 480 136868
rect 124844 136856 235262 136912
rect 235318 136856 235323 136912
rect 124844 136854 235323 136856
rect 235257 136851 235323 136854
rect 238334 136852 238340 136916
rect 238404 136914 238410 136916
rect 239630 136914 239690 136922
rect 238404 136854 239690 136914
rect 238404 136852 238410 136854
rect 3366 136778 3372 136780
rect -960 136718 3372 136778
rect -960 136628 480 136718
rect 3366 136716 3372 136718
rect 3436 136716 3442 136780
rect 59670 136036 59676 136100
rect 59740 136098 59746 136100
rect 59740 136038 60076 136098
rect 59740 136036 59746 136038
rect 313958 135900 313964 135964
rect 314028 135962 314034 135964
rect 314028 135902 360180 135962
rect 314028 135900 314034 135902
rect 239630 135834 240212 135894
rect 238518 135764 238524 135828
rect 238588 135826 238594 135828
rect 239630 135826 239690 135834
rect 238588 135766 239690 135826
rect 238588 135764 238594 135766
rect 128077 135282 128143 135285
rect 124844 135280 128143 135282
rect 124844 135224 128082 135280
rect 128138 135224 128143 135280
rect 124844 135222 128143 135224
rect 128077 135219 128143 135222
rect 280061 135148 280127 135149
rect 280061 135144 280108 135148
rect 280172 135146 280178 135148
rect 280061 135088 280066 135144
rect 280061 135084 280108 135088
rect 280172 135086 280218 135146
rect 280172 135084 280178 135086
rect 280061 135083 280127 135084
rect 357382 134812 357388 134876
rect 357452 134874 357458 134876
rect 357452 134814 360180 134874
rect 357452 134812 357458 134814
rect 239622 134744 239628 134808
rect 239692 134806 239698 134808
rect 239692 134746 240212 134806
rect 239692 134744 239698 134746
rect 280061 134738 280127 134741
rect 281942 134738 281948 134740
rect 280061 134736 281948 134738
rect 280061 134680 280066 134736
rect 280122 134680 281948 134736
rect 280061 134678 281948 134680
rect 280061 134675 280127 134678
rect 281942 134676 281948 134678
rect 282012 134676 282018 134740
rect 334566 134404 334572 134468
rect 334636 134466 334642 134468
rect 357382 134466 357388 134468
rect 334636 134406 357388 134466
rect 334636 134404 334642 134406
rect 357382 134404 357388 134406
rect 357452 134404 357458 134468
rect 57789 134194 57855 134197
rect 57789 134192 60076 134194
rect 57789 134136 57794 134192
rect 57850 134136 60076 134192
rect 57789 134134 60076 134136
rect 57789 134131 57855 134134
rect 300158 133724 300164 133788
rect 300228 133786 300234 133788
rect 300228 133726 360180 133786
rect 300228 133724 300234 133726
rect 239630 133658 240212 133718
rect 128261 133650 128327 133653
rect 124844 133648 128327 133650
rect 124844 133592 128266 133648
rect 128322 133592 128327 133648
rect 124844 133590 128327 133592
rect 128261 133587 128327 133590
rect 239438 133588 239444 133652
rect 239508 133650 239514 133652
rect 239630 133650 239690 133658
rect 239508 133590 239690 133650
rect 239508 133588 239514 133590
rect 357382 132636 357388 132700
rect 357452 132698 357458 132700
rect 357452 132638 360180 132698
rect 357452 132636 357458 132638
rect 239806 132568 239812 132632
rect 239876 132630 239882 132632
rect 239876 132570 240212 132630
rect 239876 132568 239882 132570
rect 60089 132562 60155 132565
rect 60046 132560 60155 132562
rect 60046 132504 60094 132560
rect 60150 132504 60155 132560
rect 60046 132499 60155 132504
rect 60046 132260 60106 132499
rect 127433 132018 127499 132021
rect 124844 132016 127499 132018
rect 124844 131960 127438 132016
rect 127494 131960 127499 132016
rect 124844 131958 127499 131960
rect 127433 131955 127499 131958
rect 291878 131548 291884 131612
rect 291948 131610 291954 131612
rect 291948 131550 360180 131610
rect 291948 131548 291954 131550
rect 291377 131202 291443 131205
rect 291510 131202 291516 131204
rect 291377 131200 291516 131202
rect 291377 131144 291382 131200
rect 291438 131144 291516 131200
rect 291377 131142 291516 131144
rect 291377 131139 291443 131142
rect 291510 131140 291516 131142
rect 291580 131140 291586 131204
rect 60181 130930 60247 130933
rect 60181 130928 60290 130930
rect 60181 130872 60186 130928
rect 60242 130872 60290 130928
rect 60181 130867 60290 130872
rect 60230 130356 60290 130867
rect 319294 130460 319300 130524
rect 319364 130522 319370 130524
rect 319364 130462 360180 130522
rect 319364 130460 319370 130462
rect 127341 130386 127407 130389
rect 124844 130384 127407 130386
rect 124844 130328 127346 130384
rect 127402 130328 127407 130384
rect 124844 130326 127407 130328
rect 127341 130323 127407 130326
rect 298870 129372 298876 129436
rect 298940 129434 298946 129436
rect 298940 129374 360180 129434
rect 298940 129372 298946 129374
rect 127801 128754 127867 128757
rect 124844 128752 127867 128754
rect 124844 128696 127806 128752
rect 127862 128696 127867 128752
rect 124844 128694 127867 128696
rect 127801 128691 127867 128694
rect 57329 128482 57395 128485
rect 57329 128480 60076 128482
rect 57329 128424 57334 128480
rect 57390 128424 60076 128480
rect 57329 128422 60076 128424
rect 57329 128419 57395 128422
rect 342846 128284 342852 128348
rect 342916 128346 342922 128348
rect 342916 128286 360180 128346
rect 342916 128284 342922 128286
rect 407757 128074 407823 128077
rect 404892 128072 407823 128074
rect 404892 128016 407762 128072
rect 407818 128016 407823 128072
rect 404892 128014 407823 128016
rect 407757 128011 407823 128014
rect 349654 127196 349660 127260
rect 349724 127258 349730 127260
rect 349724 127198 360180 127258
rect 349724 127196 349730 127198
rect 127249 127122 127315 127125
rect 124844 127120 127315 127122
rect 124844 127064 127254 127120
rect 127310 127064 127315 127120
rect 124844 127062 127315 127064
rect 127249 127059 127315 127062
rect 59169 126578 59235 126581
rect 59169 126576 60076 126578
rect 59169 126520 59174 126576
rect 59230 126520 60076 126576
rect 59169 126518 60076 126520
rect 59169 126515 59235 126518
rect 335854 126108 335860 126172
rect 335924 126170 335930 126172
rect 335924 126110 360180 126170
rect 335924 126108 335930 126110
rect 583520 125884 584960 126124
rect 128077 125490 128143 125493
rect 124844 125488 128143 125490
rect 124844 125432 128082 125488
rect 128138 125432 128143 125488
rect 124844 125430 128143 125432
rect 128077 125427 128143 125430
rect 293953 125490 294019 125493
rect 294270 125490 294276 125492
rect 293953 125488 294276 125490
rect 293953 125432 293958 125488
rect 294014 125432 294276 125488
rect 293953 125430 294276 125432
rect 293953 125427 294019 125430
rect 294270 125428 294276 125430
rect 294340 125428 294346 125492
rect 294822 125020 294828 125084
rect 294892 125082 294898 125084
rect 294892 125022 360180 125082
rect 294892 125020 294898 125022
rect 56501 124674 56567 124677
rect 56501 124672 60076 124674
rect 56501 124616 56506 124672
rect 56562 124616 60076 124672
rect 56501 124614 60076 124616
rect 56501 124611 56567 124614
rect 307150 123932 307156 123996
rect 307220 123994 307226 123996
rect 307220 123934 360180 123994
rect 307220 123932 307226 123934
rect 237782 123858 237788 123860
rect -960 123572 480 123812
rect 124844 123798 237788 123858
rect 237782 123796 237788 123798
rect 237852 123796 237858 123860
rect 238017 123586 238083 123589
rect 238334 123586 238340 123588
rect 238017 123584 238340 123586
rect 238017 123528 238022 123584
rect 238078 123528 238340 123584
rect 238017 123526 238340 123528
rect 238017 123523 238083 123526
rect 238334 123524 238340 123526
rect 238404 123524 238410 123588
rect 353886 122844 353892 122908
rect 353956 122906 353962 122908
rect 353956 122846 360180 122906
rect 353956 122844 353962 122846
rect 57237 122770 57303 122773
rect 57237 122768 60076 122770
rect 57237 122712 57242 122768
rect 57298 122712 60076 122768
rect 57237 122710 60076 122712
rect 57237 122707 57303 122710
rect 309726 121756 309732 121820
rect 309796 121818 309802 121820
rect 309796 121758 360180 121818
rect 309796 121756 309802 121758
rect 57237 121546 57303 121549
rect 57830 121546 57836 121548
rect 57237 121544 57836 121546
rect 57237 121488 57242 121544
rect 57298 121488 57836 121544
rect 57237 121486 57836 121488
rect 57237 121483 57303 121486
rect 57830 121484 57836 121486
rect 57900 121484 57906 121548
rect 127566 121348 127572 121412
rect 127636 121410 127642 121412
rect 287278 121410 287284 121412
rect 127636 121350 287284 121410
rect 127636 121348 127642 121350
rect 287278 121348 287284 121350
rect 287348 121348 287354 121412
rect 128118 121212 128124 121276
rect 128188 121274 128194 121276
rect 287462 121274 287468 121276
rect 128188 121214 287468 121274
rect 128188 121212 128194 121214
rect 287462 121212 287468 121214
rect 287532 121212 287538 121276
rect 127709 121138 127775 121141
rect 285765 121138 285831 121141
rect 127709 121136 285831 121138
rect 127709 121080 127714 121136
rect 127770 121080 285770 121136
rect 285826 121080 285831 121136
rect 127709 121078 285831 121080
rect 127709 121075 127775 121078
rect 285765 121075 285831 121078
rect 127893 121002 127959 121005
rect 284385 121002 284451 121005
rect 127893 121000 284451 121002
rect 127893 120944 127898 121000
rect 127954 120944 284390 121000
rect 284446 120944 284451 121000
rect 127893 120942 284451 120944
rect 127893 120939 127959 120942
rect 284385 120939 284451 120942
rect 127341 120866 127407 120869
rect 235809 120866 235875 120869
rect 127341 120864 235875 120866
rect 127341 120808 127346 120864
rect 127402 120808 235814 120864
rect 235870 120808 235875 120864
rect 127341 120806 235875 120808
rect 127341 120803 127407 120806
rect 235809 120803 235875 120806
rect 296110 120804 296116 120868
rect 296180 120866 296186 120868
rect 357566 120866 357572 120868
rect 296180 120806 357572 120866
rect 296180 120804 296186 120806
rect 357566 120804 357572 120806
rect 357636 120804 357642 120868
rect 129089 120730 129155 120733
rect 235901 120730 235967 120733
rect 129089 120728 235967 120730
rect 129089 120672 129094 120728
rect 129150 120672 235906 120728
rect 235962 120672 235967 120728
rect 129089 120670 235967 120672
rect 129089 120667 129155 120670
rect 235901 120667 235967 120670
rect 351126 120668 351132 120732
rect 351196 120730 351202 120732
rect 351196 120670 360180 120730
rect 351196 120668 351202 120670
rect 50429 120594 50495 120597
rect 86309 120594 86375 120597
rect 50429 120592 86375 120594
rect 50429 120536 50434 120592
rect 50490 120536 86314 120592
rect 86370 120536 86375 120592
rect 50429 120534 86375 120536
rect 50429 120531 50495 120534
rect 86309 120531 86375 120534
rect 234654 120532 234660 120596
rect 234724 120594 234730 120596
rect 235717 120594 235783 120597
rect 295425 120594 295491 120597
rect 234724 120592 235783 120594
rect 234724 120536 235722 120592
rect 235778 120536 235783 120592
rect 234724 120534 235783 120536
rect 234724 120532 234730 120534
rect 235717 120531 235783 120534
rect 237238 120592 295491 120594
rect 237238 120536 295430 120592
rect 295486 120536 295491 120592
rect 237238 120534 295491 120536
rect 49417 120458 49483 120461
rect 82813 120458 82879 120461
rect 49417 120456 82879 120458
rect 49417 120400 49422 120456
rect 49478 120400 82818 120456
rect 82874 120400 82879 120456
rect 49417 120398 82879 120400
rect 49417 120395 49483 120398
rect 82813 120395 82879 120398
rect 235349 120458 235415 120461
rect 237238 120458 237298 120534
rect 295425 120531 295491 120534
rect 292614 120458 292620 120460
rect 235349 120456 237298 120458
rect 235349 120400 235354 120456
rect 235410 120400 237298 120456
rect 235349 120398 237298 120400
rect 237422 120398 292620 120458
rect 235349 120395 235415 120398
rect 55121 120322 55187 120325
rect 88057 120322 88123 120325
rect 55121 120320 88123 120322
rect 55121 120264 55126 120320
rect 55182 120264 88062 120320
rect 88118 120264 88123 120320
rect 55121 120262 88123 120264
rect 55121 120259 55187 120262
rect 88057 120259 88123 120262
rect 235809 120322 235875 120325
rect 237281 120322 237347 120325
rect 235809 120320 237347 120322
rect 235809 120264 235814 120320
rect 235870 120264 237286 120320
rect 237342 120264 237347 120320
rect 235809 120262 237347 120264
rect 235809 120259 235875 120262
rect 237281 120259 237347 120262
rect 235206 120124 235212 120188
rect 235276 120186 235282 120188
rect 237422 120186 237482 120398
rect 292614 120396 292620 120398
rect 292684 120396 292690 120460
rect 237557 120322 237623 120325
rect 279969 120322 280035 120325
rect 237557 120320 280035 120322
rect 237557 120264 237562 120320
rect 237618 120264 279974 120320
rect 280030 120264 280035 120320
rect 237557 120262 280035 120264
rect 237557 120259 237623 120262
rect 279969 120259 280035 120262
rect 235276 120126 237482 120186
rect 279693 120186 279759 120189
rect 281993 120186 282059 120189
rect 279693 120184 282059 120186
rect 279693 120128 279698 120184
rect 279754 120128 281998 120184
rect 282054 120128 282059 120184
rect 279693 120126 282059 120128
rect 235276 120124 235282 120126
rect 279693 120123 279759 120126
rect 281993 120123 282059 120126
rect 47853 120050 47919 120053
rect 70393 120050 70459 120053
rect 127617 120050 127683 120053
rect 47853 120048 127683 120050
rect 47853 119992 47858 120048
rect 47914 119992 70398 120048
rect 70454 119992 127622 120048
rect 127678 119992 127683 120048
rect 47853 119990 127683 119992
rect 47853 119987 47919 119990
rect 70393 119987 70459 119990
rect 127617 119987 127683 119990
rect 238293 120050 238359 120053
rect 238518 120050 238524 120052
rect 238293 120048 238524 120050
rect 238293 119992 238298 120048
rect 238354 119992 238524 120048
rect 238293 119990 238524 119992
rect 238293 119987 238359 119990
rect 238518 119988 238524 119990
rect 238588 119988 238594 120052
rect 284293 120050 284359 120053
rect 284518 120050 284524 120052
rect 284293 120048 284524 120050
rect 284293 119992 284298 120048
rect 284354 119992 284524 120048
rect 284293 119990 284524 119992
rect 284293 119987 284359 119990
rect 284518 119988 284524 119990
rect 284588 119988 284594 120052
rect 53097 119914 53163 119917
rect 74073 119914 74139 119917
rect 53097 119912 74139 119914
rect 53097 119856 53102 119912
rect 53158 119856 74078 119912
rect 74134 119856 74139 119912
rect 53097 119854 74139 119856
rect 53097 119851 53163 119854
rect 74073 119851 74139 119854
rect 93301 119914 93367 119917
rect 126329 119914 126395 119917
rect 93301 119912 126395 119914
rect 93301 119856 93306 119912
rect 93362 119856 126334 119912
rect 126390 119856 126395 119912
rect 93301 119854 126395 119856
rect 93301 119851 93367 119854
rect 126329 119851 126395 119854
rect 127750 119852 127756 119916
rect 127820 119914 127826 119916
rect 287094 119914 287100 119916
rect 127820 119854 287100 119914
rect 127820 119852 127826 119854
rect 287094 119852 287100 119854
rect 287164 119852 287170 119916
rect 95049 119778 95115 119781
rect 126973 119778 127039 119781
rect 95049 119776 127039 119778
rect 95049 119720 95054 119776
rect 95110 119720 126978 119776
rect 127034 119720 127039 119776
rect 95049 119718 127039 119720
rect 95049 119715 95115 119718
rect 126973 119715 127039 119718
rect 127934 119716 127940 119780
rect 128004 119778 128010 119780
rect 285622 119778 285628 119780
rect 128004 119718 285628 119778
rect 128004 119716 128010 119718
rect 285622 119716 285628 119718
rect 285692 119716 285698 119780
rect 96797 119642 96863 119645
rect 127801 119642 127867 119645
rect 96797 119640 127867 119642
rect 96797 119584 96802 119640
rect 96858 119584 127806 119640
rect 127862 119584 127867 119640
rect 96797 119582 127867 119584
rect 96797 119579 96863 119582
rect 127801 119579 127867 119582
rect 127985 119642 128051 119645
rect 283005 119642 283071 119645
rect 127985 119640 283071 119642
rect 127985 119584 127990 119640
rect 128046 119584 283010 119640
rect 283066 119584 283071 119640
rect 127985 119582 283071 119584
rect 127985 119579 128051 119582
rect 283005 119579 283071 119582
rect 355174 119580 355180 119644
rect 355244 119642 355250 119644
rect 355244 119582 360180 119642
rect 355244 119580 355250 119582
rect 127433 119506 127499 119509
rect 238569 119506 238635 119509
rect 294270 119506 294276 119508
rect 127433 119504 238635 119506
rect 127433 119448 127438 119504
rect 127494 119448 238574 119504
rect 238630 119448 238635 119504
rect 127433 119446 238635 119448
rect 127433 119443 127499 119446
rect 238569 119443 238635 119446
rect 238710 119446 294276 119506
rect 48630 119308 48636 119372
rect 48700 119370 48706 119372
rect 127525 119370 127591 119373
rect 48700 119368 127591 119370
rect 48700 119312 127530 119368
rect 127586 119312 127591 119368
rect 48700 119310 127591 119312
rect 48700 119308 48706 119310
rect 127525 119307 127591 119310
rect 235758 119308 235764 119372
rect 235828 119370 235834 119372
rect 235828 119310 236194 119370
rect 235828 119308 235834 119310
rect 128261 119234 128327 119237
rect 235901 119234 235967 119237
rect 128261 119232 235967 119234
rect 128261 119176 128266 119232
rect 128322 119176 235906 119232
rect 235962 119176 235967 119232
rect 128261 119174 235967 119176
rect 236134 119234 236194 119310
rect 238150 119308 238156 119372
rect 238220 119370 238226 119372
rect 238710 119370 238770 119446
rect 294270 119444 294276 119446
rect 294340 119444 294346 119508
rect 238220 119310 238770 119370
rect 238845 119370 238911 119373
rect 291285 119370 291351 119373
rect 238845 119368 291351 119370
rect 238845 119312 238850 119368
rect 238906 119312 291290 119368
rect 291346 119312 291351 119368
rect 238845 119310 291351 119312
rect 238220 119308 238226 119310
rect 238845 119307 238911 119310
rect 291285 119307 291351 119310
rect 327574 119308 327580 119372
rect 327644 119370 327650 119372
rect 357382 119370 357388 119372
rect 327644 119310 357388 119370
rect 327644 119308 327650 119310
rect 357382 119308 357388 119310
rect 357452 119308 357458 119372
rect 291510 119234 291516 119236
rect 236134 119174 291516 119234
rect 128261 119171 128327 119174
rect 235901 119171 235967 119174
rect 291510 119172 291516 119174
rect 291580 119172 291586 119236
rect 127617 119098 127683 119101
rect 287145 119098 287211 119101
rect 127617 119096 287211 119098
rect 127617 119040 127622 119096
rect 127678 119040 287150 119096
rect 287206 119040 287211 119096
rect 127617 119038 287211 119040
rect 127617 119035 127683 119038
rect 287145 119035 287211 119038
rect 127249 118962 127315 118965
rect 235809 118962 235875 118965
rect 127249 118960 235875 118962
rect 127249 118904 127254 118960
rect 127310 118904 235814 118960
rect 235870 118904 235875 118960
rect 127249 118902 235875 118904
rect 127249 118899 127315 118902
rect 235809 118899 235875 118902
rect 235257 118826 235323 118829
rect 238845 118826 238911 118829
rect 235257 118824 238911 118826
rect 235257 118768 235262 118824
rect 235318 118768 238850 118824
rect 238906 118768 238911 118824
rect 235257 118766 238911 118768
rect 235257 118763 235323 118766
rect 238845 118763 238911 118766
rect 291561 118826 291627 118829
rect 291878 118826 291884 118828
rect 291561 118824 291884 118826
rect 291561 118768 291566 118824
rect 291622 118768 291884 118824
rect 291561 118766 291884 118768
rect 291561 118763 291627 118766
rect 291878 118764 291884 118766
rect 291948 118764 291954 118828
rect 238661 118690 238727 118693
rect 358077 118690 358143 118693
rect 238661 118688 358143 118690
rect 238661 118632 238666 118688
rect 238722 118632 358082 118688
rect 358138 118632 358143 118688
rect 238661 118630 358143 118632
rect 238661 118627 238727 118630
rect 358077 118627 358143 118630
rect 235574 118492 235580 118556
rect 235644 118554 235650 118556
rect 294454 118554 294460 118556
rect 235644 118494 294460 118554
rect 235644 118492 235650 118494
rect 294454 118492 294460 118494
rect 294524 118492 294530 118556
rect 357566 118492 357572 118556
rect 357636 118554 357642 118556
rect 357636 118494 360180 118554
rect 357636 118492 357642 118494
rect 237966 118356 237972 118420
rect 238036 118418 238042 118420
rect 271781 118418 271847 118421
rect 238036 118416 271847 118418
rect 238036 118360 271786 118416
rect 271842 118360 271847 118416
rect 238036 118358 271847 118360
rect 238036 118356 238042 118358
rect 271781 118355 271847 118358
rect 247769 118282 247835 118285
rect 282085 118282 282151 118285
rect 247769 118280 282151 118282
rect 247769 118224 247774 118280
rect 247830 118224 282090 118280
rect 282146 118224 282151 118280
rect 247769 118222 282151 118224
rect 247769 118219 247835 118222
rect 282085 118219 282151 118222
rect 21817 118146 21883 118149
rect 121453 118146 121519 118149
rect 21817 118144 121519 118146
rect 21817 118088 21822 118144
rect 21878 118088 121458 118144
rect 121514 118088 121519 118144
rect 21817 118086 121519 118088
rect 21817 118083 21883 118086
rect 121453 118083 121519 118086
rect 122281 118146 122347 118149
rect 277669 118146 277735 118149
rect 122281 118144 277735 118146
rect 122281 118088 122286 118144
rect 122342 118088 277674 118144
rect 277730 118088 277735 118144
rect 122281 118086 277735 118088
rect 122281 118083 122347 118086
rect 277669 118083 277735 118086
rect 279417 118146 279483 118149
rect 291837 118146 291903 118149
rect 279417 118144 291903 118146
rect 279417 118088 279422 118144
rect 279478 118088 291842 118144
rect 291898 118088 291903 118144
rect 279417 118086 291903 118088
rect 279417 118083 279483 118086
rect 291837 118083 291903 118086
rect 44265 118010 44331 118013
rect 251357 118010 251423 118013
rect 44265 118008 251423 118010
rect 44265 117952 44270 118008
rect 44326 117952 251362 118008
rect 251418 117952 251423 118008
rect 44265 117950 251423 117952
rect 44265 117947 44331 117950
rect 251357 117947 251423 117950
rect 265341 118010 265407 118013
rect 286225 118010 286291 118013
rect 265341 118008 286291 118010
rect 265341 117952 265346 118008
rect 265402 117952 286230 118008
rect 286286 117952 286291 118008
rect 265341 117950 286291 117952
rect 265341 117947 265407 117950
rect 286225 117947 286291 117950
rect 37181 117874 37247 117877
rect 237373 117874 237439 117877
rect 37181 117872 237439 117874
rect 37181 117816 37186 117872
rect 37242 117816 237378 117872
rect 237434 117816 237439 117872
rect 37181 117814 237439 117816
rect 37181 117811 37247 117814
rect 237373 117811 237439 117814
rect 33593 117738 33659 117741
rect 237465 117738 237531 117741
rect 33593 117736 237531 117738
rect 33593 117680 33598 117736
rect 33654 117680 237470 117736
rect 237526 117680 237531 117736
rect 33593 117678 237531 117680
rect 33593 117675 33659 117678
rect 237465 117675 237531 117678
rect 261753 117738 261819 117741
rect 280245 117738 280311 117741
rect 261753 117736 280311 117738
rect 261753 117680 261758 117736
rect 261814 117680 280250 117736
rect 280306 117680 280311 117736
rect 261753 117678 280311 117680
rect 261753 117675 261819 117678
rect 280245 117675 280311 117678
rect 40677 117602 40743 117605
rect 247033 117602 247099 117605
rect 40677 117600 247099 117602
rect 40677 117544 40682 117600
rect 40738 117544 247038 117600
rect 247094 117544 247099 117600
rect 40677 117542 247099 117544
rect 40677 117539 40743 117542
rect 247033 117539 247099 117542
rect 30097 117466 30163 117469
rect 237557 117466 237623 117469
rect 30097 117464 237623 117466
rect 30097 117408 30102 117464
rect 30158 117408 237562 117464
rect 237618 117408 237623 117464
rect 30097 117406 237623 117408
rect 30097 117403 30163 117406
rect 237557 117403 237623 117406
rect 237782 117404 237788 117468
rect 237852 117466 237858 117468
rect 264973 117466 265039 117469
rect 237852 117464 265039 117466
rect 237852 117408 264978 117464
rect 265034 117408 265039 117464
rect 237852 117406 265039 117408
rect 237852 117404 237858 117406
rect 264973 117403 265039 117406
rect 357382 117404 357388 117468
rect 357452 117466 357458 117468
rect 357452 117406 360180 117466
rect 357452 117404 357458 117406
rect 26509 117330 26575 117333
rect 234613 117330 234679 117333
rect 26509 117328 234679 117330
rect 26509 117272 26514 117328
rect 26570 117272 234618 117328
rect 234674 117272 234679 117328
rect 26509 117270 234679 117272
rect 26509 117267 26575 117270
rect 234613 117267 234679 117270
rect 271137 117330 271203 117333
rect 272885 117330 272951 117333
rect 271137 117328 272951 117330
rect 271137 117272 271142 117328
rect 271198 117272 272890 117328
rect 272946 117272 272951 117328
rect 271137 117270 272951 117272
rect 271137 117267 271203 117270
rect 272885 117267 272951 117270
rect 273897 117330 273963 117333
rect 276381 117330 276447 117333
rect 273897 117328 276447 117330
rect 273897 117272 273902 117328
rect 273958 117272 276386 117328
rect 276442 117272 276447 117328
rect 273897 117270 276447 117272
rect 273897 117267 273963 117270
rect 276381 117267 276447 117270
rect 100293 117194 100359 117197
rect 106181 117194 106247 117197
rect 100293 117192 106247 117194
rect 100293 117136 100298 117192
rect 100354 117136 106186 117192
rect 106242 117136 106247 117192
rect 100293 117134 106247 117136
rect 100293 117131 100359 117134
rect 106181 117131 106247 117134
rect 129825 117194 129891 117197
rect 191741 117194 191807 117197
rect 129825 117192 191807 117194
rect 129825 117136 129830 117192
rect 129886 117136 191746 117192
rect 191802 117136 191807 117192
rect 129825 117134 191807 117136
rect 129825 117131 129891 117134
rect 191741 117131 191807 117134
rect 46841 117058 46907 117061
rect 98545 117058 98611 117061
rect 107561 117058 107627 117061
rect 46841 117056 64890 117058
rect 46841 117000 46846 117056
rect 46902 117000 64890 117056
rect 46841 116998 64890 117000
rect 46841 116995 46907 116998
rect 64830 116922 64890 116998
rect 98545 117056 107627 117058
rect 98545 117000 98550 117056
rect 98606 117000 107566 117056
rect 107622 117000 107627 117056
rect 98545 116998 107627 117000
rect 98545 116995 98611 116998
rect 107561 116995 107627 116998
rect 131205 117058 131271 117061
rect 355501 117058 355567 117061
rect 131205 117056 355567 117058
rect 131205 117000 131210 117056
rect 131266 117000 355506 117056
rect 355562 117000 355567 117056
rect 131205 116998 355567 117000
rect 131205 116995 131271 116998
rect 355501 116995 355567 116998
rect 68829 116922 68895 116925
rect 241421 116922 241487 116925
rect 407205 116922 407271 116925
rect 64830 116920 241487 116922
rect 64830 116864 68834 116920
rect 68890 116864 241426 116920
rect 241482 116864 241487 116920
rect 64830 116862 241487 116864
rect 404892 116920 407271 116922
rect 404892 116864 407210 116920
rect 407266 116864 407271 116920
rect 404892 116862 407271 116864
rect 68829 116859 68895 116862
rect 241421 116859 241487 116862
rect 407205 116859 407271 116862
rect 190821 116786 190887 116789
rect 280889 116786 280955 116789
rect 190821 116784 280955 116786
rect 190821 116728 190826 116784
rect 190882 116728 280894 116784
rect 280950 116728 280955 116784
rect 190821 116726 280955 116728
rect 190821 116723 190887 116726
rect 280889 116723 280955 116726
rect 126973 116650 127039 116653
rect 280838 116650 280844 116652
rect 126973 116648 280844 116650
rect 126973 116592 126978 116648
rect 127034 116592 280844 116648
rect 126973 116590 280844 116592
rect 126973 116587 127039 116590
rect 280838 116588 280844 116590
rect 280908 116588 280914 116652
rect 106917 116514 106983 116517
rect 286501 116514 286567 116517
rect 106917 116512 286567 116514
rect 106917 116456 106922 116512
rect 106978 116456 286506 116512
rect 286562 116456 286567 116512
rect 106917 116454 286567 116456
rect 106917 116451 106983 116454
rect 286501 116451 286567 116454
rect 125501 116378 125567 116381
rect 212441 116378 212507 116381
rect 280613 116378 280679 116381
rect 125501 116376 212507 116378
rect 125501 116320 125506 116376
rect 125562 116320 212446 116376
rect 212502 116320 212507 116376
rect 125501 116318 212507 116320
rect 125501 116315 125567 116318
rect 212441 116315 212507 116318
rect 219390 116376 280679 116378
rect 219390 116320 280618 116376
rect 280674 116320 280679 116376
rect 219390 116318 280679 116320
rect 212165 116242 212231 116245
rect 219390 116242 219450 116318
rect 280613 116315 280679 116318
rect 302734 116316 302740 116380
rect 302804 116378 302810 116380
rect 302804 116318 360180 116378
rect 302804 116316 302810 116318
rect 212165 116240 219450 116242
rect 212165 116184 212170 116240
rect 212226 116184 219450 116240
rect 212165 116182 219450 116184
rect 240501 116242 240567 116245
rect 280337 116242 280403 116245
rect 240501 116240 280403 116242
rect 240501 116184 240506 116240
rect 240562 116184 280342 116240
rect 280398 116184 280403 116240
rect 240501 116182 280403 116184
rect 212165 116179 212231 116182
rect 240501 116179 240567 116182
rect 280337 116179 280403 116182
rect 54334 116044 54340 116108
rect 54404 116106 54410 116108
rect 291326 116106 291332 116108
rect 54404 116046 291332 116106
rect 54404 116044 54410 116046
rect 291326 116044 291332 116046
rect 291396 116044 291402 116108
rect 7557 115970 7623 115973
rect 7557 115968 120090 115970
rect 7557 115912 7562 115968
rect 7618 115912 120090 115968
rect 7557 115910 120090 115912
rect 7557 115907 7623 115910
rect 120030 115698 120090 115910
rect 125225 115834 125291 115837
rect 355317 115834 355383 115837
rect 125225 115832 355383 115834
rect 125225 115776 125230 115832
rect 125286 115776 355322 115832
rect 355378 115776 355383 115832
rect 125225 115774 355383 115776
rect 125225 115771 125291 115774
rect 355317 115771 355383 115774
rect 121269 115698 121335 115701
rect 131205 115698 131271 115701
rect 352741 115698 352807 115701
rect 120030 115696 352807 115698
rect 120030 115640 121274 115696
rect 121330 115640 131210 115696
rect 131266 115640 352746 115696
rect 352802 115640 352807 115696
rect 120030 115638 352807 115640
rect 121269 115635 121335 115638
rect 131205 115635 131271 115638
rect 352741 115635 352807 115638
rect 119521 115562 119587 115565
rect 133873 115562 133939 115565
rect 352557 115562 352623 115565
rect 119521 115560 352623 115562
rect 119521 115504 119526 115560
rect 119582 115504 133878 115560
rect 133934 115504 352562 115560
rect 352618 115504 352623 115560
rect 119521 115502 352623 115504
rect 119521 115499 119587 115502
rect 133873 115499 133939 115502
rect 352557 115499 352623 115502
rect 123569 115426 123635 115429
rect 135253 115426 135319 115429
rect 352925 115426 352991 115429
rect 123569 115424 352991 115426
rect 123569 115368 123574 115424
rect 123630 115368 135258 115424
rect 135314 115368 352930 115424
rect 352986 115368 352991 115424
rect 123569 115366 352991 115368
rect 123569 115363 123635 115366
rect 135253 115363 135319 115366
rect 352925 115363 352991 115366
rect 63585 115290 63651 115293
rect 234613 115290 234679 115293
rect 63585 115288 234679 115290
rect 63585 115232 63590 115288
rect 63646 115232 234618 115288
rect 234674 115232 234679 115288
rect 63585 115230 234679 115232
rect 63585 115227 63651 115230
rect 234613 115227 234679 115230
rect 235390 115228 235396 115292
rect 235460 115290 235466 115292
rect 291142 115290 291148 115292
rect 235460 115230 291148 115290
rect 235460 115228 235466 115230
rect 291142 115228 291148 115230
rect 291212 115228 291218 115292
rect 294638 115228 294644 115292
rect 294708 115290 294714 115292
rect 294708 115230 360180 115290
rect 294708 115228 294714 115230
rect 180241 115154 180307 115157
rect 282269 115154 282335 115157
rect 180241 115152 282335 115154
rect 180241 115096 180246 115152
rect 180302 115096 282274 115152
rect 282330 115096 282335 115152
rect 180241 115094 282335 115096
rect 180241 115091 180307 115094
rect 282269 115091 282335 115094
rect 215661 115018 215727 115021
rect 280521 115018 280587 115021
rect 215661 115016 280587 115018
rect 215661 114960 215666 115016
rect 215722 114960 280526 115016
rect 280582 114960 280587 115016
rect 215661 114958 280587 114960
rect 215661 114955 215727 114958
rect 280521 114955 280587 114958
rect 176653 114474 176719 114477
rect 280705 114474 280771 114477
rect 176653 114472 280771 114474
rect 176653 114416 176658 114472
rect 176714 114416 280710 114472
rect 280766 114416 280771 114472
rect 176653 114414 280771 114416
rect 176653 114411 176719 114414
rect 280705 114411 280771 114414
rect 166073 114338 166139 114341
rect 281758 114338 281764 114340
rect 166073 114336 281764 114338
rect 166073 114280 166078 114336
rect 166134 114280 281764 114336
rect 166073 114278 281764 114280
rect 166073 114275 166139 114278
rect 281758 114276 281764 114278
rect 281828 114276 281834 114340
rect 112805 114202 112871 114205
rect 155217 114202 155283 114205
rect 112805 114200 155283 114202
rect 112805 114144 112810 114200
rect 112866 114144 155222 114200
rect 155278 114144 155283 114200
rect 112805 114142 155283 114144
rect 112805 114139 112871 114142
rect 155217 114139 155283 114142
rect 162485 114202 162551 114205
rect 289905 114202 289971 114205
rect 162485 114200 289971 114202
rect 162485 114144 162490 114200
rect 162546 114144 289910 114200
rect 289966 114144 289971 114200
rect 162485 114142 289971 114144
rect 162485 114139 162551 114142
rect 289905 114139 289971 114142
rect 299974 114140 299980 114204
rect 300044 114202 300050 114204
rect 300044 114142 360180 114202
rect 300044 114140 300050 114142
rect 148317 114066 148383 114069
rect 286409 114066 286475 114069
rect 148317 114064 286475 114066
rect 148317 114008 148322 114064
rect 148378 114008 286414 114064
rect 286470 114008 286475 114064
rect 148317 114006 286475 114008
rect 148317 114003 148383 114006
rect 286409 114003 286475 114006
rect 137645 113930 137711 113933
rect 292757 113930 292823 113933
rect 137645 113928 292823 113930
rect 137645 113872 137650 113928
rect 137706 113872 292762 113928
rect 292818 113872 292823 113928
rect 137645 113870 292823 113872
rect 137645 113867 137711 113870
rect 292757 113867 292823 113870
rect 110505 113794 110571 113797
rect 294137 113794 294203 113797
rect 110505 113792 294203 113794
rect 110505 113736 110510 113792
rect 110566 113736 294142 113792
rect 294198 113736 294203 113792
rect 110505 113734 294203 113736
rect 110505 113731 110571 113734
rect 294137 113731 294203 113734
rect 251173 113658 251239 113661
rect 285029 113658 285095 113661
rect 251173 113656 285095 113658
rect 251173 113600 251178 113656
rect 251234 113600 285034 113656
rect 285090 113600 285095 113656
rect 251173 113598 285095 113600
rect 251173 113595 251239 113598
rect 285029 113595 285095 113598
rect 3366 113188 3372 113252
rect 3436 113250 3442 113252
rect 252461 113250 252527 113253
rect 3436 113248 252527 113250
rect 3436 113192 252466 113248
rect 252522 113192 252527 113248
rect 3436 113190 252527 113192
rect 3436 113188 3442 113190
rect 252461 113187 252527 113190
rect 357934 113052 357940 113116
rect 358004 113114 358010 113116
rect 358004 113054 360180 113114
rect 358004 113052 358010 113054
rect 170397 112842 170463 112845
rect 282177 112842 282243 112845
rect 170397 112840 282243 112842
rect 170397 112784 170402 112840
rect 170458 112784 282182 112840
rect 282238 112784 282243 112840
rect 170397 112782 282243 112784
rect 170397 112779 170463 112782
rect 282177 112779 282243 112782
rect 580206 112780 580212 112844
rect 580276 112842 580282 112844
rect 583520 112842 584960 112932
rect 580276 112782 584960 112842
rect 580276 112780 580282 112782
rect 13537 112706 13603 112709
rect 186957 112706 187023 112709
rect 13537 112704 187023 112706
rect 13537 112648 13542 112704
rect 13598 112648 186962 112704
rect 187018 112648 187023 112704
rect 13537 112646 187023 112648
rect 13537 112643 13603 112646
rect 186957 112643 187023 112646
rect 205081 112706 205147 112709
rect 280429 112706 280495 112709
rect 205081 112704 280495 112706
rect 205081 112648 205086 112704
rect 205142 112648 280434 112704
rect 280490 112648 280495 112704
rect 205081 112646 280495 112648
rect 205081 112643 205147 112646
rect 280429 112643 280495 112646
rect 356646 112644 356652 112708
rect 356716 112706 356722 112708
rect 356716 112646 360210 112706
rect 583520 112692 584960 112782
rect 356716 112644 356722 112646
rect 85665 112570 85731 112573
rect 287881 112570 287947 112573
rect 85665 112568 287947 112570
rect 85665 112512 85670 112568
rect 85726 112512 287886 112568
rect 287942 112512 287947 112568
rect 85665 112510 287947 112512
rect 85665 112507 85731 112510
rect 287881 112507 287947 112510
rect 288934 112508 288940 112572
rect 289004 112570 289010 112572
rect 289004 112510 357450 112570
rect 289004 112508 289010 112510
rect 46054 112372 46060 112436
rect 46124 112434 46130 112436
rect 291878 112434 291884 112436
rect 46124 112374 291884 112434
rect 46124 112372 46130 112374
rect 291878 112372 291884 112374
rect 291948 112372 291954 112436
rect 357390 111754 357450 112510
rect 360150 111996 360210 112646
rect 357390 111694 360210 111754
rect 222745 111482 222811 111485
rect 280153 111482 280219 111485
rect 222745 111480 280219 111482
rect 222745 111424 222750 111480
rect 222806 111424 280158 111480
rect 280214 111424 280219 111480
rect 222745 111422 280219 111424
rect 222745 111419 222811 111422
rect 280153 111419 280219 111422
rect 183737 111346 183803 111349
rect 281901 111346 281967 111349
rect 183737 111344 281967 111346
rect 183737 111288 183742 111344
rect 183798 111288 281906 111344
rect 281962 111288 281967 111344
rect 183737 111286 281967 111288
rect 183737 111283 183803 111286
rect 281901 111283 281967 111286
rect 87965 111210 88031 111213
rect 226977 111210 227043 111213
rect 87965 111208 227043 111210
rect 87965 111152 87970 111208
rect 88026 111152 226982 111208
rect 227038 111152 227043 111208
rect 87965 111150 227043 111152
rect 87965 111147 88031 111150
rect 226977 111147 227043 111150
rect 114001 111074 114067 111077
rect 287605 111074 287671 111077
rect 114001 111072 287671 111074
rect 114001 111016 114006 111072
rect 114062 111016 287610 111072
rect 287666 111016 287671 111072
rect 114001 111014 287671 111016
rect 114001 111011 114067 111014
rect 287605 111011 287671 111014
rect 305494 111012 305500 111076
rect 305564 111074 305570 111076
rect 305564 111014 357450 111074
rect 305564 111012 305570 111014
rect -960 110666 480 110756
rect 119521 110666 119587 110669
rect -960 110664 119587 110666
rect -960 110608 119526 110664
rect 119582 110608 119587 110664
rect -960 110606 119587 110608
rect -960 110516 480 110606
rect 119521 110603 119587 110606
rect 357390 110394 357450 111014
rect 360150 110908 360210 111694
rect 357390 110334 360210 110394
rect 119889 109986 119955 109989
rect 159357 109986 159423 109989
rect 119889 109984 159423 109986
rect 119889 109928 119894 109984
rect 119950 109928 159362 109984
rect 159418 109928 159423 109984
rect 119889 109926 159423 109928
rect 119889 109923 119955 109926
rect 159357 109923 159423 109926
rect 195237 109986 195303 109989
rect 281809 109986 281875 109989
rect 195237 109984 281875 109986
rect 195237 109928 195242 109984
rect 195298 109928 281814 109984
rect 281870 109928 281875 109984
rect 195237 109926 281875 109928
rect 195237 109923 195303 109926
rect 281809 109923 281875 109926
rect 18229 109850 18295 109853
rect 130377 109850 130443 109853
rect 18229 109848 130443 109850
rect 18229 109792 18234 109848
rect 18290 109792 130382 109848
rect 130438 109792 130443 109848
rect 18229 109790 130443 109792
rect 18229 109787 18295 109790
rect 130377 109787 130443 109790
rect 144729 109850 144795 109853
rect 286317 109850 286383 109853
rect 144729 109848 286383 109850
rect 144729 109792 144734 109848
rect 144790 109792 286322 109848
rect 286378 109792 286383 109848
rect 360150 109820 360210 110334
rect 144729 109790 286383 109792
rect 144729 109787 144795 109790
rect 286317 109787 286383 109790
rect 32397 109714 32463 109717
rect 284886 109714 284892 109716
rect 32397 109712 284892 109714
rect 32397 109656 32402 109712
rect 32458 109656 284892 109712
rect 32397 109654 284892 109656
rect 32397 109651 32463 109654
rect 284886 109652 284892 109654
rect 284956 109652 284962 109716
rect 295926 109652 295932 109716
rect 295996 109714 296002 109716
rect 295996 109654 357450 109714
rect 295996 109652 296002 109654
rect 357390 109034 357450 109654
rect 357390 108974 360210 109034
rect 360150 108732 360210 108974
rect 208577 108626 208643 108629
rect 285121 108626 285187 108629
rect 208577 108624 285187 108626
rect 208577 108568 208582 108624
rect 208638 108568 285126 108624
rect 285182 108568 285187 108624
rect 208577 108566 285187 108568
rect 208577 108563 208643 108566
rect 285121 108563 285187 108566
rect 98637 108490 98703 108493
rect 222837 108490 222903 108493
rect 98637 108488 222903 108490
rect 98637 108432 98642 108488
rect 98698 108432 222842 108488
rect 222898 108432 222903 108488
rect 98637 108430 222903 108432
rect 98637 108427 98703 108430
rect 222837 108427 222903 108430
rect 226333 108490 226399 108493
rect 286133 108490 286199 108493
rect 226333 108488 286199 108490
rect 226333 108432 226338 108488
rect 226394 108432 286138 108488
rect 286194 108432 286199 108488
rect 226333 108430 286199 108432
rect 226333 108427 226399 108430
rect 286133 108427 286199 108430
rect 155401 108354 155467 108357
rect 283741 108354 283807 108357
rect 155401 108352 283807 108354
rect 155401 108296 155406 108352
rect 155462 108296 283746 108352
rect 283802 108296 283807 108352
rect 155401 108294 283807 108296
rect 155401 108291 155467 108294
rect 283741 108291 283807 108294
rect 304206 107612 304212 107676
rect 304276 107674 304282 107676
rect 304276 107614 360180 107674
rect 304276 107612 304282 107614
rect 197905 107130 197971 107133
rect 283557 107130 283623 107133
rect 197905 107128 283623 107130
rect 197905 107072 197910 107128
rect 197966 107072 283562 107128
rect 283618 107072 283623 107128
rect 197905 107070 283623 107072
rect 197905 107067 197971 107070
rect 283557 107067 283623 107070
rect 18597 106994 18663 106997
rect 243353 106994 243419 106997
rect 18597 106992 243419 106994
rect 18597 106936 18602 106992
rect 18658 106936 243358 106992
rect 243414 106936 243419 106992
rect 18597 106934 243419 106936
rect 18597 106931 18663 106934
rect 243353 106931 243419 106934
rect 43069 106858 43135 106861
rect 289077 106858 289143 106861
rect 43069 106856 289143 106858
rect 43069 106800 43074 106856
rect 43130 106800 289082 106856
rect 289138 106800 289143 106856
rect 43069 106798 289143 106800
rect 43069 106795 43135 106798
rect 289077 106795 289143 106798
rect 322054 106524 322060 106588
rect 322124 106586 322130 106588
rect 322124 106526 360180 106586
rect 322124 106524 322130 106526
rect 219249 105770 219315 105773
rect 286041 105770 286107 105773
rect 407113 105770 407179 105773
rect 219249 105768 286107 105770
rect 219249 105712 219254 105768
rect 219310 105712 286046 105768
rect 286102 105712 286107 105768
rect 219249 105710 286107 105712
rect 404892 105768 407179 105770
rect 404892 105712 407118 105768
rect 407174 105712 407179 105768
rect 404892 105710 407179 105712
rect 219249 105707 219315 105710
rect 286041 105707 286107 105710
rect 407113 105707 407179 105710
rect 104525 105634 104591 105637
rect 272057 105634 272123 105637
rect 104525 105632 272123 105634
rect 104525 105576 104530 105632
rect 104586 105576 272062 105632
rect 272118 105576 272123 105632
rect 104525 105574 272123 105576
rect 104525 105571 104591 105574
rect 272057 105571 272123 105574
rect 99833 105498 99899 105501
rect 287513 105498 287579 105501
rect 99833 105496 287579 105498
rect 99833 105440 99838 105496
rect 99894 105440 287518 105496
rect 287574 105440 287579 105496
rect 99833 105438 287579 105440
rect 99833 105435 99899 105438
rect 287513 105435 287579 105438
rect 323526 105436 323532 105500
rect 323596 105498 323602 105500
rect 323596 105438 360180 105498
rect 323596 105436 323602 105438
rect 233417 104410 233483 104413
rect 285949 104410 286015 104413
rect 233417 104408 286015 104410
rect 233417 104352 233422 104408
rect 233478 104352 285954 104408
rect 286010 104352 286015 104408
rect 233417 104350 286015 104352
rect 233417 104347 233483 104350
rect 285949 104347 286015 104350
rect 311014 104348 311020 104412
rect 311084 104410 311090 104412
rect 311084 104350 360180 104410
rect 311084 104348 311090 104350
rect 101029 104274 101095 104277
rect 270861 104274 270927 104277
rect 101029 104272 270927 104274
rect 101029 104216 101034 104272
rect 101090 104216 270866 104272
rect 270922 104216 270927 104272
rect 101029 104214 270927 104216
rect 101029 104211 101095 104214
rect 270861 104211 270927 104214
rect 9949 104138 10015 104141
rect 281022 104138 281028 104140
rect 9949 104136 281028 104138
rect 9949 104080 9954 104136
rect 10010 104080 281028 104136
rect 9949 104078 281028 104080
rect 9949 104075 10015 104078
rect 281022 104076 281028 104078
rect 281092 104076 281098 104140
rect 291694 103260 291700 103324
rect 291764 103322 291770 103324
rect 291764 103262 360180 103322
rect 291764 103260 291770 103262
rect 116393 103050 116459 103053
rect 211797 103050 211863 103053
rect 116393 103048 211863 103050
rect 116393 102992 116398 103048
rect 116454 102992 211802 103048
rect 211858 102992 211863 103048
rect 116393 102990 211863 102992
rect 116393 102987 116459 102990
rect 211797 102987 211863 102990
rect 93945 102914 94011 102917
rect 268377 102914 268443 102917
rect 93945 102912 268443 102914
rect 93945 102856 93950 102912
rect 94006 102856 268382 102912
rect 268438 102856 268443 102912
rect 93945 102854 268443 102856
rect 93945 102851 94011 102854
rect 268377 102851 268443 102854
rect 46657 102778 46723 102781
rect 288893 102778 288959 102781
rect 46657 102776 288959 102778
rect 46657 102720 46662 102776
rect 46718 102720 288898 102776
rect 288954 102720 288959 102776
rect 46657 102718 288959 102720
rect 46657 102715 46723 102718
rect 288893 102715 288959 102718
rect 187325 101690 187391 101693
rect 281717 101690 281783 101693
rect 187325 101688 281783 101690
rect 187325 101632 187330 101688
rect 187386 101632 281722 101688
rect 281778 101632 281783 101688
rect 187325 101630 281783 101632
rect 187325 101627 187391 101630
rect 281717 101627 281783 101630
rect 91553 101554 91619 101557
rect 228357 101554 228423 101557
rect 91553 101552 228423 101554
rect 91553 101496 91558 101552
rect 91614 101496 228362 101552
rect 228418 101496 228423 101552
rect 91553 101494 228423 101496
rect 91553 101491 91619 101494
rect 228357 101491 228423 101494
rect 35985 101418 36051 101421
rect 288985 101418 289051 101421
rect 35985 101416 289051 101418
rect 35985 101360 35990 101416
rect 36046 101360 288990 101416
rect 289046 101360 289051 101416
rect 35985 101358 289051 101360
rect 35985 101355 36051 101358
rect 288985 101355 289051 101358
rect 239622 100676 239628 100740
rect 239692 100738 239698 100740
rect 580206 100738 580212 100740
rect 239692 100678 580212 100738
rect 239692 100676 239698 100678
rect 580206 100676 580212 100678
rect 580276 100676 580282 100740
rect 291837 100602 291903 100605
rect 407205 100602 407271 100605
rect 291837 100600 407271 100602
rect 291837 100544 291842 100600
rect 291898 100544 407210 100600
rect 407266 100544 407271 100600
rect 291837 100542 407271 100544
rect 291837 100539 291903 100542
rect 407205 100539 407271 100542
rect 102777 100194 102843 100197
rect 282361 100194 282427 100197
rect 102777 100192 282427 100194
rect 102777 100136 102782 100192
rect 102838 100136 282366 100192
rect 282422 100136 282427 100192
rect 102777 100134 282427 100136
rect 102777 100131 102843 100134
rect 282361 100131 282427 100134
rect 11697 100058 11763 100061
rect 240869 100058 240935 100061
rect 11697 100056 240935 100058
rect 11697 100000 11702 100056
rect 11758 100000 240874 100056
rect 240930 100000 240935 100056
rect 11697 99998 240935 100000
rect 11697 99995 11763 99998
rect 240869 99995 240935 99998
rect 313774 99452 313780 99516
rect 313844 99514 313850 99516
rect 583520 99514 584960 99604
rect 313844 99454 584960 99514
rect 313844 99452 313850 99454
rect 583520 99364 584960 99454
rect 86861 98970 86927 98973
rect 265985 98970 266051 98973
rect 86861 98968 266051 98970
rect 86861 98912 86866 98968
rect 86922 98912 265990 98968
rect 266046 98912 266051 98968
rect 86861 98910 266051 98912
rect 86861 98907 86927 98910
rect 265985 98907 266051 98910
rect 14733 98834 14799 98837
rect 283230 98834 283236 98836
rect 14733 98832 283236 98834
rect 14733 98776 14738 98832
rect 14794 98776 283236 98832
rect 14733 98774 283236 98776
rect 14733 98771 14799 98774
rect 283230 98772 283236 98774
rect 283300 98772 283306 98836
rect 239438 98636 239444 98700
rect 239508 98698 239514 98700
rect 580206 98698 580212 98700
rect 239508 98638 580212 98698
rect 239508 98636 239514 98638
rect 580206 98636 580212 98638
rect 580276 98636 580282 98700
rect 320817 97882 320883 97885
rect 382457 97882 382523 97885
rect 320817 97880 382523 97882
rect 320817 97824 320822 97880
rect 320878 97824 382462 97880
rect 382518 97824 382523 97880
rect 320817 97822 382523 97824
rect 320817 97819 320883 97822
rect 382457 97819 382523 97822
rect -960 97610 480 97700
rect 290590 97610 290596 97612
rect -960 97550 290596 97610
rect -960 97460 480 97550
rect 290590 97548 290596 97550
rect 290660 97548 290666 97612
rect 97441 97338 97507 97341
rect 269573 97338 269639 97341
rect 97441 97336 269639 97338
rect 97441 97280 97446 97336
rect 97502 97280 269578 97336
rect 269634 97280 269639 97336
rect 97441 97278 269639 97280
rect 97441 97275 97507 97278
rect 269573 97275 269639 97278
rect 34789 97202 34855 97205
rect 213177 97202 213243 97205
rect 34789 97200 213243 97202
rect 34789 97144 34794 97200
rect 34850 97144 213182 97200
rect 213238 97144 213243 97200
rect 34789 97142 213243 97144
rect 34789 97139 34855 97142
rect 213177 97139 213243 97142
rect 90357 95842 90423 95845
rect 267181 95842 267247 95845
rect 90357 95840 267247 95842
rect 90357 95784 90362 95840
rect 90418 95784 267186 95840
rect 267242 95784 267247 95840
rect 90357 95782 267247 95784
rect 90357 95779 90423 95782
rect 267181 95779 267247 95782
rect 201493 94754 201559 94757
rect 284753 94754 284819 94757
rect 201493 94752 284819 94754
rect 201493 94696 201498 94752
rect 201554 94696 284758 94752
rect 284814 94696 284819 94752
rect 201493 94694 284819 94696
rect 201493 94691 201559 94694
rect 284753 94691 284819 94694
rect 95141 94618 95207 94621
rect 209037 94618 209103 94621
rect 95141 94616 209103 94618
rect 95141 94560 95146 94616
rect 95202 94560 209042 94616
rect 209098 94560 209103 94616
rect 95141 94558 209103 94560
rect 95141 94555 95207 94558
rect 209037 94555 209103 94558
rect 24209 94482 24275 94485
rect 278814 94482 278820 94484
rect 24209 94480 278820 94482
rect 24209 94424 24214 94480
rect 24270 94424 278820 94480
rect 24209 94422 278820 94424
rect 24209 94419 24275 94422
rect 278814 94420 278820 94422
rect 278884 94420 278890 94484
rect 23013 93394 23079 93397
rect 141417 93394 141483 93397
rect 23013 93392 141483 93394
rect 23013 93336 23018 93392
rect 23074 93336 141422 93392
rect 141478 93336 141483 93392
rect 23013 93334 141483 93336
rect 23013 93331 23079 93334
rect 141417 93331 141483 93334
rect 141233 93258 141299 93261
rect 284937 93258 285003 93261
rect 141233 93256 285003 93258
rect 141233 93200 141238 93256
rect 141294 93200 284942 93256
rect 284998 93200 285003 93256
rect 141233 93198 285003 93200
rect 141233 93195 141299 93198
rect 284937 93195 285003 93198
rect 118785 93122 118851 93125
rect 273897 93122 273963 93125
rect 118785 93120 273963 93122
rect 118785 93064 118790 93120
rect 118846 93064 273902 93120
rect 273958 93064 273963 93120
rect 118785 93062 273963 93064
rect 118785 93059 118851 93062
rect 273897 93059 273963 93062
rect 38377 91898 38443 91901
rect 137277 91898 137343 91901
rect 38377 91896 137343 91898
rect 38377 91840 38382 91896
rect 38438 91840 137282 91896
rect 137338 91840 137343 91896
rect 38377 91838 137343 91840
rect 38377 91835 38443 91838
rect 137277 91835 137343 91838
rect 158897 91898 158963 91901
rect 284845 91898 284911 91901
rect 158897 91896 284911 91898
rect 158897 91840 158902 91896
rect 158958 91840 284850 91896
rect 284906 91840 284911 91896
rect 158897 91838 284911 91840
rect 158897 91835 158963 91838
rect 284845 91835 284911 91838
rect 115197 91762 115263 91765
rect 275553 91762 275619 91765
rect 115197 91760 275619 91762
rect 115197 91704 115202 91760
rect 115258 91704 275558 91760
rect 275614 91704 275619 91760
rect 115197 91702 275619 91704
rect 115197 91699 115263 91702
rect 275553 91699 275619 91702
rect 111609 90538 111675 90541
rect 274357 90538 274423 90541
rect 111609 90536 274423 90538
rect 111609 90480 111614 90536
rect 111670 90480 274362 90536
rect 274418 90480 274423 90536
rect 111609 90478 274423 90480
rect 111609 90475 111675 90478
rect 274357 90475 274423 90478
rect 39573 90402 39639 90405
rect 288801 90402 288867 90405
rect 39573 90400 288867 90402
rect 39573 90344 39578 90400
rect 39634 90344 288806 90400
rect 288862 90344 288867 90400
rect 39573 90342 288867 90344
rect 39573 90339 39639 90342
rect 288801 90339 288867 90342
rect 108113 89178 108179 89181
rect 271137 89178 271203 89181
rect 108113 89176 271203 89178
rect 108113 89120 108118 89176
rect 108174 89120 271142 89176
rect 271198 89120 271203 89176
rect 108113 89118 271203 89120
rect 108113 89115 108179 89118
rect 271137 89115 271203 89118
rect 28901 89042 28967 89045
rect 283649 89042 283715 89045
rect 28901 89040 283715 89042
rect 28901 88984 28906 89040
rect 28962 88984 283654 89040
rect 283710 88984 283715 89040
rect 28901 88982 283715 88984
rect 28901 88979 28967 88982
rect 283649 88979 283715 88982
rect 65609 87954 65675 87957
rect 87781 87954 87847 87957
rect 65609 87952 87847 87954
rect 65609 87896 65614 87952
rect 65670 87896 87786 87952
rect 87842 87896 87847 87952
rect 65609 87894 87847 87896
rect 65609 87891 65675 87894
rect 87781 87891 87847 87894
rect 54661 87818 54727 87821
rect 86401 87818 86467 87821
rect 54661 87816 86467 87818
rect 54661 87760 54666 87816
rect 54722 87760 86406 87816
rect 86462 87760 86467 87816
rect 54661 87758 86467 87760
rect 54661 87755 54727 87758
rect 86401 87755 86467 87758
rect 63861 87682 63927 87685
rect 84837 87682 84903 87685
rect 63861 87680 84903 87682
rect 63861 87624 63866 87680
rect 63922 87624 84842 87680
rect 84898 87624 84903 87680
rect 63861 87622 84903 87624
rect 63861 87619 63927 87622
rect 84837 87619 84903 87622
rect 62021 87546 62087 87549
rect 87597 87546 87663 87549
rect 62021 87544 87663 87546
rect 62021 87488 62026 87544
rect 62082 87488 87602 87544
rect 87658 87488 87663 87544
rect 62021 87486 87663 87488
rect 62021 87483 62087 87486
rect 87597 87483 87663 87486
rect 97257 87546 97323 87549
rect 281625 87546 281691 87549
rect 97257 87544 281691 87546
rect 97257 87488 97262 87544
rect 97318 87488 281630 87544
rect 281686 87488 281691 87544
rect 97257 87486 281691 87488
rect 97257 87483 97323 87486
rect 281625 87483 281691 87486
rect 59261 87410 59327 87413
rect 85021 87410 85087 87413
rect 59261 87408 85087 87410
rect 59261 87352 59266 87408
rect 59322 87352 85026 87408
rect 85082 87352 85087 87408
rect 59261 87350 85087 87352
rect 59261 87347 59327 87350
rect 85021 87347 85087 87350
rect 57605 87274 57671 87277
rect 86217 87274 86283 87277
rect 57605 87272 86283 87274
rect 57605 87216 57610 87272
rect 57666 87216 86222 87272
rect 86278 87216 86283 87272
rect 57605 87214 86283 87216
rect 57605 87211 57671 87214
rect 86217 87211 86283 87214
rect 56225 87138 56291 87141
rect 85205 87138 85271 87141
rect 56225 87136 85271 87138
rect 56225 87080 56230 87136
rect 56286 87080 85210 87136
rect 85266 87080 85271 87136
rect 56225 87078 85271 87080
rect 56225 87075 56291 87078
rect 85205 87075 85271 87078
rect 52913 87002 52979 87005
rect 60733 87002 60799 87005
rect 52913 87000 60799 87002
rect 52913 86944 52918 87000
rect 52974 86944 60738 87000
rect 60794 86944 60799 87000
rect 52913 86942 60799 86944
rect 52913 86939 52979 86942
rect 60733 86939 60799 86942
rect 3550 86260 3556 86324
rect 3620 86322 3626 86324
rect 228214 86322 228220 86324
rect 3620 86262 228220 86322
rect 3620 86260 3626 86262
rect 228214 86260 228220 86262
rect 228284 86260 228290 86324
rect 60733 86186 60799 86189
rect 304349 86186 304415 86189
rect 60733 86184 304415 86186
rect 60733 86128 60738 86184
rect 60794 86128 304354 86184
rect 304410 86128 304415 86184
rect 60733 86126 304415 86128
rect 60733 86123 60799 86126
rect 304349 86123 304415 86126
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 68645 86050 68711 86053
rect 275277 86050 275343 86053
rect 68645 86048 275343 86050
rect 68645 85992 68650 86048
rect 68706 85992 275282 86048
rect 275338 85992 275343 86048
rect 583520 86036 584960 86126
rect 68645 85990 275343 85992
rect 68645 85987 68711 85990
rect 275277 85987 275343 85990
rect 50981 85914 51047 85917
rect 271137 85914 271203 85917
rect 50981 85912 271203 85914
rect 50981 85856 50986 85912
rect 51042 85856 271142 85912
rect 271198 85856 271203 85912
rect 50981 85854 271203 85856
rect 50981 85851 51047 85854
rect 271137 85851 271203 85854
rect 60641 85778 60707 85781
rect 322105 85778 322171 85781
rect 60641 85776 322171 85778
rect 60641 85720 60646 85776
rect 60702 85720 322110 85776
rect 322166 85720 322171 85776
rect 60641 85718 322171 85720
rect 60641 85715 60707 85718
rect 322105 85715 322171 85718
rect 66989 85642 67055 85645
rect 336273 85642 336339 85645
rect 66989 85640 336339 85642
rect 66989 85584 66994 85640
rect 67050 85584 336278 85640
rect 336334 85584 336339 85640
rect 66989 85582 336339 85584
rect 66989 85579 67055 85582
rect 336273 85579 336339 85582
rect 80743 85098 80809 85101
rect 364609 85098 364675 85101
rect 80743 85096 364675 85098
rect 80743 85040 80748 85096
rect 80804 85040 364614 85096
rect 364670 85040 364675 85096
rect 80743 85038 364675 85040
rect 80743 85035 80809 85038
rect 364609 85035 364675 85038
rect 77615 84962 77681 84965
rect 357525 84962 357591 84965
rect 77615 84960 357591 84962
rect 77615 84904 77620 84960
rect 77676 84904 357530 84960
rect 357586 84904 357591 84960
rect 77615 84902 357591 84904
rect 77615 84899 77681 84902
rect 357525 84899 357591 84902
rect 69795 84826 69861 84829
rect 282177 84826 282243 84829
rect 69795 84824 282243 84826
rect -960 84690 480 84780
rect 69795 84768 69800 84824
rect 69856 84768 282182 84824
rect 282238 84768 282243 84824
rect 69795 84766 282243 84768
rect 69795 84763 69861 84766
rect 282177 84763 282243 84766
rect 3550 84690 3556 84692
rect -960 84630 3556 84690
rect -960 84540 480 84630
rect 3550 84628 3556 84630
rect 3620 84628 3626 84692
rect 71359 84690 71425 84693
rect 343357 84690 343423 84693
rect 71359 84688 343423 84690
rect 71359 84632 71364 84688
rect 71420 84632 343362 84688
rect 343418 84632 343423 84688
rect 71359 84630 343423 84632
rect 71359 84627 71425 84630
rect 343357 84627 343423 84630
rect 79179 84554 79245 84557
rect 361113 84554 361179 84557
rect 79179 84552 361179 84554
rect 79179 84496 79184 84552
rect 79240 84496 361118 84552
rect 361174 84496 361179 84552
rect 79179 84494 361179 84496
rect 79179 84491 79245 84494
rect 361113 84491 361179 84494
rect 82307 84280 82373 84285
rect 82307 84224 82312 84280
rect 82368 84224 82373 84280
rect 82307 84219 82373 84224
rect 82310 84146 82370 84219
rect 82310 84086 84210 84146
rect 84150 83466 84210 84086
rect 368197 83466 368263 83469
rect 84150 83464 368263 83466
rect 84150 83408 368202 83464
rect 368258 83408 368263 83464
rect 84150 83406 368263 83408
rect 368197 83403 368263 83406
rect 435357 83058 435423 83061
rect 84916 83056 435423 83058
rect 84916 83000 435362 83056
rect 435418 83000 435423 83056
rect 84916 82998 435423 83000
rect 435357 82995 435423 82998
rect 85205 82106 85271 82109
rect 311433 82106 311499 82109
rect 85205 82104 311499 82106
rect 85205 82048 85210 82104
rect 85266 82048 311438 82104
rect 311494 82048 311499 82104
rect 85205 82046 311499 82048
rect 85205 82043 85271 82046
rect 311433 82043 311499 82046
rect 48129 81698 48195 81701
rect 432597 81698 432663 81701
rect 48129 81696 50140 81698
rect 48129 81640 48134 81696
rect 48190 81640 50140 81696
rect 48129 81638 50140 81640
rect 84916 81696 432663 81698
rect 84916 81640 432602 81696
rect 432658 81640 432663 81696
rect 84916 81638 432663 81640
rect 48129 81635 48195 81638
rect 432597 81635 432663 81638
rect 85021 80746 85087 80749
rect 318517 80746 318583 80749
rect 85021 80744 318583 80746
rect 85021 80688 85026 80744
rect 85082 80688 318522 80744
rect 318578 80688 318583 80744
rect 85021 80686 318583 80688
rect 85021 80683 85087 80686
rect 318517 80683 318583 80686
rect 48221 80338 48287 80341
rect 428549 80338 428615 80341
rect 48221 80336 50140 80338
rect 48221 80280 48226 80336
rect 48282 80280 50140 80336
rect 48221 80278 50140 80280
rect 84916 80336 428615 80338
rect 84916 80280 428554 80336
rect 428610 80280 428615 80336
rect 84916 80278 428615 80280
rect 48221 80275 48287 80278
rect 428549 80275 428615 80278
rect 173157 79522 173223 79525
rect 282729 79522 282795 79525
rect 173157 79520 282795 79522
rect 173157 79464 173162 79520
rect 173218 79464 282734 79520
rect 282790 79464 282795 79520
rect 173157 79462 282795 79464
rect 173157 79459 173223 79462
rect 282729 79459 282795 79462
rect 84837 79386 84903 79389
rect 329189 79386 329255 79389
rect 84837 79384 329255 79386
rect 84837 79328 84842 79384
rect 84898 79328 329194 79384
rect 329250 79328 329255 79384
rect 84837 79326 329255 79328
rect 84837 79323 84903 79326
rect 329189 79323 329255 79326
rect 49325 78978 49391 78981
rect 105537 78978 105603 78981
rect 49325 78976 50140 78978
rect 49325 78920 49330 78976
rect 49386 78920 50140 78976
rect 49325 78918 50140 78920
rect 84916 78976 105603 78978
rect 84916 78920 105542 78976
rect 105598 78920 105603 78976
rect 84916 78918 105603 78920
rect 49325 78915 49391 78918
rect 105537 78915 105603 78918
rect 130561 77890 130627 77893
rect 283465 77890 283531 77893
rect 130561 77888 283531 77890
rect 130561 77832 130566 77888
rect 130622 77832 283470 77888
rect 283526 77832 283531 77888
rect 130561 77830 283531 77832
rect 130561 77827 130627 77830
rect 283465 77827 283531 77830
rect 421557 77618 421623 77621
rect 84916 77616 421623 77618
rect 50294 77349 50354 77588
rect 84916 77560 421562 77616
rect 421618 77560 421623 77616
rect 84916 77558 421623 77560
rect 421557 77555 421623 77558
rect 50245 77344 50354 77349
rect 50245 77288 50250 77344
rect 50306 77288 50354 77344
rect 50245 77286 50354 77288
rect 50245 77283 50311 77286
rect 134149 76530 134215 76533
rect 283373 76530 283439 76533
rect 134149 76528 283439 76530
rect 134149 76472 134154 76528
rect 134210 76472 283378 76528
rect 283434 76472 283439 76528
rect 134149 76470 283439 76472
rect 134149 76467 134215 76470
rect 283373 76467 283439 76470
rect 49601 76258 49667 76261
rect 417417 76258 417483 76261
rect 49601 76256 50140 76258
rect 49601 76200 49606 76256
rect 49662 76200 50140 76256
rect 49601 76198 50140 76200
rect 84916 76256 417483 76258
rect 84916 76200 417422 76256
rect 417478 76200 417483 76256
rect 84916 76198 417483 76200
rect 49601 76195 49667 76198
rect 417417 76195 417483 76198
rect 414657 74898 414723 74901
rect 84916 74896 414723 74898
rect 50294 74629 50354 74868
rect 84916 74840 414662 74896
rect 414718 74840 414723 74896
rect 84916 74838 414723 74840
rect 414657 74835 414723 74838
rect 50294 74624 50403 74629
rect 50294 74568 50342 74624
rect 50398 74568 50403 74624
rect 50294 74566 50403 74568
rect 50337 74563 50403 74566
rect 151813 73810 151879 73813
rect 285857 73810 285923 73813
rect 151813 73808 285923 73810
rect 151813 73752 151818 73808
rect 151874 73752 285862 73808
rect 285918 73752 285923 73808
rect 151813 73750 285923 73752
rect 151813 73747 151879 73750
rect 285857 73747 285923 73750
rect 49509 73538 49575 73541
rect 450537 73538 450603 73541
rect 49509 73536 50140 73538
rect 49509 73480 49514 73536
rect 49570 73480 50140 73536
rect 49509 73478 50140 73480
rect 84916 73536 450603 73538
rect 84916 73480 450542 73536
rect 450598 73480 450603 73536
rect 84916 73478 450603 73480
rect 49509 73475 49575 73478
rect 450537 73475 450603 73478
rect 580206 72932 580212 72996
rect 580276 72994 580282 72996
rect 583520 72994 584960 73084
rect 580276 72934 584960 72994
rect 580276 72932 580282 72934
rect 583520 72844 584960 72934
rect 89161 72450 89227 72453
rect 287421 72450 287487 72453
rect 89161 72448 287487 72450
rect 89161 72392 89166 72448
rect 89222 72392 287426 72448
rect 287482 72392 287487 72448
rect 89161 72390 287487 72392
rect 89161 72387 89227 72390
rect 287421 72387 287487 72390
rect 447777 72178 447843 72181
rect 84916 72176 447843 72178
rect 50110 71909 50170 72148
rect 84916 72120 447782 72176
rect 447838 72120 447843 72176
rect 84916 72118 447843 72120
rect 447777 72115 447843 72118
rect 50110 71904 50219 71909
rect 50110 71848 50158 71904
rect 50214 71848 50219 71904
rect 50110 71846 50219 71848
rect 50153 71843 50219 71846
rect -960 71634 480 71724
rect 7557 71634 7623 71637
rect -960 71632 7623 71634
rect -960 71576 7562 71632
rect 7618 71576 7623 71632
rect -960 71574 7623 71576
rect -960 71484 480 71574
rect 7557 71571 7623 71574
rect 49417 70818 49483 70821
rect 443637 70818 443703 70821
rect 49417 70816 50140 70818
rect 49417 70760 49422 70816
rect 49478 70760 50140 70816
rect 49417 70758 50140 70760
rect 84916 70816 443703 70818
rect 84916 70760 443642 70816
rect 443698 70760 443703 70816
rect 84916 70758 443703 70760
rect 49417 70755 49483 70758
rect 443637 70755 443703 70758
rect 278037 69458 278103 69461
rect 84916 69456 278103 69458
rect 50478 69053 50538 69428
rect 84916 69400 278042 69456
rect 278098 69400 278103 69456
rect 84916 69398 278103 69400
rect 278037 69395 278103 69398
rect 50429 69048 50538 69053
rect 50429 68992 50434 69048
rect 50490 68992 50538 69048
rect 50429 68990 50538 68992
rect 50429 68987 50495 68990
rect 49233 68098 49299 68101
rect 422937 68098 423003 68101
rect 49233 68096 50140 68098
rect 49233 68040 49238 68096
rect 49294 68040 50140 68096
rect 49233 68038 50140 68040
rect 84916 68096 423003 68098
rect 84916 68040 422942 68096
rect 422998 68040 423003 68096
rect 84916 68038 423003 68040
rect 49233 68035 49299 68038
rect 422937 68035 423003 68038
rect 49049 66738 49115 66741
rect 436737 66738 436803 66741
rect 49049 66736 50140 66738
rect 49049 66680 49054 66736
rect 49110 66680 50140 66736
rect 49049 66678 50140 66680
rect 84916 66736 436803 66738
rect 84916 66680 436742 66736
rect 436798 66680 436803 66736
rect 84916 66678 436803 66680
rect 49049 66675 49115 66678
rect 436737 66675 436803 66678
rect 47669 65378 47735 65381
rect 431217 65378 431283 65381
rect 47669 65376 50140 65378
rect 47669 65320 47674 65376
rect 47730 65320 50140 65376
rect 47669 65318 50140 65320
rect 84916 65376 431283 65378
rect 84916 65320 431222 65376
rect 431278 65320 431283 65376
rect 84916 65318 431283 65320
rect 47669 65315 47735 65318
rect 431217 65315 431283 65318
rect 96245 64154 96311 64157
rect 284661 64154 284727 64157
rect 96245 64152 284727 64154
rect 96245 64096 96250 64152
rect 96306 64096 284666 64152
rect 284722 64096 284727 64152
rect 96245 64094 284727 64096
rect 96245 64091 96311 64094
rect 284661 64091 284727 64094
rect 47945 64018 48011 64021
rect 429837 64018 429903 64021
rect 47945 64016 50140 64018
rect 47945 63960 47950 64016
rect 48006 63960 50140 64016
rect 47945 63958 50140 63960
rect 84916 64016 429903 64018
rect 84916 63960 429842 64016
rect 429898 63960 429903 64016
rect 84916 63958 429903 63960
rect 47945 63955 48011 63958
rect 429837 63955 429903 63958
rect 90449 62794 90515 62797
rect 281574 62794 281580 62796
rect 90449 62792 281580 62794
rect 90449 62736 90454 62792
rect 90510 62736 281580 62792
rect 90449 62734 281580 62736
rect 90449 62731 90515 62734
rect 281574 62732 281580 62734
rect 281644 62732 281650 62796
rect 47577 62658 47643 62661
rect 425697 62658 425763 62661
rect 47577 62656 50140 62658
rect 47577 62600 47582 62656
rect 47638 62600 50140 62656
rect 47577 62598 50140 62600
rect 84916 62656 425763 62658
rect 84916 62600 425702 62656
rect 425758 62600 425763 62656
rect 84916 62598 425763 62600
rect 47577 62595 47643 62598
rect 425697 62595 425763 62598
rect 124673 61434 124739 61437
rect 288709 61434 288775 61437
rect 124673 61432 288775 61434
rect 124673 61376 124678 61432
rect 124734 61376 288714 61432
rect 288770 61376 288775 61432
rect 124673 61374 288775 61376
rect 124673 61371 124739 61374
rect 288709 61371 288775 61374
rect 48037 61298 48103 61301
rect 418797 61298 418863 61301
rect 48037 61296 50140 61298
rect 48037 61240 48042 61296
rect 48098 61240 50140 61296
rect 48037 61238 50140 61240
rect 84916 61296 418863 61298
rect 84916 61240 418802 61296
rect 418858 61240 418863 61296
rect 84916 61238 418863 61240
rect 48037 61235 48103 61238
rect 418797 61235 418863 61238
rect 121085 60074 121151 60077
rect 288617 60074 288683 60077
rect 121085 60072 288683 60074
rect 121085 60016 121090 60072
rect 121146 60016 288622 60072
rect 288678 60016 288683 60072
rect 121085 60014 288683 60016
rect 121085 60011 121151 60014
rect 288617 60011 288683 60014
rect 47853 59938 47919 59941
rect 307109 59938 307175 59941
rect 47853 59936 50140 59938
rect 47853 59880 47858 59936
rect 47914 59880 50140 59936
rect 47853 59878 50140 59880
rect 84916 59936 307175 59938
rect 84916 59880 307114 59936
rect 307170 59880 307175 59936
rect 84916 59878 307175 59880
rect 47853 59875 47919 59878
rect 307109 59875 307175 59878
rect 306966 59604 306972 59668
rect 307036 59666 307042 59668
rect 583520 59666 584960 59756
rect 307036 59606 584960 59666
rect 307036 59604 307042 59606
rect 583520 59516 584960 59606
rect 117589 58714 117655 58717
rect 288525 58714 288591 58717
rect 117589 58712 288591 58714
rect -960 58578 480 58668
rect 117589 58656 117594 58712
rect 117650 58656 288530 58712
rect 288586 58656 288591 58712
rect 117589 58654 288591 58656
rect 117589 58651 117655 58654
rect 288525 58651 288591 58654
rect 46054 58578 46060 58580
rect -960 58518 46060 58578
rect -960 58428 480 58518
rect 46054 58516 46060 58518
rect 46124 58516 46130 58580
rect 47761 58578 47827 58581
rect 324957 58578 325023 58581
rect 47761 58576 50140 58578
rect 47761 58520 47766 58576
rect 47822 58520 50140 58576
rect 47761 58518 50140 58520
rect 84916 58576 325023 58578
rect 84916 58520 324962 58576
rect 325018 58520 325023 58576
rect 84916 58518 325023 58520
rect 47761 58515 47827 58518
rect 324957 58515 325023 58518
rect 123477 57354 123543 57357
rect 199377 57354 199443 57357
rect 123477 57352 199443 57354
rect 123477 57296 123482 57352
rect 123538 57296 199382 57352
rect 199438 57296 199443 57352
rect 123477 57294 199443 57296
rect 123477 57291 123543 57294
rect 199377 57291 199443 57294
rect 411897 57218 411963 57221
rect 84916 57216 411963 57218
rect 50478 56677 50538 57188
rect 84916 57160 411902 57216
rect 411958 57160 411963 57216
rect 84916 57158 411963 57160
rect 411897 57155 411963 57158
rect 50478 56672 50587 56677
rect 50478 56616 50526 56672
rect 50582 56616 50587 56672
rect 50478 56614 50587 56616
rect 50521 56611 50587 56614
rect 47485 55858 47551 55861
rect 105537 55858 105603 55861
rect 467465 55858 467531 55861
rect 47485 55856 50140 55858
rect 47485 55800 47490 55856
rect 47546 55800 50140 55856
rect 47485 55798 50140 55800
rect 105537 55856 467531 55858
rect 105537 55800 105542 55856
rect 105598 55800 467470 55856
rect 467526 55800 467531 55856
rect 105537 55798 467531 55800
rect 47485 55795 47551 55798
rect 105537 55795 105603 55798
rect 467465 55795 467531 55798
rect 84886 55722 84946 55760
rect 287697 55722 287763 55725
rect 84886 55720 287763 55722
rect 84886 55664 287702 55720
rect 287758 55664 287763 55720
rect 84886 55662 287763 55664
rect 287697 55659 287763 55662
rect 49141 54498 49207 54501
rect 266997 54498 267063 54501
rect 49141 54496 50140 54498
rect 49141 54440 49146 54496
rect 49202 54440 50140 54496
rect 49141 54438 50140 54440
rect 84916 54496 267063 54498
rect 84916 54440 267002 54496
rect 267058 54440 267063 54496
rect 84916 54438 267063 54440
rect 49141 54435 49207 54438
rect 266997 54435 267063 54438
rect 85573 53274 85639 53277
rect 138657 53274 138723 53277
rect 84886 53272 138723 53274
rect 84886 53216 85578 53272
rect 85634 53216 138662 53272
rect 138718 53216 138723 53272
rect 84886 53214 138723 53216
rect 84886 53108 84946 53214
rect 85573 53211 85639 53214
rect 138657 53211 138723 53214
rect 307109 53274 307175 53277
rect 421373 53274 421439 53277
rect 307109 53272 421439 53274
rect 307109 53216 307114 53272
rect 307170 53216 421378 53272
rect 421434 53216 421439 53272
rect 307109 53214 421439 53216
rect 307109 53211 307175 53214
rect 421373 53211 421439 53214
rect 86401 53138 86467 53141
rect 307937 53138 308003 53141
rect 86401 53136 308003 53138
rect 50478 52594 50538 53108
rect 86401 53080 86406 53136
rect 86462 53080 307942 53136
rect 307998 53080 308003 53136
rect 86401 53078 308003 53080
rect 86401 53075 86467 53078
rect 307937 53075 308003 53078
rect 50613 52594 50679 52597
rect 50478 52592 50679 52594
rect 50478 52536 50618 52592
rect 50674 52536 50679 52592
rect 50478 52534 50679 52536
rect 50613 52531 50679 52534
rect 86217 51778 86283 51781
rect 315021 51778 315087 51781
rect 86217 51776 315087 51778
rect 57830 51444 57836 51508
rect 57900 51506 57906 51508
rect 57900 51446 64890 51506
rect 57900 51444 57906 51446
rect 64830 51370 64890 51446
rect 84334 51370 84394 51748
rect 86217 51720 86222 51776
rect 86278 51720 315026 51776
rect 315082 51720 315087 51776
rect 86217 51718 315087 51720
rect 86217 51715 86283 51718
rect 315021 51715 315087 51718
rect 84469 51506 84535 51509
rect 215937 51506 216003 51509
rect 84469 51504 216003 51506
rect 84469 51448 84474 51504
rect 84530 51448 215942 51504
rect 215998 51448 216003 51504
rect 84469 51446 216003 51448
rect 84469 51443 84535 51446
rect 215937 51443 216003 51446
rect 64830 51310 84394 51370
rect 82077 50282 82143 50285
rect 287329 50282 287395 50285
rect 82077 50280 287395 50282
rect 82077 50224 82082 50280
rect 82138 50224 287334 50280
rect 287390 50224 287395 50280
rect 82077 50222 287395 50224
rect 82077 50219 82143 50222
rect 287329 50219 287395 50222
rect 48221 49330 48287 49333
rect 268837 49330 268903 49333
rect 48221 49328 268903 49330
rect 48221 49272 48226 49328
rect 48282 49272 268842 49328
rect 268898 49272 268903 49328
rect 48221 49270 268903 49272
rect 48221 49267 48287 49270
rect 268837 49267 268903 49270
rect 67909 49194 67975 49197
rect 291469 49194 291535 49197
rect 67909 49192 291535 49194
rect 67909 49136 67914 49192
rect 67970 49136 291474 49192
rect 291530 49136 291535 49192
rect 67909 49134 291535 49136
rect 67909 49131 67975 49134
rect 291469 49131 291535 49134
rect 49049 49058 49115 49061
rect 517145 49058 517211 49061
rect 49049 49056 517211 49058
rect 49049 49000 49054 49056
rect 49110 49000 517150 49056
rect 517206 49000 517211 49056
rect 49049 48998 517211 49000
rect 49049 48995 49115 48998
rect 517145 48995 517211 48998
rect 47945 48922 48011 48925
rect 576117 48922 576183 48925
rect 47945 48920 576183 48922
rect 47945 48864 47950 48920
rect 48006 48864 576122 48920
rect 576178 48864 576183 48920
rect 47945 48862 576183 48864
rect 47945 48859 48011 48862
rect 576117 48859 576183 48862
rect 60641 47970 60707 47973
rect 62757 47970 62823 47973
rect 60641 47968 62823 47970
rect 60641 47912 60646 47968
rect 60702 47912 62762 47968
rect 62818 47912 62823 47968
rect 60641 47910 62823 47912
rect 60641 47907 60707 47910
rect 62757 47907 62823 47910
rect 50981 47834 51047 47837
rect 439497 47834 439563 47837
rect 50981 47832 439563 47834
rect 50981 47776 50986 47832
rect 51042 47776 439502 47832
rect 439558 47776 439563 47832
rect 50981 47774 439563 47776
rect 50981 47771 51047 47774
rect 439497 47771 439563 47774
rect 52361 47698 52427 47701
rect 442257 47698 442323 47701
rect 52361 47696 442323 47698
rect 52361 47640 52366 47696
rect 52422 47640 442262 47696
rect 442318 47640 442323 47696
rect 52361 47638 442323 47640
rect 52361 47635 52427 47638
rect 442257 47635 442323 47638
rect 53741 47562 53807 47565
rect 446397 47562 446463 47565
rect 53741 47560 446463 47562
rect 53741 47504 53746 47560
rect 53802 47504 446402 47560
rect 446458 47504 446463 47560
rect 53741 47502 446463 47504
rect 53741 47499 53807 47502
rect 446397 47499 446463 47502
rect 64781 47018 64847 47021
rect 65609 47018 65675 47021
rect 64781 47016 65675 47018
rect 64781 46960 64786 47016
rect 64842 46960 65614 47016
rect 65670 46960 65675 47016
rect 64781 46958 65675 46960
rect 64781 46955 64847 46958
rect 65609 46955 65675 46958
rect 74441 47018 74507 47021
rect 75177 47018 75243 47021
rect 74441 47016 75243 47018
rect 74441 46960 74446 47016
rect 74502 46960 75182 47016
rect 75238 46960 75243 47016
rect 74441 46958 75243 46960
rect 74441 46955 74507 46958
rect 75177 46955 75243 46958
rect 56501 46338 56567 46341
rect 481725 46338 481791 46341
rect 56501 46336 481791 46338
rect 56501 46280 56506 46336
rect 56562 46280 481730 46336
rect 481786 46280 481791 46336
rect 56501 46278 481791 46280
rect 56501 46275 56567 46278
rect 481725 46275 481791 46278
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 565 46202 631 46205
rect 57830 46202 57836 46204
rect 565 46200 57836 46202
rect 565 46144 570 46200
rect 626 46144 57836 46200
rect 565 46142 57836 46144
rect 565 46139 631 46142
rect 57830 46140 57836 46142
rect 57900 46140 57906 46204
rect 74993 46202 75059 46205
rect 287237 46202 287303 46205
rect 74993 46200 287303 46202
rect 74993 46144 74998 46200
rect 75054 46144 287242 46200
rect 287298 46144 287303 46200
rect 583520 46188 584960 46278
rect 74993 46142 287303 46144
rect 74993 46139 75059 46142
rect 287237 46139 287303 46142
rect -960 45522 480 45612
rect 231158 45522 231164 45524
rect -960 45462 231164 45522
rect -960 45372 480 45462
rect 231158 45460 231164 45462
rect 231228 45460 231234 45524
rect 53741 44978 53807 44981
rect 280654 44978 280660 44980
rect 53741 44976 280660 44978
rect 53741 44920 53746 44976
rect 53802 44920 280660 44976
rect 53741 44918 280660 44920
rect 53741 44915 53807 44918
rect 280654 44916 280660 44918
rect 280724 44916 280730 44980
rect 49325 44842 49391 44845
rect 549069 44842 549135 44845
rect 49325 44840 549135 44842
rect 49325 44784 49330 44840
rect 49386 44784 549074 44840
rect 549130 44784 549135 44840
rect 49325 44782 549135 44784
rect 49325 44779 49391 44782
rect 549069 44779 549135 44782
rect 47669 43618 47735 43621
rect 284937 43618 285003 43621
rect 47669 43616 285003 43618
rect 47669 43560 47674 43616
rect 47730 43560 284942 43616
rect 284998 43560 285003 43616
rect 47669 43558 285003 43560
rect 47669 43555 47735 43558
rect 284937 43555 285003 43558
rect 63309 43482 63375 43485
rect 499389 43482 499455 43485
rect 63309 43480 499455 43482
rect 63309 43424 63314 43480
rect 63370 43424 499394 43480
rect 499450 43424 499455 43480
rect 63309 43422 499455 43424
rect 63309 43419 63375 43422
rect 499389 43419 499455 43422
rect 48129 42258 48195 42261
rect 289077 42258 289143 42261
rect 48129 42256 289143 42258
rect 48129 42200 48134 42256
rect 48190 42200 289082 42256
rect 289138 42200 289143 42256
rect 48129 42198 289143 42200
rect 48129 42195 48195 42198
rect 289077 42195 289143 42198
rect 66069 42122 66135 42125
rect 506473 42122 506539 42125
rect 66069 42120 506539 42122
rect 66069 42064 66074 42120
rect 66130 42064 506478 42120
rect 506534 42064 506539 42120
rect 66069 42062 506539 42064
rect 66069 42059 66135 42062
rect 506473 42059 506539 42062
rect 77109 40762 77175 40765
rect 389449 40762 389515 40765
rect 77109 40760 389515 40762
rect 77109 40704 77114 40760
rect 77170 40704 389454 40760
rect 389510 40704 389515 40760
rect 77109 40702 389515 40704
rect 77109 40699 77175 40702
rect 389449 40699 389515 40702
rect 68829 40626 68895 40629
rect 512637 40626 512703 40629
rect 68829 40624 512703 40626
rect 68829 40568 68834 40624
rect 68890 40568 512642 40624
rect 512698 40568 512703 40624
rect 68829 40566 512703 40568
rect 68829 40563 68895 40566
rect 512637 40563 512703 40566
rect 81249 39402 81315 39405
rect 400121 39402 400187 39405
rect 81249 39400 400187 39402
rect 81249 39344 81254 39400
rect 81310 39344 400126 39400
rect 400182 39344 400187 39400
rect 81249 39342 400187 39344
rect 81249 39339 81315 39342
rect 400121 39339 400187 39342
rect 49233 39266 49299 39269
rect 520733 39266 520799 39269
rect 49233 39264 520799 39266
rect 49233 39208 49238 39264
rect 49294 39208 520738 39264
rect 520794 39208 520799 39264
rect 49233 39206 520799 39208
rect 49233 39203 49299 39206
rect 520733 39203 520799 39206
rect 84009 38042 84075 38045
rect 407205 38042 407271 38045
rect 84009 38040 407271 38042
rect 84009 37984 84014 38040
rect 84070 37984 407210 38040
rect 407266 37984 407271 38040
rect 84009 37982 407271 37984
rect 84009 37979 84075 37982
rect 407205 37979 407271 37982
rect 50429 37906 50495 37909
rect 524229 37906 524295 37909
rect 50429 37904 524295 37906
rect 50429 37848 50434 37904
rect 50490 37848 524234 37904
rect 524290 37848 524295 37904
rect 50429 37846 524295 37848
rect 50429 37843 50495 37846
rect 524229 37843 524295 37846
rect 51349 36682 51415 36685
rect 254025 36682 254091 36685
rect 51349 36680 254091 36682
rect 51349 36624 51354 36680
rect 51410 36624 254030 36680
rect 254086 36624 254091 36680
rect 51349 36622 254091 36624
rect 51349 36619 51415 36622
rect 254025 36619 254091 36622
rect 49417 36546 49483 36549
rect 527817 36546 527883 36549
rect 49417 36544 527883 36546
rect 49417 36488 49422 36544
rect 49478 36488 527822 36544
rect 527878 36488 527883 36544
rect 49417 36486 527883 36488
rect 49417 36483 49483 36486
rect 527817 36483 527883 36486
rect 55857 35322 55923 35325
rect 255221 35322 255287 35325
rect 55857 35320 255287 35322
rect 55857 35264 55862 35320
rect 55918 35264 255226 35320
rect 255282 35264 255287 35320
rect 55857 35262 255287 35264
rect 55857 35259 55923 35262
rect 255221 35259 255287 35262
rect 49509 35186 49575 35189
rect 534901 35186 534967 35189
rect 49509 35184 534967 35186
rect 49509 35128 49514 35184
rect 49570 35128 534906 35184
rect 534962 35128 534967 35184
rect 49509 35126 534967 35128
rect 49509 35123 49575 35126
rect 534901 35123 534967 35126
rect 62849 33962 62915 33965
rect 257613 33962 257679 33965
rect 62849 33960 257679 33962
rect 62849 33904 62854 33960
rect 62910 33904 257618 33960
rect 257674 33904 257679 33960
rect 62849 33902 257679 33904
rect 62849 33899 62915 33902
rect 257613 33899 257679 33902
rect 50337 33826 50403 33829
rect 538397 33826 538463 33829
rect 50337 33824 538463 33826
rect 50337 33768 50342 33824
rect 50398 33768 538402 33824
rect 538458 33768 538463 33824
rect 50337 33766 538463 33768
rect 50337 33763 50403 33766
rect 538397 33763 538463 33766
rect 239806 33084 239812 33148
rect 239876 33146 239882 33148
rect 583520 33146 584960 33236
rect 239876 33086 584960 33146
rect 239876 33084 239882 33086
rect 583520 32996 584960 33086
rect 56041 32738 56107 32741
rect 210417 32738 210483 32741
rect 56041 32736 210483 32738
rect 56041 32680 56046 32736
rect 56102 32680 210422 32736
rect 210478 32680 210483 32736
rect 56041 32678 210483 32680
rect 56041 32675 56107 32678
rect 210417 32675 210483 32678
rect 50613 32602 50679 32605
rect 297265 32602 297331 32605
rect 50613 32600 297331 32602
rect -960 32466 480 32556
rect 50613 32544 50618 32600
rect 50674 32544 297270 32600
rect 297326 32544 297331 32600
rect 50613 32542 297331 32544
rect 50613 32539 50679 32542
rect 297265 32539 297331 32542
rect 123569 32466 123635 32469
rect -960 32464 123635 32466
rect -960 32408 123574 32464
rect 123630 32408 123635 32464
rect -960 32406 123635 32408
rect -960 32316 480 32406
rect 123569 32403 123635 32406
rect 72601 31106 72667 31109
rect 261201 31106 261267 31109
rect 72601 31104 261267 31106
rect 72601 31048 72606 31104
rect 72662 31048 261206 31104
rect 261262 31048 261267 31104
rect 72601 31046 261267 31048
rect 72601 31043 72667 31046
rect 261201 31043 261267 31046
rect 49601 30970 49667 30973
rect 541985 30970 542051 30973
rect 49601 30968 542051 30970
rect 49601 30912 49606 30968
rect 49662 30912 541990 30968
rect 542046 30912 542051 30968
rect 49601 30910 542051 30912
rect 49601 30907 49667 30910
rect 541985 30907 542051 30910
rect 83273 29882 83339 29885
rect 264789 29882 264855 29885
rect 83273 29880 264855 29882
rect 83273 29824 83278 29880
rect 83334 29824 264794 29880
rect 264850 29824 264855 29880
rect 83273 29822 264855 29824
rect 83273 29819 83339 29822
rect 264789 29819 264855 29822
rect 50429 29746 50495 29749
rect 284702 29746 284708 29748
rect 50429 29744 284708 29746
rect 50429 29688 50434 29744
rect 50490 29688 284708 29744
rect 50429 29686 284708 29688
rect 50429 29683 50495 29686
rect 284702 29684 284708 29686
rect 284772 29684 284778 29748
rect 50245 29610 50311 29613
rect 545481 29610 545547 29613
rect 50245 29608 545547 29610
rect 50245 29552 50250 29608
rect 50306 29552 545486 29608
rect 545542 29552 545547 29608
rect 50245 29550 545547 29552
rect 50245 29547 50311 29550
rect 545481 29547 545547 29550
rect 76189 28386 76255 28389
rect 262397 28386 262463 28389
rect 76189 28384 262463 28386
rect 76189 28328 76194 28384
rect 76250 28328 262402 28384
rect 262458 28328 262463 28384
rect 76189 28326 262463 28328
rect 76189 28323 76255 28326
rect 262397 28323 262463 28326
rect 49141 28250 49207 28253
rect 552657 28250 552723 28253
rect 49141 28248 552723 28250
rect 49141 28192 49146 28248
rect 49202 28192 552662 28248
rect 552718 28192 552723 28248
rect 49141 28190 552723 28192
rect 49141 28187 49207 28190
rect 552657 28187 552723 28190
rect 69105 27026 69171 27029
rect 260005 27026 260071 27029
rect 69105 27024 260071 27026
rect 69105 26968 69110 27024
rect 69166 26968 260010 27024
rect 260066 26968 260071 27024
rect 69105 26966 260071 26968
rect 69105 26963 69171 26966
rect 260005 26963 260071 26966
rect 50521 26890 50587 26893
rect 559741 26890 559807 26893
rect 50521 26888 559807 26890
rect 50521 26832 50526 26888
rect 50582 26832 559746 26888
rect 559802 26832 559807 26888
rect 50521 26830 559807 26832
rect 50521 26827 50587 26830
rect 559741 26827 559807 26830
rect 65517 25666 65583 25669
rect 258809 25666 258875 25669
rect 65517 25664 258875 25666
rect 65517 25608 65522 25664
rect 65578 25608 258814 25664
rect 258870 25608 258875 25664
rect 65517 25606 258875 25608
rect 65517 25603 65583 25606
rect 258809 25603 258875 25606
rect 47761 25530 47827 25533
rect 562317 25530 562383 25533
rect 47761 25528 562383 25530
rect 47761 25472 47766 25528
rect 47822 25472 562322 25528
rect 562378 25472 562383 25528
rect 47761 25470 562383 25472
rect 47761 25467 47827 25470
rect 562317 25467 562383 25470
rect 58433 24306 58499 24309
rect 256417 24306 256483 24309
rect 58433 24304 256483 24306
rect 58433 24248 58438 24304
rect 58494 24248 256422 24304
rect 256478 24248 256483 24304
rect 58433 24246 256483 24248
rect 58433 24243 58499 24246
rect 256417 24243 256483 24246
rect 47853 24170 47919 24173
rect 566825 24170 566891 24173
rect 47853 24168 566891 24170
rect 47853 24112 47858 24168
rect 47914 24112 566830 24168
rect 566886 24112 566891 24168
rect 47853 24110 566891 24112
rect 47853 24107 47919 24110
rect 566825 24107 566891 24110
rect 51717 22946 51783 22949
rect 252829 22946 252895 22949
rect 51717 22944 252895 22946
rect 51717 22888 51722 22944
rect 51778 22888 252834 22944
rect 252890 22888 252895 22944
rect 51717 22886 252895 22888
rect 51717 22883 51783 22886
rect 252829 22883 252895 22886
rect 71497 22810 71563 22813
rect 285806 22810 285812 22812
rect 71497 22808 285812 22810
rect 71497 22752 71502 22808
rect 71558 22752 285812 22808
rect 71497 22750 285812 22752
rect 71497 22747 71563 22750
rect 285806 22748 285812 22750
rect 285876 22748 285882 22812
rect 48037 22674 48103 22677
rect 570321 22674 570387 22677
rect 48037 22672 570387 22674
rect 48037 22616 48042 22672
rect 48098 22616 570326 22672
rect 570382 22616 570387 22672
rect 48037 22614 570387 22616
rect 48037 22611 48103 22614
rect 570321 22611 570387 22614
rect 80697 21450 80763 21453
rect 396533 21450 396599 21453
rect 80697 21448 396599 21450
rect 80697 21392 80702 21448
rect 80758 21392 396538 21448
rect 396594 21392 396599 21448
rect 80697 21390 396599 21392
rect 80697 21387 80763 21390
rect 396533 21387 396599 21390
rect 47577 21314 47643 21317
rect 573909 21314 573975 21317
rect 47577 21312 573975 21314
rect 47577 21256 47582 21312
rect 47638 21256 573914 21312
rect 573970 21256 573975 21312
rect 47577 21254 573975 21256
rect 47577 21251 47643 21254
rect 573909 21251 573975 21254
rect 8753 20226 8819 20229
rect 142797 20226 142863 20229
rect 8753 20224 142863 20226
rect 8753 20168 8758 20224
rect 8814 20168 142802 20224
rect 142858 20168 142863 20224
rect 8753 20166 142863 20168
rect 8753 20163 8819 20166
rect 142797 20163 142863 20166
rect 63217 20090 63283 20093
rect 206277 20090 206343 20093
rect 63217 20088 206343 20090
rect 63217 20032 63222 20088
rect 63278 20032 206282 20088
rect 206338 20032 206343 20088
rect 63217 20030 206343 20032
rect 63217 20027 63283 20030
rect 206277 20027 206343 20030
rect 55029 19954 55095 19957
rect 290181 19954 290247 19957
rect 55029 19952 290247 19954
rect 55029 19896 55034 19952
rect 55090 19896 290186 19952
rect 290242 19896 290247 19952
rect 55029 19894 290247 19896
rect 55029 19891 55095 19894
rect 290181 19891 290247 19894
rect 298686 19756 298692 19820
rect 298756 19818 298762 19820
rect 583520 19818 584960 19908
rect 298756 19758 584960 19818
rect 298756 19756 298762 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3366 19410 3372 19412
rect -960 19350 3372 19410
rect -960 19260 480 19350
rect 3366 19348 3372 19350
rect 3436 19348 3442 19412
rect 79317 18730 79383 18733
rect 393037 18730 393103 18733
rect 79317 18728 393103 18730
rect 79317 18672 79322 18728
rect 79378 18672 393042 18728
rect 393098 18672 393103 18728
rect 79317 18670 393103 18672
rect 79317 18667 79383 18670
rect 393037 18667 393103 18670
rect 47485 18594 47551 18597
rect 555417 18594 555483 18597
rect 47485 18592 555483 18594
rect 47485 18536 47490 18592
rect 47546 18536 555422 18592
rect 555478 18536 555483 18592
rect 47485 18534 555483 18536
rect 47485 18531 47551 18534
rect 555417 18531 555483 18534
rect 70301 17506 70367 17509
rect 233877 17506 233943 17509
rect 70301 17504 233943 17506
rect 70301 17448 70306 17504
rect 70362 17448 233882 17504
rect 233938 17448 233943 17504
rect 70301 17446 233943 17448
rect 70301 17443 70367 17446
rect 233877 17443 233943 17446
rect 83457 17370 83523 17373
rect 403617 17370 403683 17373
rect 83457 17368 403683 17370
rect 83457 17312 83462 17368
rect 83518 17312 403622 17368
rect 403678 17312 403683 17368
rect 83457 17310 403683 17312
rect 83457 17307 83523 17310
rect 403617 17307 403683 17310
rect 4061 17234 4127 17237
rect 31017 17234 31083 17237
rect 4061 17232 31083 17234
rect 4061 17176 4066 17232
rect 4122 17176 31022 17232
rect 31078 17176 31083 17232
rect 4061 17174 31083 17176
rect 4061 17171 4127 17174
rect 31017 17171 31083 17174
rect 50153 17234 50219 17237
rect 531313 17234 531379 17237
rect 50153 17232 531379 17234
rect 50153 17176 50158 17232
rect 50214 17176 531318 17232
rect 531374 17176 531379 17232
rect 50153 17174 531379 17176
rect 50153 17171 50219 17174
rect 531313 17171 531379 17174
rect 27705 16146 27771 16149
rect 151077 16146 151143 16149
rect 27705 16144 151143 16146
rect 27705 16088 27710 16144
rect 27766 16088 151082 16144
rect 151138 16088 151143 16144
rect 27705 16086 151143 16088
rect 27705 16083 27771 16086
rect 151077 16083 151143 16086
rect 76557 16010 76623 16013
rect 385953 16010 386019 16013
rect 76557 16008 386019 16010
rect 76557 15952 76562 16008
rect 76618 15952 385958 16008
rect 386014 15952 386019 16008
rect 76557 15950 386019 15952
rect 76557 15947 76623 15950
rect 385953 15947 386019 15950
rect 67449 15874 67515 15877
rect 510061 15874 510127 15877
rect 67449 15872 510127 15874
rect 67449 15816 67454 15872
rect 67510 15816 510066 15872
rect 510122 15816 510127 15872
rect 67449 15814 510127 15816
rect 67449 15811 67515 15814
rect 510061 15811 510127 15814
rect 80881 14786 80947 14789
rect 214557 14786 214623 14789
rect 80881 14784 214623 14786
rect 80881 14728 80886 14784
rect 80942 14728 214562 14784
rect 214618 14728 214623 14784
rect 80881 14726 214623 14728
rect 80881 14723 80947 14726
rect 214557 14723 214623 14726
rect 72969 14650 73035 14653
rect 378869 14650 378935 14653
rect 72969 14648 378935 14650
rect 72969 14592 72974 14648
rect 73030 14592 378874 14648
rect 378930 14592 378935 14648
rect 72969 14590 378935 14592
rect 72969 14587 73035 14590
rect 378869 14587 378935 14590
rect 65609 14514 65675 14517
rect 502977 14514 503043 14517
rect 65609 14512 503043 14514
rect 65609 14456 65614 14512
rect 65670 14456 502982 14512
rect 503038 14456 503043 14512
rect 65609 14454 503043 14456
rect 65609 14451 65675 14454
rect 502977 14451 503043 14454
rect 77385 13290 77451 13293
rect 188337 13290 188403 13293
rect 77385 13288 188403 13290
rect 77385 13232 77390 13288
rect 77446 13232 188342 13288
rect 188398 13232 188403 13288
rect 77385 13230 188403 13232
rect 77385 13227 77451 13230
rect 188337 13227 188403 13230
rect 75177 13154 75243 13157
rect 382365 13154 382431 13157
rect 75177 13152 382431 13154
rect 75177 13096 75182 13152
rect 75238 13096 382370 13152
rect 382426 13096 382431 13152
rect 75177 13094 382431 13096
rect 75177 13091 75243 13094
rect 382365 13091 382431 13094
rect 61929 13018 61995 13021
rect 495893 13018 495959 13021
rect 61929 13016 495959 13018
rect 61929 12960 61934 13016
rect 61990 12960 495898 13016
rect 495954 12960 495959 13016
rect 61929 12958 495959 12960
rect 61929 12955 61995 12958
rect 495893 12955 495959 12958
rect 73797 11930 73863 11933
rect 220077 11930 220143 11933
rect 73797 11928 220143 11930
rect 73797 11872 73802 11928
rect 73858 11872 220082 11928
rect 220138 11872 220143 11928
rect 73797 11870 220143 11872
rect 73797 11867 73863 11870
rect 220077 11867 220143 11870
rect 72417 11794 72483 11797
rect 375281 11794 375347 11797
rect 72417 11792 375347 11794
rect 72417 11736 72422 11792
rect 72478 11736 375286 11792
rect 375342 11736 375347 11792
rect 72417 11734 375347 11736
rect 72417 11731 72483 11734
rect 375281 11731 375347 11734
rect 62757 11658 62823 11661
rect 492305 11658 492371 11661
rect 62757 11656 492371 11658
rect 62757 11600 62762 11656
rect 62818 11600 492310 11656
rect 492366 11600 492371 11656
rect 62757 11598 492371 11600
rect 62757 11595 62823 11598
rect 492305 11595 492371 11598
rect 52545 10434 52611 10437
rect 140037 10434 140103 10437
rect 52545 10432 140103 10434
rect 52545 10376 52550 10432
rect 52606 10376 140042 10432
rect 140098 10376 140103 10432
rect 52545 10374 140103 10376
rect 52545 10371 52611 10374
rect 140037 10371 140103 10374
rect 59169 10298 59235 10301
rect 488809 10298 488875 10301
rect 59169 10296 488875 10298
rect 59169 10240 59174 10296
rect 59230 10240 488814 10296
rect 488870 10240 488875 10296
rect 59169 10238 488875 10240
rect 59169 10235 59235 10238
rect 488809 10235 488875 10238
rect 66713 9210 66779 9213
rect 224217 9210 224283 9213
rect 66713 9208 224283 9210
rect 66713 9152 66718 9208
rect 66774 9152 224222 9208
rect 224278 9152 224283 9208
rect 66713 9150 224283 9152
rect 66713 9147 66779 9150
rect 224217 9147 224283 9150
rect 87781 9074 87847 9077
rect 332685 9074 332751 9077
rect 87781 9072 332751 9074
rect 87781 9016 87786 9072
rect 87842 9016 332690 9072
rect 332746 9016 332751 9072
rect 87781 9014 332751 9016
rect 87781 9011 87847 9014
rect 332685 9011 332751 9014
rect 2865 8938 2931 8941
rect 35157 8938 35223 8941
rect 2865 8936 35223 8938
rect 2865 8880 2870 8936
rect 2926 8880 35162 8936
rect 35218 8880 35223 8936
rect 2865 8878 35223 8880
rect 2865 8875 2931 8878
rect 35157 8875 35223 8878
rect 57789 8938 57855 8941
rect 485221 8938 485287 8941
rect 57789 8936 485287 8938
rect 57789 8880 57794 8936
rect 57850 8880 485226 8936
rect 485282 8880 485287 8936
rect 57789 8878 485287 8880
rect 57789 8875 57855 8878
rect 485221 8875 485287 8878
rect 59629 7850 59695 7853
rect 146937 7850 147003 7853
rect 59629 7848 147003 7850
rect 59629 7792 59634 7848
rect 59690 7792 146942 7848
rect 146998 7792 147003 7848
rect 59629 7790 147003 7792
rect 59629 7787 59695 7790
rect 146937 7787 147003 7790
rect 4102 7652 4108 7716
rect 4172 7714 4178 7716
rect 234654 7714 234660 7716
rect 4172 7654 234660 7714
rect 4172 7652 4178 7654
rect 234654 7652 234660 7654
rect 234724 7652 234730 7716
rect 237005 7714 237071 7717
rect 285673 7714 285739 7717
rect 237005 7712 285739 7714
rect 237005 7656 237010 7712
rect 237066 7656 285678 7712
rect 285734 7656 285739 7712
rect 237005 7654 285739 7656
rect 237005 7651 237071 7654
rect 285673 7651 285739 7654
rect 324957 7714 325023 7717
rect 417877 7714 417943 7717
rect 324957 7712 417943 7714
rect 324957 7656 324962 7712
rect 325018 7656 417882 7712
rect 417938 7656 417943 7712
rect 324957 7654 417943 7656
rect 324957 7651 325023 7654
rect 417877 7651 417943 7654
rect 87597 7578 87663 7581
rect 325601 7578 325667 7581
rect 87597 7576 325667 7578
rect 87597 7520 87602 7576
rect 87658 7520 325606 7576
rect 325662 7520 325667 7576
rect 87597 7518 325667 7520
rect 87597 7515 87663 7518
rect 325601 7515 325667 7518
rect 422937 7578 423003 7581
rect 442625 7578 442691 7581
rect 422937 7576 442691 7578
rect 422937 7520 422942 7576
rect 422998 7520 442630 7576
rect 442686 7520 442691 7576
rect 422937 7518 442691 7520
rect 422937 7515 423003 7518
rect 442625 7515 442691 7518
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 4102 6490 4108 6492
rect -960 6430 4108 6490
rect -960 6340 480 6430
rect 4102 6428 4108 6430
rect 4172 6428 4178 6492
rect 79685 6490 79751 6493
rect 263593 6490 263659 6493
rect 79685 6488 263659 6490
rect 79685 6432 79690 6488
rect 79746 6432 263598 6488
rect 263654 6432 263659 6488
rect 583520 6476 584960 6566
rect 79685 6430 263659 6432
rect 79685 6427 79751 6430
rect 263593 6427 263659 6430
rect 31293 6354 31359 6357
rect 238109 6354 238175 6357
rect 31293 6352 238175 6354
rect 31293 6296 31298 6352
rect 31354 6296 238114 6352
rect 238170 6296 238175 6352
rect 31293 6294 238175 6296
rect 31293 6291 31359 6294
rect 238109 6291 238175 6294
rect 12341 6218 12407 6221
rect 242065 6218 242131 6221
rect 12341 6216 242131 6218
rect 12341 6160 12346 6216
rect 12402 6160 242070 6216
rect 242126 6160 242131 6216
rect 12341 6158 242131 6160
rect 12341 6155 12407 6158
rect 242065 6155 242131 6158
rect 266997 6218 267063 6221
rect 283097 6218 283163 6221
rect 266997 6216 283163 6218
rect 266997 6160 267002 6216
rect 267058 6160 283102 6216
rect 283158 6160 283163 6216
rect 266997 6158 283163 6160
rect 266997 6155 267063 6158
rect 283097 6155 283163 6158
rect 278037 5674 278103 5677
rect 286593 5674 286659 5677
rect 278037 5672 286659 5674
rect 278037 5616 278042 5672
rect 278098 5616 286598 5672
rect 286654 5616 286659 5672
rect 278037 5614 286659 5616
rect 278037 5611 278103 5614
rect 286593 5611 286659 5614
rect 1669 5266 1735 5269
rect 85573 5266 85639 5269
rect 1669 5264 85639 5266
rect 1669 5208 1674 5264
rect 1730 5208 85578 5264
rect 85634 5208 85639 5264
rect 1669 5206 85639 5208
rect 1669 5203 1735 5206
rect 85573 5203 85639 5206
rect 48957 5130 49023 5133
rect 197997 5130 198063 5133
rect 48957 5128 198063 5130
rect 48957 5072 48962 5128
rect 49018 5072 198002 5128
rect 198058 5072 198063 5128
rect 48957 5070 198063 5072
rect 48957 5067 49023 5070
rect 197997 5067 198063 5070
rect 78581 4994 78647 4997
rect 287053 4994 287119 4997
rect 78581 4992 287119 4994
rect 78581 4936 78586 4992
rect 78642 4936 287058 4992
rect 287114 4936 287119 4992
rect 78581 4934 287119 4936
rect 78581 4931 78647 4934
rect 287053 4931 287119 4934
rect 431217 4994 431283 4997
rect 435541 4994 435607 4997
rect 431217 4992 435607 4994
rect 431217 4936 431222 4992
rect 431278 4936 435546 4992
rect 435602 4936 435607 4992
rect 431217 4934 435607 4936
rect 431217 4931 431283 4934
rect 435541 4931 435607 4934
rect 71037 4858 71103 4861
rect 279509 4858 279575 4861
rect 71037 4856 279575 4858
rect 71037 4800 71042 4856
rect 71098 4800 279514 4856
rect 279570 4800 279575 4856
rect 71037 4798 279575 4800
rect 71037 4795 71103 4798
rect 279509 4795 279575 4798
rect 287697 4858 287763 4861
rect 410793 4858 410859 4861
rect 287697 4856 410859 4858
rect 287697 4800 287702 4856
rect 287758 4800 410798 4856
rect 410854 4800 410859 4856
rect 287697 4798 410859 4800
rect 287697 4795 287763 4798
rect 410793 4795 410859 4798
rect 411897 4858 411963 4861
rect 414289 4858 414355 4861
rect 411897 4856 414355 4858
rect 411897 4800 411902 4856
rect 411958 4800 414294 4856
rect 414350 4800 414355 4856
rect 411897 4798 414355 4800
rect 411897 4795 411963 4798
rect 414289 4795 414355 4798
rect 418797 4858 418863 4861
rect 424961 4858 425027 4861
rect 418797 4856 425027 4858
rect 418797 4800 418802 4856
rect 418858 4800 424966 4856
rect 425022 4800 425027 4856
rect 418797 4798 425027 4800
rect 418797 4795 418863 4798
rect 424961 4795 425027 4798
rect 429837 4858 429903 4861
rect 432045 4858 432111 4861
rect 429837 4856 432111 4858
rect 429837 4800 429842 4856
rect 429898 4800 432050 4856
rect 432106 4800 432111 4856
rect 429837 4798 432111 4800
rect 429837 4795 429903 4798
rect 432045 4795 432111 4798
rect 450537 4858 450603 4861
rect 453297 4858 453363 4861
rect 450537 4856 453363 4858
rect 450537 4800 450542 4856
rect 450598 4800 453302 4856
rect 453358 4800 453363 4856
rect 450537 4798 453363 4800
rect 450537 4795 450603 4798
rect 453297 4795 453363 4798
rect 425697 4178 425763 4181
rect 428457 4178 428523 4181
rect 425697 4176 428523 4178
rect 425697 4120 425702 4176
rect 425758 4120 428462 4176
rect 428518 4120 428523 4176
rect 425697 4118 428523 4120
rect 425697 4115 425763 4118
rect 428457 4115 428523 4118
rect 436737 4178 436803 4181
rect 439129 4178 439195 4181
rect 436737 4176 439195 4178
rect 436737 4120 436742 4176
rect 436798 4120 439134 4176
rect 439190 4120 439195 4176
rect 436737 4118 439195 4120
rect 436737 4115 436803 4118
rect 439129 4115 439195 4118
rect 443637 4178 443703 4181
rect 446213 4178 446279 4181
rect 443637 4176 446279 4178
rect 443637 4120 443642 4176
rect 443698 4120 446218 4176
rect 446274 4120 446279 4176
rect 443637 4118 446279 4120
rect 443637 4115 443703 4118
rect 446213 4115 446279 4118
rect 447777 4178 447843 4181
rect 449801 4178 449867 4181
rect 447777 4176 449867 4178
rect 447777 4120 447782 4176
rect 447838 4120 449806 4176
rect 449862 4120 449867 4176
rect 447777 4118 449867 4120
rect 447777 4115 447843 4118
rect 449801 4115 449867 4118
rect 54937 4042 55003 4045
rect 55857 4042 55923 4045
rect 54937 4040 55923 4042
rect 54937 3984 54942 4040
rect 54998 3984 55862 4040
rect 55918 3984 55923 4040
rect 54937 3982 55923 3984
rect 54937 3979 55003 3982
rect 55857 3979 55923 3982
rect 258257 4042 258323 4045
rect 282913 4042 282979 4045
rect 258257 4040 282979 4042
rect 258257 3984 258262 4040
rect 258318 3984 282918 4040
rect 282974 3984 282979 4040
rect 258257 3982 282979 3984
rect 258257 3979 258323 3982
rect 282913 3979 282979 3982
rect 439497 4042 439563 4045
rect 442901 4042 442967 4045
rect 439497 4040 442967 4042
rect 439497 3984 439502 4040
rect 439558 3984 442906 4040
rect 442962 3984 442967 4040
rect 439497 3982 442967 3984
rect 439497 3979 439563 3982
rect 442901 3979 442967 3982
rect 576117 4042 576183 4045
rect 577405 4042 577471 4045
rect 576117 4040 577471 4042
rect 576117 3984 576122 4040
rect 576178 3984 577410 4040
rect 577466 3984 577471 4040
rect 576117 3982 577471 3984
rect 576117 3979 576183 3982
rect 577405 3979 577471 3982
rect 109309 3906 109375 3909
rect 126421 3906 126487 3909
rect 109309 3904 126487 3906
rect 109309 3848 109314 3904
rect 109370 3848 126426 3904
rect 126482 3848 126487 3904
rect 109309 3846 126487 3848
rect 109309 3843 109375 3846
rect 126421 3843 126487 3846
rect 229829 3906 229895 3909
rect 247677 3906 247743 3909
rect 229829 3904 247743 3906
rect 229829 3848 229834 3904
rect 229890 3848 247682 3904
rect 247738 3848 247743 3904
rect 229829 3846 247743 3848
rect 229829 3843 229895 3846
rect 247677 3843 247743 3846
rect 254669 3906 254735 3909
rect 280797 3906 280863 3909
rect 254669 3904 280863 3906
rect 254669 3848 254674 3904
rect 254730 3848 280802 3904
rect 280858 3848 280863 3904
rect 254669 3846 280863 3848
rect 254669 3843 254735 3846
rect 280797 3843 280863 3846
rect 421557 3906 421623 3909
rect 463969 3906 464035 3909
rect 421557 3904 464035 3906
rect 421557 3848 421562 3904
rect 421618 3848 463974 3904
rect 464030 3848 464035 3904
rect 421557 3846 464035 3848
rect 421557 3843 421623 3846
rect 463969 3843 464035 3846
rect 105721 3770 105787 3773
rect 126237 3770 126303 3773
rect 105721 3768 126303 3770
rect 105721 3712 105726 3768
rect 105782 3712 126242 3768
rect 126298 3712 126303 3768
rect 105721 3710 126303 3712
rect 105721 3707 105787 3710
rect 126237 3707 126303 3710
rect 247585 3770 247651 3773
rect 280981 3770 281047 3773
rect 247585 3768 281047 3770
rect 247585 3712 247590 3768
rect 247646 3712 280986 3768
rect 281042 3712 281047 3768
rect 247585 3710 281047 3712
rect 247585 3707 247651 3710
rect 280981 3707 281047 3710
rect 428549 3770 428615 3773
rect 471053 3770 471119 3773
rect 428549 3768 471119 3770
rect 428549 3712 428554 3768
rect 428610 3712 471058 3768
rect 471114 3712 471119 3768
rect 428549 3710 471119 3712
rect 428549 3707 428615 3710
rect 471053 3707 471119 3710
rect 64321 3634 64387 3637
rect 90449 3634 90515 3637
rect 64321 3632 90515 3634
rect 64321 3576 64326 3632
rect 64382 3576 90454 3632
rect 90510 3576 90515 3632
rect 64321 3574 90515 3576
rect 64321 3571 64387 3574
rect 90449 3571 90515 3574
rect 92749 3634 92815 3637
rect 97257 3634 97323 3637
rect 92749 3632 97323 3634
rect 92749 3576 92754 3632
rect 92810 3576 97262 3632
rect 97318 3576 97323 3632
rect 92749 3574 97323 3576
rect 92749 3571 92815 3574
rect 97257 3571 97323 3574
rect 102225 3634 102291 3637
rect 126605 3634 126671 3637
rect 102225 3632 126671 3634
rect 102225 3576 102230 3632
rect 102286 3576 126610 3632
rect 126666 3576 126671 3632
rect 102225 3574 126671 3576
rect 102225 3571 102291 3574
rect 126605 3571 126671 3574
rect 169569 3634 169635 3637
rect 170397 3634 170463 3637
rect 169569 3632 170463 3634
rect 169569 3576 169574 3632
rect 169630 3576 170402 3632
rect 170458 3576 170463 3632
rect 169569 3574 170463 3576
rect 169569 3571 169635 3574
rect 170397 3571 170463 3574
rect 194409 3634 194475 3637
rect 195237 3634 195303 3637
rect 194409 3632 195303 3634
rect 194409 3576 194414 3632
rect 194470 3576 195242 3632
rect 195298 3576 195303 3632
rect 194409 3574 195303 3576
rect 194409 3571 194475 3574
rect 195237 3571 195303 3574
rect 244089 3634 244155 3637
rect 271137 3634 271203 3637
rect 272425 3634 272491 3637
rect 244089 3632 270970 3634
rect 244089 3576 244094 3632
rect 244150 3576 270970 3632
rect 244089 3574 270970 3576
rect 244089 3571 244155 3574
rect 7649 3498 7715 3501
rect 11697 3498 11763 3501
rect 7649 3496 11763 3498
rect 7649 3440 7654 3496
rect 7710 3440 11702 3496
rect 11758 3440 11763 3496
rect 7649 3438 11763 3440
rect 7649 3435 7715 3438
rect 11697 3435 11763 3438
rect 17033 3498 17099 3501
rect 18597 3498 18663 3501
rect 17033 3496 18663 3498
rect 17033 3440 17038 3496
rect 17094 3440 18602 3496
rect 18658 3440 18663 3496
rect 17033 3438 18663 3440
rect 17033 3435 17099 3438
rect 18597 3435 18663 3438
rect 47853 3498 47919 3501
rect 51717 3498 51783 3501
rect 47853 3496 51783 3498
rect 47853 3440 47858 3496
rect 47914 3440 51722 3496
rect 51778 3440 51783 3496
rect 47853 3438 51783 3440
rect 47853 3435 47919 3438
rect 51717 3435 51783 3438
rect 62021 3498 62087 3501
rect 62849 3498 62915 3501
rect 102777 3498 102843 3501
rect 62021 3496 62915 3498
rect 62021 3440 62026 3496
rect 62082 3440 62854 3496
rect 62910 3440 62915 3496
rect 62021 3438 62915 3440
rect 62021 3435 62087 3438
rect 62849 3435 62915 3438
rect 62990 3496 102843 3498
rect 62990 3440 102782 3496
rect 102838 3440 102843 3496
rect 62990 3438 102843 3440
rect 60825 3362 60891 3365
rect 62990 3362 63050 3438
rect 102777 3435 102843 3438
rect 103329 3498 103395 3501
rect 270585 3498 270651 3501
rect 103329 3496 270651 3498
rect 103329 3440 103334 3496
rect 103390 3440 270590 3496
rect 270646 3440 270651 3496
rect 103329 3438 270651 3440
rect 103329 3435 103395 3438
rect 270585 3435 270651 3438
rect 270910 3362 270970 3574
rect 271137 3632 272491 3634
rect 271137 3576 271142 3632
rect 271198 3576 272430 3632
rect 272486 3576 272491 3632
rect 271137 3574 272491 3576
rect 271137 3571 271203 3574
rect 272425 3571 272491 3574
rect 284937 3634 285003 3637
rect 293677 3634 293743 3637
rect 284937 3632 293743 3634
rect 284937 3576 284942 3632
rect 284998 3576 293682 3632
rect 293738 3576 293743 3632
rect 284937 3574 293743 3576
rect 284937 3571 285003 3574
rect 293677 3571 293743 3574
rect 435357 3634 435423 3637
rect 478137 3634 478203 3637
rect 435357 3632 478203 3634
rect 435357 3576 435362 3632
rect 435418 3576 478142 3632
rect 478198 3576 478203 3632
rect 435357 3574 478203 3576
rect 435357 3571 435423 3574
rect 478137 3571 478203 3574
rect 271045 3498 271111 3501
rect 283281 3498 283347 3501
rect 271045 3496 283347 3498
rect 271045 3440 271050 3496
rect 271106 3440 283286 3496
rect 283342 3440 283347 3496
rect 271045 3438 283347 3440
rect 271045 3435 271111 3438
rect 283281 3435 283347 3438
rect 289077 3498 289143 3501
rect 300761 3498 300827 3501
rect 289077 3496 300827 3498
rect 289077 3440 289082 3496
rect 289138 3440 300766 3496
rect 300822 3440 300827 3496
rect 289077 3438 300827 3440
rect 289077 3435 289143 3438
rect 300761 3435 300827 3438
rect 417417 3498 417483 3501
rect 460381 3498 460447 3501
rect 417417 3496 460447 3498
rect 417417 3440 417422 3496
rect 417478 3440 460386 3496
rect 460442 3440 460447 3496
rect 417417 3438 460447 3440
rect 417417 3435 417483 3438
rect 460381 3435 460447 3438
rect 512637 3498 512703 3501
rect 513557 3498 513623 3501
rect 512637 3496 513623 3498
rect 512637 3440 512642 3496
rect 512698 3440 513562 3496
rect 513618 3440 513623 3496
rect 512637 3438 513623 3440
rect 512637 3435 512703 3438
rect 513557 3435 513623 3438
rect 562317 3498 562383 3501
rect 563237 3498 563303 3501
rect 562317 3496 563303 3498
rect 562317 3440 562322 3496
rect 562378 3440 563242 3496
rect 563298 3440 563303 3496
rect 562317 3438 563303 3440
rect 562317 3435 562383 3438
rect 563237 3435 563303 3438
rect 279417 3362 279483 3365
rect 60825 3360 63050 3362
rect 60825 3304 60830 3360
rect 60886 3304 63050 3360
rect 60825 3302 63050 3304
rect 64830 3302 258090 3362
rect 270910 3360 279483 3362
rect 270910 3304 279422 3360
rect 279478 3304 279483 3360
rect 270910 3302 279483 3304
rect 60825 3299 60891 3302
rect 57237 3226 57303 3229
rect 64830 3226 64890 3302
rect 57237 3224 64890 3226
rect 57237 3168 57242 3224
rect 57298 3168 64890 3224
rect 57237 3166 64890 3168
rect 258030 3226 258090 3302
rect 279417 3299 279483 3302
rect 282177 3362 282243 3365
rect 339861 3362 339927 3365
rect 282177 3360 339927 3362
rect 282177 3304 282182 3360
rect 282238 3304 339866 3360
rect 339922 3304 339927 3360
rect 282177 3302 339927 3304
rect 282177 3299 282243 3302
rect 339861 3299 339927 3302
rect 442257 3362 442323 3365
rect 582189 3362 582255 3365
rect 442257 3360 582255 3362
rect 442257 3304 442262 3360
rect 442318 3304 582194 3360
rect 582250 3304 582255 3360
rect 442257 3302 582255 3304
rect 442257 3299 442323 3302
rect 582189 3299 582255 3302
rect 280061 3226 280127 3229
rect 258030 3224 280127 3226
rect 258030 3168 280066 3224
rect 280122 3168 280127 3224
rect 258030 3166 280127 3168
rect 57237 3163 57303 3166
rect 280061 3163 280127 3166
rect 432597 3226 432663 3229
rect 474549 3226 474615 3229
rect 432597 3224 474615 3226
rect 432597 3168 432602 3224
rect 432658 3168 474554 3224
rect 474610 3168 474615 3224
rect 432597 3166 474615 3168
rect 432597 3163 432663 3166
rect 474549 3163 474615 3166
rect 414657 3090 414723 3093
rect 456885 3090 456951 3093
rect 414657 3088 456951 3090
rect 414657 3032 414662 3088
rect 414718 3032 456890 3088
rect 456946 3032 456951 3088
rect 414657 3030 456951 3032
rect 414657 3027 414723 3030
rect 456885 3027 456951 3030
rect 19425 2818 19491 2821
rect 271781 2818 271847 2821
rect 19425 2816 271847 2818
rect 19425 2760 19430 2816
rect 19486 2760 271786 2816
rect 271842 2760 271847 2816
rect 19425 2758 271847 2760
rect 19425 2755 19491 2758
rect 271781 2755 271847 2758
<< via3 >>
rect 558132 683844 558196 683908
rect 30420 671196 30484 671260
rect 15700 658140 15764 658204
rect 179276 655012 179340 655076
rect 450492 655012 450556 655076
rect 175044 653108 175108 653172
rect 480300 653108 480364 653172
rect 176516 649980 176580 650044
rect 476620 649980 476684 650044
rect 550772 649844 550836 649908
rect 44036 648212 44100 648276
rect 377628 648212 377692 648276
rect 176332 647260 176396 647324
rect 547644 647260 547708 647324
rect 176148 645900 176212 645964
rect 54892 645356 54956 645420
rect 296852 645356 296916 645420
rect 48636 643588 48700 643652
rect 297036 643588 297100 643652
rect 46796 643316 46860 643380
rect 550036 643044 550100 643108
rect 177068 641684 177132 641748
rect 294828 641140 294892 641204
rect 479380 641140 479444 641204
rect 177252 640324 177316 640388
rect 177804 640324 177868 640388
rect 297036 640188 297100 640252
rect 47900 639644 47964 639708
rect 296852 639644 296916 639708
rect 31524 639372 31588 639436
rect 291884 639372 291948 639436
rect 294644 639372 294708 639436
rect 478092 639372 478156 639436
rect 294460 638012 294524 638076
rect 482140 638012 482204 638076
rect 34284 637876 34348 637940
rect 291700 637876 291764 637940
rect 292068 637876 292132 637940
rect 483612 637876 483676 637940
rect 177436 637604 177500 637668
rect 32996 637196 33060 637260
rect 178908 637060 178972 637124
rect 48084 636652 48148 636716
rect 48452 636516 48516 636580
rect 179092 636380 179156 636444
rect 55996 635836 56060 635900
rect 377812 635836 377876 635900
rect 296668 635428 296732 635492
rect 47716 635292 47780 635356
rect 296484 635292 296548 635356
rect 127572 634068 127636 634132
rect 249012 634068 249076 634132
rect 127572 633660 127636 633724
rect 249012 633660 249076 633724
rect 179276 632164 179340 632228
rect 179092 631076 179156 631140
rect 555372 630804 555436 630868
rect 178908 628900 178972 628964
rect 57652 628764 57716 628828
rect 57836 627676 57900 627740
rect 58940 626588 59004 626652
rect 291148 626452 291212 626516
rect 377628 626452 377692 626516
rect 176148 625636 176212 625700
rect 296852 625636 296916 625700
rect 177252 624548 177316 624612
rect 297036 624548 297100 624612
rect 294828 624004 294892 624068
rect 550772 624004 550836 624068
rect 294644 623188 294708 623252
rect 177620 622372 177684 622436
rect 288388 622372 288452 622436
rect 292068 621556 292132 621620
rect 177068 621284 177132 621348
rect 543780 621284 543844 621348
rect 294460 620740 294524 620804
rect 59124 620196 59188 620260
rect 177252 620196 177316 620260
rect 298140 619924 298204 619988
rect 546540 619924 546604 619988
rect 29132 619108 29196 619172
rect 58756 619108 58820 619172
rect 175044 619108 175108 619172
rect 290596 619108 290660 619172
rect 550956 618564 551020 618628
rect 172652 618292 172716 618356
rect 295380 618292 295444 618356
rect 177436 618020 177500 618084
rect 175228 617476 175292 617540
rect 287100 617476 287164 617540
rect 176332 616932 176396 616996
rect 173940 616660 174004 616724
rect 295932 616660 295996 616724
rect 176516 615844 176580 615908
rect 282132 615844 282196 615908
rect 291884 615844 291948 615908
rect 288572 615028 288636 615092
rect 377812 615028 377876 615092
rect 177804 614756 177868 614820
rect 291700 614756 291764 614820
rect 541020 614484 541084 614548
rect 294828 614212 294892 614276
rect 177436 613668 177500 613732
rect 280660 613396 280724 613460
rect 542860 613124 542924 613188
rect 177068 612580 177132 612644
rect 294460 612580 294524 612644
rect 284892 611764 284956 611828
rect 541204 611764 541268 611828
rect 177804 611492 177868 611556
rect 177620 611356 177684 611420
rect 256740 610948 256804 611012
rect 177252 610676 177316 610740
rect 59676 610404 59740 610468
rect 177988 610404 178052 610468
rect 286180 610404 286244 610468
rect 543412 610404 543476 610468
rect 298324 610132 298388 610196
rect 177436 609724 177500 609788
rect 176700 609316 176764 609380
rect 294644 609316 294708 609380
rect 178172 609044 178236 609108
rect 177804 608500 177868 608564
rect 290780 608500 290844 608564
rect 177252 608228 177316 608292
rect 299612 607684 299676 607748
rect 543044 607684 543108 607748
rect 177068 607140 177132 607204
rect 177804 607140 177868 607204
rect 296668 607140 296732 607204
rect 177988 607004 178052 607068
rect 298508 606868 298572 606932
rect 543228 606324 543292 606388
rect 26740 606052 26804 606116
rect 177068 606052 177132 606116
rect 292620 606052 292684 606116
rect 299428 605236 299492 605300
rect 177620 604964 177684 605028
rect 297036 604964 297100 605028
rect 539364 604964 539428 605028
rect 176700 604420 176764 604484
rect 299244 604420 299308 604484
rect 299612 604420 299676 604484
rect 166764 603876 166828 603940
rect 287652 603604 287716 603668
rect 539548 603604 539612 603668
rect 177436 602788 177500 602852
rect 298692 602924 298756 602988
rect 299428 602924 299492 602988
rect 255268 602516 255332 602580
rect 299428 601972 299492 602036
rect 298140 601836 298204 601900
rect 177252 601700 177316 601764
rect 538260 601700 538324 601764
rect 295012 601156 295076 601220
rect 294828 601020 294892 601084
rect 295748 600340 295812 600404
rect 538812 600340 538876 600404
rect 539548 600340 539612 600404
rect 500172 599660 500236 599724
rect 296300 599388 296364 599452
rect 256740 598844 256804 598908
rect 256924 598708 256988 598772
rect 504220 598028 504284 598092
rect 256740 597892 256804 597956
rect 506980 598028 507044 598092
rect 533292 598028 533356 598092
rect 534580 598028 534644 598092
rect 295380 597484 295444 597548
rect 299428 597484 299492 597548
rect 296116 597076 296180 597140
rect 178540 596396 178604 596460
rect 299796 596396 299860 596460
rect 295748 596260 295812 596324
rect 296300 596260 296364 596324
rect 296668 596124 296732 596188
rect 299060 595444 299124 595508
rect 298324 594764 298388 594828
rect 291700 594628 291764 594692
rect 283972 593812 284036 593876
rect 298876 592860 298940 592924
rect 281028 592180 281092 592244
rect 298508 592044 298572 592108
rect 285260 591364 285324 591428
rect 580212 590956 580276 591020
rect 294460 590548 294524 590612
rect 294828 590276 294892 590340
rect 283788 589596 283852 589660
rect 294644 589188 294708 589252
rect 294460 588916 294524 588980
rect 289308 588100 289372 588164
rect 294644 587284 294708 587348
rect 178724 586740 178788 586804
rect 287836 586468 287900 586532
rect 295012 586528 295076 586532
rect 295012 586472 295026 586528
rect 295026 586472 295076 586528
rect 295012 586468 295076 586472
rect 290964 585652 291028 585716
rect 290596 585108 290660 585172
rect 288204 584836 288268 584900
rect 286364 584020 286428 584084
rect 285076 583204 285140 583268
rect 283420 582388 283484 582452
rect 283604 581572 283668 581636
rect 290964 581088 291028 581092
rect 290964 581032 290978 581088
rect 290978 581032 291028 581088
rect 290964 581028 291028 581032
rect 290780 580892 290844 580956
rect 290964 580756 291028 580820
rect 289492 579804 289556 579868
rect 293172 579124 293236 579188
rect 290596 578308 290660 578372
rect 287100 578172 287164 578236
rect 551140 577628 551204 577692
rect 288020 577492 288084 577556
rect 379468 577492 379532 577556
rect 296668 577356 296732 577420
rect 292068 576676 292132 576740
rect 296668 576676 296732 576740
rect 257108 575860 257172 575924
rect 256924 575452 256988 575516
rect 291884 575044 291948 575108
rect 285444 574228 285508 574292
rect 382228 574228 382292 574292
rect 256740 572732 256804 572796
rect 257108 572596 257172 572660
rect 257108 571780 257172 571844
rect 166580 571236 166644 571300
rect 286548 571236 286612 571300
rect 299244 571100 299308 571164
rect 256924 570964 256988 571028
rect 171548 570012 171612 570076
rect 299244 570012 299308 570076
rect 177252 569876 177316 569940
rect 294828 569936 294892 569940
rect 294828 569880 294878 569936
rect 294878 569880 294892 569936
rect 294828 569876 294892 569880
rect 295012 569332 295076 569396
rect 177252 569060 177316 569124
rect 292620 568516 292684 568580
rect 292988 568244 293052 568308
rect 175044 567972 175108 568036
rect 296668 567428 296732 567492
rect 296668 567020 296732 567084
rect 2820 566884 2884 566948
rect 179828 566816 179892 566880
rect 179460 565796 179524 565860
rect 176516 564708 176580 564772
rect 289124 564708 289188 564772
rect 288388 564436 288452 564500
rect 288940 563620 289004 563684
rect 179828 563076 179892 563140
rect 288572 563076 288636 563140
rect 292252 562532 292316 562596
rect 180380 562464 180444 562528
rect 291148 562260 291212 562324
rect 172652 561580 172716 561644
rect 180564 561376 180628 561440
rect 255820 560628 255884 560692
rect 177988 560356 178052 560420
rect 57652 560280 57716 560284
rect 57652 560224 57666 560280
rect 57666 560224 57716 560280
rect 57652 560220 57716 560224
rect 59124 560220 59188 560284
rect 166764 560280 166828 560284
rect 166764 560224 166814 560280
rect 166814 560224 166828 560280
rect 166764 560220 166828 560224
rect 175228 560220 175292 560284
rect 255084 560492 255148 560556
rect 58756 559404 58820 559468
rect 59860 558996 59924 559060
rect 512132 558996 512196 559060
rect 173940 558860 174004 558924
rect 180564 558920 180628 558924
rect 180564 558864 180614 558920
rect 180614 558864 180628 558920
rect 180564 558860 180628 558864
rect 180380 558724 180444 558788
rect 295012 558452 295076 558516
rect 523172 558452 523236 558516
rect 256924 558180 256988 558244
rect 515260 558180 515324 558244
rect 296668 557772 296732 557836
rect 53604 557636 53668 557700
rect 32812 557500 32876 557564
rect 294644 557364 294708 557428
rect 499068 557364 499132 557428
rect 296668 557228 296732 557292
rect 299060 557228 299124 557292
rect 505140 557228 505204 557292
rect 289308 557092 289372 557156
rect 525380 557092 525444 557156
rect 178724 556548 178788 556612
rect 47532 556140 47596 556204
rect 288388 556140 288452 556204
rect 35756 554916 35820 554980
rect 55812 554916 55876 554980
rect 30972 554780 31036 554844
rect 507900 554840 507964 554844
rect 507900 554784 507914 554840
rect 507914 554784 507964 554840
rect 507900 554780 507964 554784
rect 522988 554840 523052 554844
rect 522988 554784 523038 554840
rect 523038 554784 523052 554840
rect 522988 554780 523052 554784
rect 177252 554644 177316 554708
rect 58572 554372 58636 554436
rect 33916 554236 33980 554300
rect 54524 554100 54588 554164
rect 178540 554100 178604 554164
rect 18460 553828 18524 553892
rect 35572 553828 35636 553892
rect 40724 553556 40788 553620
rect 39804 553420 39868 553484
rect 30052 552196 30116 552260
rect 291148 551652 291212 551716
rect 59676 551516 59740 551580
rect 292068 551516 292132 551580
rect 539548 551652 539612 551716
rect 179460 551380 179524 551444
rect 59124 550836 59188 550900
rect 32444 550700 32508 550764
rect 509188 550760 509252 550764
rect 509188 550704 509238 550760
rect 509238 550704 509252 550760
rect 509188 550700 509252 550704
rect 296484 550564 296548 550628
rect 502380 550564 502444 550628
rect 296484 550216 296548 550220
rect 296484 550160 296534 550216
rect 296534 550160 296548 550216
rect 296484 550156 296548 550160
rect 298876 550020 298940 550084
rect 511028 550020 511092 550084
rect 176516 549808 176580 549812
rect 176516 549752 176566 549808
rect 176566 549752 176580 549808
rect 176516 549748 176580 549752
rect 36860 549340 36924 549404
rect 288572 549068 288636 549132
rect 290964 549068 291028 549132
rect 514156 549068 514220 549132
rect 289492 548932 289556 548996
rect 529060 548932 529124 548996
rect 30236 548388 30300 548452
rect 506612 547844 506676 547908
rect 283972 547572 284036 547636
rect 498700 547572 498764 547636
rect 37044 547436 37108 547500
rect 292252 547436 292316 547500
rect 293172 547436 293236 547500
rect 519308 547436 519372 547500
rect 175044 547164 175108 547228
rect 29868 546484 29932 546548
rect 282868 546484 282932 546548
rect 292620 546484 292684 546548
rect 503668 546544 503732 546548
rect 503668 546488 503718 546544
rect 503718 546488 503732 546544
rect 503668 546484 503732 546488
rect 255084 546348 255148 546412
rect 284892 546212 284956 546276
rect 508268 546212 508332 546276
rect 34100 546076 34164 546140
rect 286548 546076 286612 546140
rect 288204 546076 288268 546140
rect 497412 546076 497476 546140
rect 27476 545668 27540 545732
rect 382228 545668 382292 545732
rect 296300 544988 296364 545052
rect 502564 544988 502628 545052
rect 28764 543764 28828 543828
rect 292988 543356 293052 543420
rect 516180 543356 516244 543420
rect 296668 542404 296732 542468
rect 29132 542268 29196 542332
rect 58388 542132 58452 542196
rect 296300 542268 296364 542332
rect 285260 541996 285324 542060
rect 532740 541996 532804 542060
rect 32628 541860 32692 541924
rect 288572 541860 288636 541924
rect 294460 541860 294524 541924
rect 539732 541860 539796 541924
rect 171548 541724 171612 541788
rect 29684 541044 29748 541108
rect 506796 541044 506860 541108
rect 295932 540908 295996 540972
rect 502932 540908 502996 540972
rect 510660 540636 510724 540700
rect 521700 539744 521764 539748
rect 521700 539688 521714 539744
rect 521714 539688 521764 539744
rect 521700 539684 521764 539688
rect 33732 539548 33796 539612
rect 521884 539548 521948 539612
rect 282132 539140 282196 539204
rect 514340 539140 514404 539204
rect 58940 538052 59004 538116
rect 283788 537780 283852 537844
rect 534028 537780 534092 537844
rect 580396 537780 580460 537844
rect 31340 537644 31404 537708
rect 286180 537644 286244 537708
rect 290596 537644 290660 537708
rect 520412 537644 520476 537708
rect 166580 537508 166644 537572
rect 35388 537372 35452 537436
rect 379468 537372 379532 537436
rect 298692 536556 298756 536620
rect 518388 536556 518452 536620
rect 299244 536420 299308 536484
rect 526116 536420 526180 536484
rect 291700 536284 291764 536348
rect 519492 536284 519556 536348
rect 58756 535740 58820 535804
rect 535500 535468 535564 535532
rect 255820 534924 255884 534988
rect 57836 534788 57900 534852
rect 499620 534168 499684 534172
rect 499620 534112 499634 534168
rect 499634 534112 499684 534168
rect 499620 534108 499684 534112
rect 287652 533700 287716 533764
rect 498884 533700 498948 533764
rect 510476 532748 510540 532812
rect 514708 532808 514772 532812
rect 514708 532752 514758 532808
rect 514758 532752 514772 532808
rect 514708 532748 514772 532752
rect 518940 532808 519004 532812
rect 518940 532752 518990 532808
rect 518990 532752 519004 532808
rect 518940 532748 519004 532752
rect 177436 532612 177500 532676
rect 52316 531796 52380 531860
rect 296852 531796 296916 531860
rect 499804 531388 499868 531452
rect 522068 531388 522132 531452
rect 525748 531448 525812 531452
rect 525748 531392 525798 531448
rect 525798 531392 525812 531448
rect 525748 531388 525812 531392
rect 529980 531388 530044 531452
rect 61884 530436 61948 530500
rect 50844 530300 50908 530364
rect 43852 530164 43916 530228
rect 36676 529892 36740 529956
rect 53788 529816 53852 529820
rect 53788 529760 53802 529816
rect 53802 529760 53852 529816
rect 53788 529756 53852 529760
rect 286364 529484 286428 529548
rect 497596 529484 497660 529548
rect 61332 529348 61396 529412
rect 501276 529212 501340 529276
rect 450492 529076 450556 529140
rect 42564 528532 42628 528596
rect 501644 528532 501708 528596
rect 26004 528124 26068 528188
rect 476620 527988 476684 528052
rect 536788 527988 536852 528052
rect 49740 527172 49804 527236
rect 55076 527232 55140 527236
rect 55076 527176 55126 527232
rect 55126 527176 55140 527232
rect 55076 527172 55140 527176
rect 511948 527232 512012 527236
rect 511948 527176 511998 527232
rect 511998 527176 512012 527232
rect 511948 527172 512012 527176
rect 514892 527172 514956 527236
rect 518020 527172 518084 527236
rect 523540 527172 523604 527236
rect 44956 526764 45020 526828
rect 291148 526764 291212 526828
rect 288020 526628 288084 526692
rect 512316 526900 512380 526964
rect 296116 526764 296180 526828
rect 502748 526764 502812 526828
rect 501460 526492 501524 526556
rect 257108 526084 257172 526148
rect 514524 526084 514588 526148
rect 35204 525948 35268 526012
rect 41092 525812 41156 525876
rect 514340 525812 514404 525876
rect 177620 525676 177684 525740
rect 280660 525540 280724 525604
rect 499436 525540 499500 525604
rect 44772 525404 44836 525468
rect 289124 525404 289188 525468
rect 285076 525268 285140 525332
rect 530164 525268 530228 525332
rect 46428 525132 46492 525196
rect 282868 525132 282932 525196
rect 285444 525132 285508 525196
rect 535684 525132 535748 525196
rect 41276 524996 41340 525060
rect 36492 524860 36556 524924
rect 42380 524724 42444 524788
rect 39436 524452 39500 524516
rect 512500 524452 512564 524516
rect 548380 524452 548444 524516
rect 54708 524316 54772 524380
rect 296484 524316 296548 524380
rect 480300 524316 480364 524380
rect 281028 524180 281092 524244
rect 527404 524180 527468 524244
rect 37412 524044 37476 524108
rect 288940 524044 289004 524108
rect 283604 523908 283668 523972
rect 536972 523908 537036 523972
rect 44588 523772 44652 523836
rect 46612 523500 46676 523564
rect 288388 523500 288452 523564
rect 177804 523364 177868 523428
rect 39252 523228 39316 523292
rect 57652 523152 57716 523156
rect 57652 523096 57702 523152
rect 57702 523096 57716 523152
rect 57652 523092 57716 523096
rect 503852 523092 503916 523156
rect 517836 523092 517900 523156
rect 525932 523092 525996 523156
rect 483612 522956 483676 523020
rect 519124 522956 519188 523020
rect 482140 522820 482204 522884
rect 520228 522820 520292 522884
rect 37228 522684 37292 522748
rect 478092 522684 478156 522748
rect 479380 522548 479444 522612
rect 525196 522548 525260 522612
rect 39620 522276 39684 522340
rect 292620 522276 292684 522340
rect 43484 521868 43548 521932
rect 500724 521868 500788 521932
rect 43668 521732 43732 521796
rect 499252 521732 499316 521796
rect 518204 521732 518268 521796
rect 498700 521596 498764 521660
rect 500540 521596 500604 521660
rect 530532 521596 530596 521660
rect 299796 521324 299860 521388
rect 503116 521324 503180 521388
rect 287836 521188 287900 521252
rect 505324 521188 505388 521252
rect 527220 521188 527284 521252
rect 508084 521052 508148 521116
rect 57836 520916 57900 520980
rect 254532 520916 254596 520980
rect 283420 520916 283484 520980
rect 531452 520916 531516 520980
rect 497596 520780 497660 520844
rect 508452 520780 508516 520844
rect 499436 520644 499500 520708
rect 500356 520644 500420 520708
rect 40908 520508 40972 520572
rect 499436 520508 499500 520572
rect 291884 520372 291948 520436
rect 538444 520372 538508 520436
rect 50292 520236 50356 520300
rect 51212 520236 51276 520300
rect 52132 520236 52196 520300
rect 59676 520236 59740 520300
rect 61332 520236 61396 520300
rect 61884 520296 61948 520300
rect 61884 520240 61898 520296
rect 61898 520240 61948 520296
rect 61884 520236 61948 520240
rect 497412 520236 497476 520300
rect 499988 520236 500052 520300
rect 499436 520100 499500 520164
rect 502932 520236 502996 520300
rect 515076 520236 515140 520300
rect 55444 519964 55508 520028
rect 501092 519964 501156 520028
rect 529244 519964 529308 520028
rect 500540 519692 500604 519756
rect 50660 519556 50724 519620
rect 500724 519556 500788 519620
rect 504036 519556 504100 519620
rect 507164 519692 507228 519756
rect 526300 519692 526364 519756
rect 516364 519556 516428 519620
rect 500356 519420 500420 519484
rect 522252 519420 522316 519484
rect 51580 519284 51644 519348
rect 511212 519284 511276 519348
rect 44036 518740 44100 518804
rect 31156 514932 31220 514996
rect 30420 514796 30484 514860
rect 514708 514720 514772 514724
rect 514708 514664 514722 514720
rect 514722 514664 514772 514720
rect 514708 514660 514772 514664
rect 55996 514388 56060 514452
rect 55628 513980 55692 514044
rect 510844 513436 510908 513500
rect 53788 513300 53852 513364
rect 504036 511940 504100 512004
rect 504036 511804 504100 511868
rect 50660 510580 50724 510644
rect 57652 510580 57716 510644
rect 43852 509492 43916 509556
rect 57652 508540 57716 508604
rect 41276 507316 41340 507380
rect 41276 506500 41340 506564
rect 49740 506500 49804 506564
rect 57652 505684 57716 505748
rect 57468 505276 57532 505340
rect 514708 505336 514772 505340
rect 514708 505280 514722 505336
rect 514722 505280 514772 505336
rect 514708 505276 514772 505280
rect 35572 505140 35636 505204
rect 51028 503644 51092 503708
rect 55444 503644 55508 503708
rect 54524 503508 54588 503572
rect 58572 502964 58636 503028
rect 40724 502420 40788 502484
rect 38884 502284 38948 502348
rect 36676 501876 36740 501940
rect 22692 501740 22756 501804
rect 39804 501332 39868 501396
rect 55628 500652 55692 500716
rect 52132 499836 52196 499900
rect 57468 499156 57532 499220
rect 57652 498884 57716 498948
rect 42380 498068 42444 498132
rect 36492 497524 36556 497588
rect 55996 497116 56060 497180
rect 42748 496980 42812 497044
rect 43484 496708 43548 496772
rect 57652 496436 57716 496500
rect 32444 495892 32508 495956
rect 35204 495348 35268 495412
rect 40908 494804 40972 494868
rect 39068 494668 39132 494732
rect 46428 494668 46492 494732
rect 57284 494668 57348 494732
rect 39252 494260 39316 494324
rect 44404 493988 44468 494052
rect 59676 493716 59740 493780
rect 44588 493172 44652 493236
rect 35756 492084 35820 492148
rect 46060 491812 46124 491876
rect 42564 491540 42628 491604
rect 39252 491132 39316 491196
rect 39436 490452 39500 490516
rect 35388 489364 35452 489428
rect 30972 488276 31036 488340
rect 499436 488276 499500 488340
rect 55812 487732 55876 487796
rect 27476 487188 27540 487252
rect 29684 486100 29748 486164
rect 29868 485556 29932 485620
rect 30052 485012 30116 485076
rect 522252 484740 522316 484804
rect 580580 484604 580644 484668
rect 33732 484468 33796 484532
rect 508268 484196 508332 484260
rect 36860 483924 36924 483988
rect 507164 483924 507228 483988
rect 37228 483380 37292 483444
rect 50292 482836 50356 482900
rect 500172 482896 500236 482900
rect 500172 482840 500222 482896
rect 500222 482840 500236 482896
rect 500172 482836 500236 482840
rect 500540 482156 500604 482220
rect 512500 482156 512564 482220
rect 529244 481476 529308 481540
rect 501460 481340 501524 481404
rect 503116 481340 503180 481404
rect 512132 481340 512196 481404
rect 518388 481204 518452 481268
rect 526300 480796 526364 480860
rect 502564 480388 502628 480452
rect 511212 480252 511276 480316
rect 502380 480116 502444 480180
rect 502748 479300 502812 479364
rect 502932 479028 502996 479092
rect 55996 478892 56060 478956
rect 505140 478756 505204 478820
rect 519492 478484 519556 478548
rect 516364 478212 516428 478276
rect 511028 477940 511092 478004
rect 527404 477668 527468 477732
rect 532740 477396 532804 477460
rect 534028 476852 534092 476916
rect 539732 476580 539796 476644
rect 525380 476308 525444 476372
rect 51580 476172 51644 476236
rect 505324 475764 505388 475828
rect 46060 475356 46124 475420
rect 54340 475356 54404 475420
rect 500356 475220 500420 475284
rect 508452 474948 508516 475012
rect 530164 474676 530228 474740
rect 500356 474540 500420 474604
rect 531452 474404 531516 474468
rect 536972 474132 537036 474196
rect 514156 473860 514220 473924
rect 529060 473588 529124 473652
rect 519308 473316 519372 473380
rect 538628 473180 538692 473244
rect 520412 473044 520476 473108
rect 512316 472772 512380 472836
rect 539548 472500 539612 472564
rect 538444 471956 538508 472020
rect 535684 471684 535748 471748
rect 547092 471412 547156 471476
rect 514524 470868 514588 470932
rect 515260 470596 515324 470660
rect 526116 470324 526180 470388
rect 523172 470052 523236 470116
rect 516180 469780 516244 469844
rect 523540 467876 523604 467940
rect 3372 462572 3436 462636
rect 46796 458356 46860 458420
rect 48636 457812 48700 457876
rect 54892 456180 54956 456244
rect 47900 455636 47964 455700
rect 47716 455092 47780 455156
rect 48452 454548 48516 454612
rect 501276 454548 501340 454612
rect 33916 454004 33980 454068
rect 58756 453460 58820 453524
rect 536788 453460 536852 453524
rect 54340 452916 54404 452980
rect 26004 452372 26068 452436
rect 28764 451828 28828 451892
rect 48084 451284 48148 451348
rect 31524 450740 31588 450804
rect 34284 450196 34348 450260
rect 54708 449652 54772 449716
rect 3740 449516 3804 449580
rect 32996 449108 33060 449172
rect 57284 448564 57348 448628
rect 31340 448020 31404 448084
rect 53604 447476 53668 447540
rect 59124 446932 59188 446996
rect 58388 446388 58452 446452
rect 59860 445844 59924 445908
rect 52316 445300 52380 445364
rect 41092 444756 41156 444820
rect 57836 444212 57900 444276
rect 39620 443668 39684 443732
rect 44772 443124 44836 443188
rect 37412 442580 37476 442644
rect 37044 442036 37108 442100
rect 32812 441492 32876 441556
rect 34100 440948 34164 441012
rect 32628 440404 32692 440468
rect 47532 439860 47596 439924
rect 46612 439316 46676 439380
rect 44956 438772 45020 438836
rect 525196 436052 525260 436116
rect 519124 435236 519188 435300
rect 520228 434964 520292 435028
rect 544332 418236 544396 418300
rect 41276 417012 41340 417076
rect 39252 416468 39316 416532
rect 39068 415924 39132 415988
rect 42380 415380 42444 415444
rect 30236 414836 30300 414900
rect 38884 414292 38948 414356
rect 44404 413748 44468 413812
rect 3924 410484 3988 410548
rect 2820 398108 2884 398172
rect 3556 397428 3620 397492
rect 357940 390220 358004 390284
rect 543228 390220 543292 390284
rect 501092 389948 501156 390012
rect 543228 389132 543292 389196
rect 345612 388588 345676 388652
rect 538812 388588 538876 388652
rect 500356 388044 500420 388108
rect 349660 387908 349724 387972
rect 361620 386820 361684 386884
rect 362908 386820 362972 386884
rect 360148 386684 360212 386748
rect 360332 386412 360396 386476
rect 349844 385732 349908 385796
rect 356652 384780 356716 384844
rect 543780 384780 543844 384844
rect 351132 384644 351196 384708
rect 546540 384644 546604 384708
rect 346900 384508 346964 384572
rect 550956 384508 551020 384572
rect 354628 383964 354692 384028
rect 353892 383828 353956 383892
rect 358124 383012 358188 383076
rect 3740 382876 3804 382940
rect 137140 382876 137204 382940
rect 356836 382196 356900 382260
rect 355180 381924 355244 381988
rect 550036 381924 550100 381988
rect 338620 381788 338684 381852
rect 550772 381788 550836 381852
rect 239812 380156 239876 380220
rect 580212 380156 580276 380220
rect 355548 379340 355612 379404
rect 538628 379340 538692 379404
rect 547644 379340 547708 379404
rect 352972 379204 353036 379268
rect 234476 377436 234540 377500
rect 354076 376484 354140 376548
rect 550588 376484 550652 376548
rect 357204 375396 357268 375460
rect 284892 375124 284956 375188
rect 282132 374716 282196 374780
rect 538260 374716 538324 374780
rect 282316 373356 282380 373420
rect 541020 373356 541084 373420
rect 351316 371996 351380 372060
rect 543228 371996 543292 372060
rect 542676 371316 542740 371380
rect 287836 371180 287900 371244
rect 282684 370500 282748 370564
rect 541204 370500 541268 370564
rect 282500 369004 282564 369068
rect 539364 369004 539428 369068
rect 352788 367644 352852 367708
rect 542860 367644 542924 367708
rect 234292 366420 234356 366484
rect 357020 365332 357084 365396
rect 543412 365332 543476 365396
rect 354260 365196 354324 365260
rect 542676 365196 542740 365260
rect 580212 365060 580276 365124
rect 234108 364924 234172 364988
rect 355364 363564 355428 363628
rect 543044 363564 543108 363628
rect 239628 362204 239692 362268
rect 580396 362204 580460 362268
rect 239444 360980 239508 361044
rect 580580 360980 580644 361044
rect 43668 360844 43732 360908
rect 282868 357504 282932 357508
rect 282868 357448 282918 357504
rect 282918 357448 282932 357504
rect 282868 357444 282932 357448
rect 3372 355948 3436 356012
rect 530532 355948 530596 356012
rect 533292 355948 533356 356012
rect 534580 355948 534644 356012
rect 284340 355056 284404 355060
rect 284340 355000 284354 355056
rect 284354 355000 284404 355056
rect 284340 354996 284404 355000
rect 31156 354588 31220 354652
rect 504220 354316 504284 354380
rect 506980 354180 507044 354244
rect 3924 353908 3988 353972
rect 283052 353908 283116 353972
rect 235764 353772 235828 353836
rect 231164 353500 231228 353564
rect 285812 353500 285876 353564
rect 239260 353364 239324 353428
rect 50844 352548 50908 352612
rect 229876 351112 229940 351116
rect 229876 351056 229926 351112
rect 229926 351056 229940 351112
rect 229876 351052 229940 351056
rect 235212 349148 235276 349212
rect 298140 349208 298204 349212
rect 298140 349152 298154 349208
rect 298154 349152 298204 349208
rect 298140 349148 298204 349152
rect 361620 349012 361684 349076
rect 362908 348876 362972 348940
rect 227484 347924 227548 347988
rect 299428 347924 299492 347988
rect 226932 347788 226996 347852
rect 299612 347788 299676 347852
rect 223436 347516 223500 347580
rect 288572 347516 288636 347580
rect 224356 346836 224420 346900
rect 279004 346836 279068 346900
rect 227116 346700 227180 346764
rect 291332 346700 291396 346764
rect 214788 346564 214852 346628
rect 48084 346428 48148 346492
rect 226196 346156 226260 346220
rect 290780 346156 290844 346220
rect 360148 345748 360212 345812
rect 217548 345612 217612 345676
rect 280660 345612 280724 345676
rect 284524 345612 284588 345676
rect 228220 345476 228284 345540
rect 287652 345476 287716 345540
rect 4108 345340 4172 345404
rect 222700 345340 222764 345404
rect 227300 345340 227364 345404
rect 288388 345340 288452 345404
rect 217364 344932 217428 344996
rect 218652 344796 218716 344860
rect 306420 344796 306484 344860
rect 224540 343844 224604 343908
rect 303660 343844 303724 343908
rect 214604 342756 214668 342820
rect 231348 342756 231412 342820
rect 295564 342756 295628 342820
rect 214420 342484 214484 342548
rect 224724 342484 224788 342548
rect 295380 342484 295444 342548
rect 220308 341940 220372 342004
rect 224908 341532 224972 341596
rect 279556 341532 279620 341596
rect 222884 341124 222948 341188
rect 280292 341124 280356 341188
rect 286916 341124 286980 341188
rect 231532 340988 231596 341052
rect 290596 340988 290660 341052
rect 211660 340852 211724 340916
rect 296484 340852 296548 340916
rect 221228 340580 221292 340644
rect 279924 340580 279988 340644
rect 221044 340308 221108 340372
rect 267596 340308 267660 340372
rect 279740 340308 279804 340372
rect 215892 340172 215956 340236
rect 237972 340172 238036 340236
rect 238156 340172 238220 340236
rect 280108 340172 280172 340236
rect 217180 339628 217244 339692
rect 296852 339628 296916 339692
rect 219940 339492 220004 339556
rect 230244 339492 230308 339556
rect 238156 339492 238220 339556
rect 256004 339492 256068 339556
rect 274588 339492 274652 339556
rect 218836 338948 218900 339012
rect 279004 339356 279068 339420
rect 256004 338948 256068 339012
rect 274588 338948 274652 339012
rect 303844 338948 303908 339012
rect 4108 338676 4172 338740
rect 230980 338676 231044 338740
rect 279924 338812 279988 338876
rect 267596 338540 267660 338604
rect 291516 338540 291580 338604
rect 220492 338404 220556 338468
rect 294644 338404 294708 338468
rect 216076 338268 216140 338332
rect 224172 338132 224236 338196
rect 301820 338132 301884 338196
rect 279556 337996 279620 338060
rect 290780 337996 290844 338060
rect 279740 337860 279804 337924
rect 220124 337724 220188 337788
rect 290964 337724 291028 337788
rect 285996 336636 286060 336700
rect 3556 326300 3620 326364
rect 522068 315828 522132 315892
rect 580396 312020 580460 312084
rect 234108 309844 234172 309908
rect 521884 309844 521948 309908
rect 280476 309300 280540 309364
rect 214788 306172 214852 306236
rect 284524 303316 284588 303380
rect 294460 301684 294524 301748
rect 55076 301412 55140 301476
rect 291148 300596 291212 300660
rect 292620 300052 292684 300116
rect 287836 299372 287900 299436
rect 223068 298556 223132 298620
rect 216628 298012 216692 298076
rect 287284 297876 287348 297940
rect 287100 297332 287164 297396
rect 217548 296924 217612 296988
rect 285628 296788 285692 296852
rect 287468 296244 287532 296308
rect 217364 295292 217428 295356
rect 220308 293660 220372 293724
rect 3372 293116 3436 293180
rect 284524 291348 284588 291412
rect 220492 290396 220556 290460
rect 226196 289716 226260 289780
rect 357204 289172 357268 289236
rect 226012 288764 226076 288828
rect 354076 288628 354140 288692
rect 352972 288084 353036 288148
rect 355548 287540 355612 287604
rect 228220 287132 228284 287196
rect 234476 286996 234540 287060
rect 355180 285908 355244 285972
rect 231532 285500 231596 285564
rect 48084 284956 48148 285020
rect 234292 284820 234356 284884
rect 354260 284276 354324 284340
rect 235764 283732 235828 283796
rect 356836 283188 356900 283252
rect 224908 282372 224972 282436
rect 224908 282236 224972 282300
rect 358124 282100 358188 282164
rect 349844 281012 349908 281076
rect 222884 280604 222948 280668
rect 354444 280604 354508 280668
rect 518940 279924 519004 279988
rect 353892 279380 353956 279444
rect 338620 278292 338684 278356
rect 356652 277204 356716 277268
rect 351132 276660 351196 276724
rect 542860 276660 542924 276724
rect 580396 276660 580460 276724
rect 346900 276116 346964 276180
rect 220124 275708 220188 275772
rect 349660 275572 349724 275636
rect 351316 275028 351380 275092
rect 282316 274484 282380 274548
rect 227484 274076 227548 274140
rect 352788 273940 352852 274004
rect 282684 273396 282748 273460
rect 357020 272852 357084 272916
rect 226932 272444 226996 272508
rect 282132 272308 282196 272372
rect 355364 271764 355428 271828
rect 357940 271220 358004 271284
rect 227116 270812 227180 270876
rect 282500 270676 282564 270740
rect 345612 270132 345676 270196
rect 227300 269180 227364 269244
rect 518204 267956 518268 268020
rect 231348 267548 231412 267612
rect 211660 265916 211724 265980
rect 215892 264284 215956 264348
rect 216076 262652 216140 262716
rect 518020 261972 518084 262036
rect 284892 260068 284956 260132
rect 508452 258844 508516 258908
rect 224356 257756 224420 257820
rect 223620 256668 223684 256732
rect 221044 256124 221108 256188
rect 220860 255308 220924 255372
rect 224540 254492 224604 254556
rect 48636 254084 48700 254148
rect 223804 253948 223868 254012
rect 224724 252860 224788 252924
rect 230060 252452 230124 252516
rect 230244 251228 230308 251292
rect 224172 249596 224236 249660
rect 288572 249460 288636 249524
rect 238340 246740 238404 246804
rect 218836 246332 218900 246396
rect 197860 245652 197924 245716
rect 287652 245652 287716 245716
rect 290596 245108 290660 245172
rect 231164 244700 231228 244764
rect 285996 244020 286060 244084
rect 280292 243476 280356 243540
rect 221228 243068 221292 243132
rect 210556 242388 210620 242452
rect 290780 241844 290844 241908
rect 218652 241436 218716 241500
rect 299428 241300 299492 241364
rect 3556 241028 3620 241092
rect 299612 240756 299676 240820
rect 291332 240212 291396 240276
rect 288388 239668 288452 239732
rect 237788 239124 237852 239188
rect 295564 239124 295628 239188
rect 296668 238580 296732 238644
rect 237604 238036 237668 238100
rect 296852 238036 296916 238100
rect 238156 236948 238220 237012
rect 237972 235996 238036 236060
rect 59124 235860 59188 235924
rect 291516 235316 291580 235380
rect 60412 235180 60476 235244
rect 238340 235180 238404 235244
rect 237972 234772 238036 234836
rect 303660 234772 303724 234836
rect 295380 234228 295444 234292
rect 58572 233684 58636 233748
rect 280292 233684 280356 233748
rect 301820 233140 301884 233204
rect 303844 232052 303908 232116
rect 237420 231508 237484 231572
rect 285812 231508 285876 231572
rect 60044 231100 60108 231164
rect 237604 231100 237668 231164
rect 294644 230964 294708 231028
rect 306420 230420 306484 230484
rect 3372 228244 3436 228308
rect 214788 228244 214852 228308
rect 58940 226884 59004 226948
rect 237420 226884 237484 226948
rect 238524 226400 238588 226404
rect 238524 226344 238574 226400
rect 238574 226344 238588 226400
rect 238524 226340 238588 226344
rect 60228 225524 60292 225588
rect 237788 225524 237852 225588
rect 3556 218588 3620 218652
rect 213132 218588 213196 218652
rect 281764 214644 281828 214708
rect 286916 210020 286980 210084
rect 280844 208660 280908 208724
rect 58756 207572 58820 207636
rect 237972 207572 238036 207636
rect 282132 204852 282196 204916
rect 234660 201860 234724 201924
rect 285812 199956 285876 200020
rect 281580 198868 281644 198932
rect 281948 197780 282012 197844
rect 280660 197236 280724 197300
rect 284708 196692 284772 196756
rect 60596 195196 60660 195260
rect 238156 195196 238220 195260
rect 284892 193972 284956 194036
rect 18460 193836 18524 193900
rect 237972 193836 238036 193900
rect 15700 192476 15764 192540
rect 237420 192476 237484 192540
rect 283236 191796 283300 191860
rect 281028 191252 281092 191316
rect 26740 190980 26804 191044
rect 238156 190980 238220 191044
rect 302924 190164 302988 190228
rect 57468 189620 57532 189684
rect 210556 189620 210620 189684
rect 346900 189620 346964 189684
rect 345612 189076 345676 189140
rect 3372 188804 3436 188868
rect 327764 188532 327828 188596
rect 22692 188260 22756 188324
rect 238340 188260 238404 188324
rect 290780 187988 290844 188052
rect 237420 187716 237484 187780
rect 313964 187444 314028 187508
rect 57652 186900 57716 186964
rect 197860 186900 197924 186964
rect 338620 186900 338684 186964
rect 300164 186356 300228 186420
rect 334572 185812 334636 185876
rect 3372 185540 3436 185604
rect 235396 185540 235460 185604
rect 291884 185268 291948 185332
rect 319300 184724 319364 184788
rect 3372 184452 3436 184516
rect 134380 184452 134444 184516
rect 298876 184180 298940 184244
rect 342852 183636 342916 183700
rect 349660 183092 349724 183156
rect 335860 182548 335924 182612
rect 59676 182004 59740 182068
rect 294828 182004 294892 182068
rect 60412 181732 60476 181796
rect 307156 181460 307220 181524
rect 407620 181324 407684 181388
rect 214604 180916 214668 180980
rect 353892 180916 353956 180980
rect 525748 180508 525812 180572
rect 309732 180372 309796 180436
rect 535500 180372 535564 180436
rect 529980 180236 530044 180300
rect 517836 180100 517900 180164
rect 57652 179828 57716 179892
rect 351132 179828 351196 179892
rect 514892 179964 514956 180028
rect 57836 179480 57900 179484
rect 57836 179424 57886 179480
rect 57886 179424 57900 179480
rect 57836 179420 57900 179424
rect 214420 179148 214484 179212
rect 504036 179284 504100 179348
rect 334756 179148 334820 179212
rect 510660 179012 510724 179076
rect 503668 178876 503732 178940
rect 296116 178740 296180 178804
rect 503116 178740 503180 178804
rect 355180 178604 355244 178668
rect 327580 178196 327644 178260
rect 522988 177924 523052 177988
rect 512132 177788 512196 177852
rect 217180 177652 217244 177716
rect 302740 177652 302804 177716
rect 521700 177652 521764 177716
rect 515076 177516 515140 177580
rect 525932 177380 525996 177444
rect 499804 177244 499868 177308
rect 294644 177108 294708 177172
rect 299980 176564 300044 176628
rect 510476 176564 510540 176628
rect 57652 176428 57716 176492
rect 527220 176428 527284 176492
rect 509004 176292 509068 176356
rect 57836 176020 57900 176084
rect 216628 176156 216692 176220
rect 510844 176156 510908 176220
rect 289492 176020 289556 176084
rect 499620 176020 499684 176084
rect 356652 175476 356716 175540
rect 57836 175204 57900 175268
rect 506796 175204 506860 175268
rect 500172 175068 500236 175132
rect 288940 174932 289004 174996
rect 501644 174932 501708 174996
rect 503852 174796 503916 174860
rect 507900 174660 507964 174724
rect 289492 174524 289556 174588
rect 357940 174524 358004 174588
rect 506612 174524 506676 174588
rect 226196 174388 226260 174452
rect 305500 174388 305564 174452
rect 514708 174388 514772 174452
rect 57468 174116 57532 174180
rect 295932 173844 295996 173908
rect 304212 173300 304276 173364
rect 219940 172756 220004 172820
rect 322060 172756 322124 172820
rect 57284 172348 57348 172412
rect 57652 172212 57716 172276
rect 323532 172212 323596 172276
rect 231164 171668 231228 171732
rect 311020 171668 311084 171732
rect 220860 171124 220924 171188
rect 291700 171124 291764 171188
rect 228220 170580 228284 170644
rect 57836 170308 57900 170372
rect 282132 169764 282196 169828
rect 223804 169628 223868 169692
rect 134380 169492 134444 169556
rect 290596 169492 290660 169556
rect 360332 169084 360396 169148
rect 291332 168948 291396 169012
rect 59860 168676 59924 168740
rect 60228 168404 60292 168468
rect 235396 168404 235460 168468
rect 223620 167860 223684 167924
rect 213132 167316 213196 167380
rect 58572 167044 58636 167108
rect 60044 166500 60108 166564
rect 214788 166364 214852 166428
rect 229876 166228 229940 166292
rect 283052 166228 283116 166292
rect 284340 165684 284404 165748
rect 230980 165140 231044 165204
rect 60596 164596 60660 164660
rect 222700 164596 222764 164660
rect 282868 164596 282932 164660
rect 298140 164052 298204 164116
rect 224908 163100 224972 163164
rect 137140 162964 137204 163028
rect 59124 162692 59188 162756
rect 59308 162692 59372 162756
rect 293356 162012 293420 162076
rect 580212 162012 580276 162076
rect 238340 161876 238404 161940
rect 230060 161332 230124 161396
rect 58756 160788 58820 160852
rect 237972 160788 238036 160852
rect 58756 160108 58820 160172
rect 235580 159700 235644 159764
rect 238156 159700 238220 159764
rect 508084 159156 508148 159220
rect 57652 158884 57716 158948
rect 57836 158748 57900 158812
rect 235764 158068 235828 158132
rect 558132 158068 558196 158132
rect 555372 157524 555436 157588
rect 58572 156980 58636 157044
rect 551140 156980 551204 157044
rect 58388 156572 58452 156636
rect 235212 156572 235276 156636
rect 235396 156436 235460 156500
rect 548380 156436 548444 156500
rect 58572 155892 58636 155956
rect 234660 155892 234724 155956
rect 547092 155892 547156 155956
rect 544332 155348 544396 155412
rect 58940 155076 59004 155140
rect 235212 154804 235276 154868
rect 293356 154804 293420 154868
rect 57468 154396 57532 154460
rect 542860 154260 542924 154324
rect 508452 153716 508516 153780
rect 57284 153172 57348 153236
rect 334756 152628 334820 152692
rect 306420 152084 306484 152148
rect 238156 151540 238220 151604
rect 313780 151540 313844 151604
rect 58756 151268 58820 151332
rect 306420 150996 306484 151060
rect 580212 150996 580276 151060
rect 306972 150860 307036 150924
rect 298692 150452 298756 150516
rect 237972 149908 238036 149972
rect 54340 149772 54404 149836
rect 59124 149364 59188 149428
rect 127572 148276 127636 148340
rect 58572 147460 58636 147524
rect 127756 146644 127820 146708
rect 239812 145624 239876 145688
rect 58388 145556 58452 145620
rect 127940 145012 128004 145076
rect 57652 144740 57716 144804
rect 239628 144536 239692 144600
rect 407620 144740 407684 144804
rect 57836 143652 57900 143716
rect 239812 143448 239876 143512
rect 128124 143380 128188 143444
rect 302924 142700 302988 142764
rect 239628 142360 239692 142424
rect 57652 141748 57716 141812
rect 238524 141340 238588 141404
rect 327764 141340 327828 141404
rect 357388 141340 357452 141404
rect 346900 140252 346964 140316
rect 290780 139980 290844 140044
rect 357572 139980 357636 140044
rect 57468 139844 57532 139908
rect 580212 139300 580276 139364
rect 345612 139164 345676 139228
rect 59860 138484 59924 138548
rect 357388 138076 357452 138140
rect 338620 137260 338684 137324
rect 357388 137260 357452 137324
rect 357572 136988 357636 137052
rect 238340 136852 238404 136916
rect 3372 136716 3436 136780
rect 59676 136036 59740 136100
rect 313964 135900 314028 135964
rect 238524 135764 238588 135828
rect 280108 135144 280172 135148
rect 280108 135088 280122 135144
rect 280122 135088 280172 135144
rect 280108 135084 280172 135088
rect 357388 134812 357452 134876
rect 239628 134744 239692 134808
rect 281948 134676 282012 134740
rect 334572 134404 334636 134468
rect 357388 134404 357452 134468
rect 300164 133724 300228 133788
rect 239444 133588 239508 133652
rect 357388 132636 357452 132700
rect 239812 132568 239876 132632
rect 291884 131548 291948 131612
rect 291516 131140 291580 131204
rect 319300 130460 319364 130524
rect 298876 129372 298940 129436
rect 342852 128284 342916 128348
rect 349660 127196 349724 127260
rect 335860 126108 335924 126172
rect 294276 125428 294340 125492
rect 294828 125020 294892 125084
rect 307156 123932 307220 123996
rect 237788 123796 237852 123860
rect 238340 123524 238404 123588
rect 353892 122844 353956 122908
rect 309732 121756 309796 121820
rect 57836 121484 57900 121548
rect 127572 121348 127636 121412
rect 287284 121348 287348 121412
rect 128124 121212 128188 121276
rect 287468 121212 287532 121276
rect 296116 120804 296180 120868
rect 357572 120804 357636 120868
rect 351132 120668 351196 120732
rect 234660 120532 234724 120596
rect 235212 120124 235276 120188
rect 292620 120396 292684 120460
rect 238524 119988 238588 120052
rect 284524 119988 284588 120052
rect 127756 119852 127820 119916
rect 287100 119852 287164 119916
rect 127940 119716 128004 119780
rect 285628 119716 285692 119780
rect 355180 119580 355244 119644
rect 48636 119308 48700 119372
rect 235764 119308 235828 119372
rect 238156 119308 238220 119372
rect 294276 119444 294340 119508
rect 327580 119308 327644 119372
rect 357388 119308 357452 119372
rect 291516 119172 291580 119236
rect 291884 118764 291948 118828
rect 235580 118492 235644 118556
rect 294460 118492 294524 118556
rect 357572 118492 357636 118556
rect 237972 118356 238036 118420
rect 237788 117404 237852 117468
rect 357388 117404 357452 117468
rect 280844 116588 280908 116652
rect 302740 116316 302804 116380
rect 54340 116044 54404 116108
rect 291332 116044 291396 116108
rect 235396 115228 235460 115292
rect 291148 115228 291212 115292
rect 294644 115228 294708 115292
rect 281764 114276 281828 114340
rect 299980 114140 300044 114204
rect 3372 113188 3436 113252
rect 357940 113052 358004 113116
rect 580212 112780 580276 112844
rect 356652 112644 356716 112708
rect 288940 112508 289004 112572
rect 46060 112372 46124 112436
rect 291884 112372 291948 112436
rect 305500 111012 305564 111076
rect 284892 109652 284956 109716
rect 295932 109652 295996 109716
rect 304212 107612 304276 107676
rect 322060 106524 322124 106588
rect 323532 105436 323596 105500
rect 311020 104348 311084 104412
rect 281028 104076 281092 104140
rect 291700 103260 291764 103324
rect 239628 100676 239692 100740
rect 580212 100676 580276 100740
rect 313780 99452 313844 99516
rect 283236 98772 283300 98836
rect 239444 98636 239508 98700
rect 580212 98636 580276 98700
rect 290596 97548 290660 97612
rect 278820 94420 278884 94484
rect 3556 86260 3620 86324
rect 228220 86260 228284 86324
rect 3556 84628 3620 84692
rect 580212 72932 580276 72996
rect 281580 62732 281644 62796
rect 306972 59604 307036 59668
rect 46060 58516 46124 58580
rect 57836 51444 57900 51508
rect 57836 46140 57900 46204
rect 231164 45460 231228 45524
rect 280660 44916 280724 44980
rect 239812 33084 239876 33148
rect 284708 29684 284772 29748
rect 285812 22748 285876 22812
rect 298692 19756 298756 19820
rect 3372 19348 3436 19412
rect 4108 7652 4172 7716
rect 234660 7652 234724 7716
rect 4108 6428 4172 6492
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 677494 -8106 711002
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 -8106 677494
rect -8726 677174 -8106 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 -8106 677174
rect -8726 641494 -8106 676938
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 -8106 641494
rect -8726 641174 -8106 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 -8106 641174
rect -8726 605494 -8106 640938
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 -8106 605494
rect -8726 605174 -8106 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 -8106 605174
rect -8726 569494 -8106 604938
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 -8106 569494
rect -8726 569174 -8106 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 -8106 569174
rect -8726 533494 -8106 568938
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 -8106 533494
rect -8726 533174 -8106 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 -8106 533174
rect -8726 497494 -8106 532938
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 -8106 497494
rect -8726 497174 -8106 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 -8106 497174
rect -8726 461494 -8106 496938
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 -8106 461494
rect -8726 461174 -8106 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 -8106 461174
rect -8726 425494 -8106 460938
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 -8106 425494
rect -8726 425174 -8106 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 -8106 425174
rect -8726 389494 -8106 424938
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 -8106 389494
rect -8726 389174 -8106 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 -8106 389174
rect -8726 353494 -8106 388938
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 -8106 353494
rect -8726 353174 -8106 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 -8106 353174
rect -8726 317494 -8106 352938
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 -8106 317494
rect -8726 317174 -8106 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 -8106 317174
rect -8726 281494 -8106 316938
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 -8106 281494
rect -8726 281174 -8106 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 -8106 281174
rect -8726 245494 -8106 280938
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 -8106 245494
rect -8726 245174 -8106 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 -8106 245174
rect -8726 209494 -8106 244938
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 -8106 209494
rect -8726 209174 -8106 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 -8106 209174
rect -8726 173494 -8106 208938
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 -8106 173494
rect -8726 173174 -8106 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 -8106 173174
rect -8726 137494 -8106 172938
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 -8106 137494
rect -8726 137174 -8106 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 -8106 137174
rect -8726 101494 -8106 136938
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 -8106 101494
rect -8726 101174 -8106 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 -8106 101174
rect -8726 65494 -8106 100938
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 -8106 65494
rect -8726 65174 -8106 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 -8106 65174
rect -8726 29494 -8106 64938
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 -8106 29494
rect -8726 29174 -8106 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 -8106 29174
rect -8726 -7066 -8106 28938
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 673774 -7146 710042
rect -7766 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 -7146 673774
rect -7766 673454 -7146 673538
rect -7766 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 -7146 673454
rect -7766 637774 -7146 673218
rect -7766 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 -7146 637774
rect -7766 637454 -7146 637538
rect -7766 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 -7146 637454
rect -7766 601774 -7146 637218
rect -7766 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 -7146 601774
rect -7766 601454 -7146 601538
rect -7766 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 -7146 601454
rect -7766 565774 -7146 601218
rect -7766 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 -7146 565774
rect -7766 565454 -7146 565538
rect -7766 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 -7146 565454
rect -7766 529774 -7146 565218
rect -7766 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 -7146 529774
rect -7766 529454 -7146 529538
rect -7766 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 -7146 529454
rect -7766 493774 -7146 529218
rect -7766 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 -7146 493774
rect -7766 493454 -7146 493538
rect -7766 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 -7146 493454
rect -7766 457774 -7146 493218
rect -7766 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 -7146 457774
rect -7766 457454 -7146 457538
rect -7766 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 -7146 457454
rect -7766 421774 -7146 457218
rect -7766 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 -7146 421774
rect -7766 421454 -7146 421538
rect -7766 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 -7146 421454
rect -7766 385774 -7146 421218
rect -7766 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 -7146 385774
rect -7766 385454 -7146 385538
rect -7766 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 -7146 385454
rect -7766 349774 -7146 385218
rect -7766 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 -7146 349774
rect -7766 349454 -7146 349538
rect -7766 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 -7146 349454
rect -7766 313774 -7146 349218
rect -7766 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 -7146 313774
rect -7766 313454 -7146 313538
rect -7766 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 -7146 313454
rect -7766 277774 -7146 313218
rect -7766 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 -7146 277774
rect -7766 277454 -7146 277538
rect -7766 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 -7146 277454
rect -7766 241774 -7146 277218
rect -7766 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 -7146 241774
rect -7766 241454 -7146 241538
rect -7766 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 -7146 241454
rect -7766 205774 -7146 241218
rect -7766 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 -7146 205774
rect -7766 205454 -7146 205538
rect -7766 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 -7146 205454
rect -7766 169774 -7146 205218
rect -7766 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 -7146 169774
rect -7766 169454 -7146 169538
rect -7766 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 -7146 169454
rect -7766 133774 -7146 169218
rect -7766 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 -7146 133774
rect -7766 133454 -7146 133538
rect -7766 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 -7146 133454
rect -7766 97774 -7146 133218
rect -7766 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 -7146 97774
rect -7766 97454 -7146 97538
rect -7766 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 -7146 97454
rect -7766 61774 -7146 97218
rect -7766 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 -7146 61774
rect -7766 61454 -7146 61538
rect -7766 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 -7146 61454
rect -7766 25774 -7146 61218
rect -7766 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 -7146 25774
rect -7766 25454 -7146 25538
rect -7766 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 -7146 25454
rect -7766 -6106 -7146 25218
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 670054 -6186 709082
rect -6806 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 -6186 670054
rect -6806 669734 -6186 669818
rect -6806 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 -6186 669734
rect -6806 634054 -6186 669498
rect -6806 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 -6186 634054
rect -6806 633734 -6186 633818
rect -6806 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 -6186 633734
rect -6806 598054 -6186 633498
rect -6806 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 -6186 598054
rect -6806 597734 -6186 597818
rect -6806 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 -6186 597734
rect -6806 562054 -6186 597498
rect -6806 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 -6186 562054
rect -6806 561734 -6186 561818
rect -6806 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 -6186 561734
rect -6806 526054 -6186 561498
rect -6806 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 -6186 526054
rect -6806 525734 -6186 525818
rect -6806 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 -6186 525734
rect -6806 490054 -6186 525498
rect -6806 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 -6186 490054
rect -6806 489734 -6186 489818
rect -6806 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 -6186 489734
rect -6806 454054 -6186 489498
rect -6806 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 -6186 454054
rect -6806 453734 -6186 453818
rect -6806 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 -6186 453734
rect -6806 418054 -6186 453498
rect -6806 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 -6186 418054
rect -6806 417734 -6186 417818
rect -6806 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 -6186 417734
rect -6806 382054 -6186 417498
rect -6806 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 -6186 382054
rect -6806 381734 -6186 381818
rect -6806 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 -6186 381734
rect -6806 346054 -6186 381498
rect -6806 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 -6186 346054
rect -6806 345734 -6186 345818
rect -6806 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 -6186 345734
rect -6806 310054 -6186 345498
rect -6806 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 -6186 310054
rect -6806 309734 -6186 309818
rect -6806 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 -6186 309734
rect -6806 274054 -6186 309498
rect -6806 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 -6186 274054
rect -6806 273734 -6186 273818
rect -6806 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 -6186 273734
rect -6806 238054 -6186 273498
rect -6806 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 -6186 238054
rect -6806 237734 -6186 237818
rect -6806 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 -6186 237734
rect -6806 202054 -6186 237498
rect -6806 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 -6186 202054
rect -6806 201734 -6186 201818
rect -6806 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 -6186 201734
rect -6806 166054 -6186 201498
rect -6806 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 -6186 166054
rect -6806 165734 -6186 165818
rect -6806 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 -6186 165734
rect -6806 130054 -6186 165498
rect -6806 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 -6186 130054
rect -6806 129734 -6186 129818
rect -6806 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 -6186 129734
rect -6806 94054 -6186 129498
rect -6806 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 -6186 94054
rect -6806 93734 -6186 93818
rect -6806 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 -6186 93734
rect -6806 58054 -6186 93498
rect -6806 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 -6186 58054
rect -6806 57734 -6186 57818
rect -6806 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 -6186 57734
rect -6806 22054 -6186 57498
rect -6806 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 -6186 22054
rect -6806 21734 -6186 21818
rect -6806 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 -6186 21734
rect -6806 -5146 -6186 21498
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 666334 -5226 708122
rect -5846 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 -5226 666334
rect -5846 666014 -5226 666098
rect -5846 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 -5226 666014
rect -5846 630334 -5226 665778
rect -5846 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 -5226 630334
rect -5846 630014 -5226 630098
rect -5846 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 -5226 630014
rect -5846 594334 -5226 629778
rect -5846 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 -5226 594334
rect -5846 594014 -5226 594098
rect -5846 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 -5226 594014
rect -5846 558334 -5226 593778
rect -5846 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 -5226 558334
rect -5846 558014 -5226 558098
rect -5846 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 -5226 558014
rect -5846 522334 -5226 557778
rect -5846 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 -5226 522334
rect -5846 522014 -5226 522098
rect -5846 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 -5226 522014
rect -5846 486334 -5226 521778
rect -5846 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 -5226 486334
rect -5846 486014 -5226 486098
rect -5846 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 -5226 486014
rect -5846 450334 -5226 485778
rect -5846 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 -5226 450334
rect -5846 450014 -5226 450098
rect -5846 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 -5226 450014
rect -5846 414334 -5226 449778
rect -5846 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 -5226 414334
rect -5846 414014 -5226 414098
rect -5846 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 -5226 414014
rect -5846 378334 -5226 413778
rect -5846 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 -5226 378334
rect -5846 378014 -5226 378098
rect -5846 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 -5226 378014
rect -5846 342334 -5226 377778
rect -5846 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 -5226 342334
rect -5846 342014 -5226 342098
rect -5846 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 -5226 342014
rect -5846 306334 -5226 341778
rect -5846 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 -5226 306334
rect -5846 306014 -5226 306098
rect -5846 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 -5226 306014
rect -5846 270334 -5226 305778
rect -5846 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 -5226 270334
rect -5846 270014 -5226 270098
rect -5846 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 -5226 270014
rect -5846 234334 -5226 269778
rect -5846 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 -5226 234334
rect -5846 234014 -5226 234098
rect -5846 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 -5226 234014
rect -5846 198334 -5226 233778
rect -5846 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 -5226 198334
rect -5846 198014 -5226 198098
rect -5846 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 -5226 198014
rect -5846 162334 -5226 197778
rect -5846 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 -5226 162334
rect -5846 162014 -5226 162098
rect -5846 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 -5226 162014
rect -5846 126334 -5226 161778
rect -5846 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 -5226 126334
rect -5846 126014 -5226 126098
rect -5846 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 -5226 126014
rect -5846 90334 -5226 125778
rect -5846 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 -5226 90334
rect -5846 90014 -5226 90098
rect -5846 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 -5226 90014
rect -5846 54334 -5226 89778
rect -5846 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 -5226 54334
rect -5846 54014 -5226 54098
rect -5846 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 -5226 54014
rect -5846 18334 -5226 53778
rect -5846 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 -5226 18334
rect -5846 18014 -5226 18098
rect -5846 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 -5226 18014
rect -5846 -4186 -5226 17778
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 698614 -4266 707162
rect -4886 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 -4266 698614
rect -4886 698294 -4266 698378
rect -4886 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 -4266 698294
rect -4886 662614 -4266 698058
rect -4886 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 -4266 662614
rect -4886 662294 -4266 662378
rect -4886 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 -4266 662294
rect -4886 626614 -4266 662058
rect -4886 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 -4266 626614
rect -4886 626294 -4266 626378
rect -4886 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 -4266 626294
rect -4886 590614 -4266 626058
rect -4886 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 -4266 590614
rect -4886 590294 -4266 590378
rect -4886 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 -4266 590294
rect -4886 554614 -4266 590058
rect -4886 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 -4266 554614
rect -4886 554294 -4266 554378
rect -4886 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 -4266 554294
rect -4886 518614 -4266 554058
rect -4886 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 -4266 518614
rect -4886 518294 -4266 518378
rect -4886 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 -4266 518294
rect -4886 482614 -4266 518058
rect -4886 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 -4266 482614
rect -4886 482294 -4266 482378
rect -4886 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 -4266 482294
rect -4886 446614 -4266 482058
rect -4886 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 -4266 446614
rect -4886 446294 -4266 446378
rect -4886 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 -4266 446294
rect -4886 410614 -4266 446058
rect -4886 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 -4266 410614
rect -4886 410294 -4266 410378
rect -4886 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 -4266 410294
rect -4886 374614 -4266 410058
rect -4886 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 -4266 374614
rect -4886 374294 -4266 374378
rect -4886 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 -4266 374294
rect -4886 338614 -4266 374058
rect -4886 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 -4266 338614
rect -4886 338294 -4266 338378
rect -4886 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 -4266 338294
rect -4886 302614 -4266 338058
rect -4886 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 -4266 302614
rect -4886 302294 -4266 302378
rect -4886 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 -4266 302294
rect -4886 266614 -4266 302058
rect -4886 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 -4266 266614
rect -4886 266294 -4266 266378
rect -4886 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 -4266 266294
rect -4886 230614 -4266 266058
rect -4886 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 -4266 230614
rect -4886 230294 -4266 230378
rect -4886 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 -4266 230294
rect -4886 194614 -4266 230058
rect -4886 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 -4266 194614
rect -4886 194294 -4266 194378
rect -4886 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 -4266 194294
rect -4886 158614 -4266 194058
rect -4886 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 -4266 158614
rect -4886 158294 -4266 158378
rect -4886 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 -4266 158294
rect -4886 122614 -4266 158058
rect -4886 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 -4266 122614
rect -4886 122294 -4266 122378
rect -4886 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 -4266 122294
rect -4886 86614 -4266 122058
rect -4886 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 -4266 86614
rect -4886 86294 -4266 86378
rect -4886 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 -4266 86294
rect -4886 50614 -4266 86058
rect -4886 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 -4266 50614
rect -4886 50294 -4266 50378
rect -4886 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 -4266 50294
rect -4886 14614 -4266 50058
rect -4886 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 -4266 14614
rect -4886 14294 -4266 14378
rect -4886 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 -4266 14294
rect -4886 -3226 -4266 14058
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 694894 -3306 706202
rect -3926 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 -3306 694894
rect -3926 694574 -3306 694658
rect -3926 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 -3306 694574
rect -3926 658894 -3306 694338
rect -3926 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 -3306 658894
rect -3926 658574 -3306 658658
rect -3926 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 -3306 658574
rect -3926 622894 -3306 658338
rect -3926 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 -3306 622894
rect -3926 622574 -3306 622658
rect -3926 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 -3306 622574
rect -3926 586894 -3306 622338
rect -3926 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 -3306 586894
rect -3926 586574 -3306 586658
rect -3926 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 -3306 586574
rect -3926 550894 -3306 586338
rect -3926 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 -3306 550894
rect -3926 550574 -3306 550658
rect -3926 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 -3306 550574
rect -3926 514894 -3306 550338
rect -3926 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 -3306 514894
rect -3926 514574 -3306 514658
rect -3926 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 -3306 514574
rect -3926 478894 -3306 514338
rect -3926 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 -3306 478894
rect -3926 478574 -3306 478658
rect -3926 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 -3306 478574
rect -3926 442894 -3306 478338
rect -3926 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 -3306 442894
rect -3926 442574 -3306 442658
rect -3926 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 -3306 442574
rect -3926 406894 -3306 442338
rect -3926 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 -3306 406894
rect -3926 406574 -3306 406658
rect -3926 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 -3306 406574
rect -3926 370894 -3306 406338
rect -3926 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 -3306 370894
rect -3926 370574 -3306 370658
rect -3926 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 -3306 370574
rect -3926 334894 -3306 370338
rect -3926 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 -3306 334894
rect -3926 334574 -3306 334658
rect -3926 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 -3306 334574
rect -3926 298894 -3306 334338
rect -3926 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 -3306 298894
rect -3926 298574 -3306 298658
rect -3926 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 -3306 298574
rect -3926 262894 -3306 298338
rect -3926 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 -3306 262894
rect -3926 262574 -3306 262658
rect -3926 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 -3306 262574
rect -3926 226894 -3306 262338
rect -3926 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 -3306 226894
rect -3926 226574 -3306 226658
rect -3926 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 -3306 226574
rect -3926 190894 -3306 226338
rect -3926 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 -3306 190894
rect -3926 190574 -3306 190658
rect -3926 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 -3306 190574
rect -3926 154894 -3306 190338
rect -3926 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 -3306 154894
rect -3926 154574 -3306 154658
rect -3926 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 -3306 154574
rect -3926 118894 -3306 154338
rect -3926 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 -3306 118894
rect -3926 118574 -3306 118658
rect -3926 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 -3306 118574
rect -3926 82894 -3306 118338
rect -3926 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 -3306 82894
rect -3926 82574 -3306 82658
rect -3926 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 -3306 82574
rect -3926 46894 -3306 82338
rect -3926 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 -3306 46894
rect -3926 46574 -3306 46658
rect -3926 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 -3306 46574
rect -3926 10894 -3306 46338
rect -3926 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 -3306 10894
rect -3926 10574 -3306 10658
rect -3926 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 -3306 10574
rect -3926 -2266 -3306 10338
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 691174 -2346 705242
rect -2966 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 -2346 691174
rect -2966 690854 -2346 690938
rect -2966 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 -2346 690854
rect -2966 655174 -2346 690618
rect -2966 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 -2346 655174
rect -2966 654854 -2346 654938
rect -2966 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 -2346 654854
rect -2966 619174 -2346 654618
rect -2966 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 -2346 619174
rect -2966 618854 -2346 618938
rect -2966 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 -2346 618854
rect -2966 583174 -2346 618618
rect -2966 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 -2346 583174
rect -2966 582854 -2346 582938
rect -2966 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 -2346 582854
rect -2966 547174 -2346 582618
rect -2966 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 -2346 547174
rect -2966 546854 -2346 546938
rect -2966 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 -2346 546854
rect -2966 511174 -2346 546618
rect -2966 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 -2346 511174
rect -2966 510854 -2346 510938
rect -2966 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 -2346 510854
rect -2966 475174 -2346 510618
rect -2966 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 -2346 475174
rect -2966 474854 -2346 474938
rect -2966 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 -2346 474854
rect -2966 439174 -2346 474618
rect -2966 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 -2346 439174
rect -2966 438854 -2346 438938
rect -2966 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 -2346 438854
rect -2966 403174 -2346 438618
rect -2966 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 -2346 403174
rect -2966 402854 -2346 402938
rect -2966 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 -2346 402854
rect -2966 367174 -2346 402618
rect -2966 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 -2346 367174
rect -2966 366854 -2346 366938
rect -2966 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 -2346 366854
rect -2966 331174 -2346 366618
rect -2966 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 -2346 331174
rect -2966 330854 -2346 330938
rect -2966 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 -2346 330854
rect -2966 295174 -2346 330618
rect -2966 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 -2346 295174
rect -2966 294854 -2346 294938
rect -2966 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 -2346 294854
rect -2966 259174 -2346 294618
rect -2966 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 -2346 259174
rect -2966 258854 -2346 258938
rect -2966 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 -2346 258854
rect -2966 223174 -2346 258618
rect -2966 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 -2346 223174
rect -2966 222854 -2346 222938
rect -2966 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 -2346 222854
rect -2966 187174 -2346 222618
rect -2966 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 -2346 187174
rect -2966 186854 -2346 186938
rect -2966 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 -2346 186854
rect -2966 151174 -2346 186618
rect -2966 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 -2346 151174
rect -2966 150854 -2346 150938
rect -2966 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 -2346 150854
rect -2966 115174 -2346 150618
rect -2966 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 -2346 115174
rect -2966 114854 -2346 114938
rect -2966 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 -2346 114854
rect -2966 79174 -2346 114618
rect -2966 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 -2346 79174
rect -2966 78854 -2346 78938
rect -2966 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 -2346 78854
rect -2966 43174 -2346 78618
rect -2966 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 -2346 43174
rect -2966 42854 -2346 42938
rect -2966 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 -2346 42854
rect -2966 7174 -2346 42618
rect -2966 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 -2346 7174
rect -2966 6854 -2346 6938
rect -2966 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 -2346 6854
rect -2966 -1306 -2346 6618
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 711590
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 5514 705798 6134 711590
rect 5514 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 6134 705798
rect 5514 705478 6134 705562
rect 5514 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 6134 705478
rect 5514 691174 6134 705242
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 2819 566948 2885 566949
rect 2819 566884 2820 566948
rect 2884 566884 2885 566948
rect 2819 566883 2885 566884
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 2822 398173 2882 566883
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 3371 462636 3437 462637
rect 3371 462572 3372 462636
rect 3436 462572 3437 462636
rect 3371 462571 3437 462572
rect 2819 398172 2885 398173
rect 2819 398108 2820 398172
rect 2884 398108 2885 398172
rect 2819 398107 2885 398108
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 3374 356013 3434 462571
rect 3739 449580 3805 449581
rect 3739 449516 3740 449580
rect 3804 449516 3805 449580
rect 3739 449515 3805 449516
rect 3555 397492 3621 397493
rect 3555 397428 3556 397492
rect 3620 397428 3621 397492
rect 3555 397427 3621 397428
rect 3371 356012 3437 356013
rect 3371 355948 3372 356012
rect 3436 355948 3437 356012
rect 3371 355947 3437 355948
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 3558 326365 3618 397427
rect 3742 382941 3802 449515
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 3923 410548 3989 410549
rect 3923 410484 3924 410548
rect 3988 410484 3989 410548
rect 3923 410483 3989 410484
rect 3739 382940 3805 382941
rect 3739 382876 3740 382940
rect 3804 382876 3805 382940
rect 3739 382875 3805 382876
rect 3926 353973 3986 410483
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 3923 353972 3989 353973
rect 3923 353908 3924 353972
rect 3988 353908 3989 353972
rect 3923 353907 3989 353908
rect 4107 345404 4173 345405
rect 4107 345340 4108 345404
rect 4172 345340 4173 345404
rect 4107 345339 4173 345340
rect 4110 338741 4170 345339
rect 4107 338740 4173 338741
rect 4107 338676 4108 338740
rect 4172 338676 4173 338740
rect 4107 338675 4173 338676
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 3555 326364 3621 326365
rect 3555 326300 3556 326364
rect 3620 326300 3621 326364
rect 3555 326299 3621 326300
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 3371 293180 3437 293181
rect 3371 293116 3372 293180
rect 3436 293116 3437 293180
rect 3371 293115 3437 293116
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 3374 228309 3434 293115
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 3555 241092 3621 241093
rect 3555 241028 3556 241092
rect 3620 241028 3621 241092
rect 3555 241027 3621 241028
rect 3371 228308 3437 228309
rect 3371 228244 3372 228308
rect 3436 228244 3437 228308
rect 3371 228243 3437 228244
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 3558 218653 3618 241027
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 3555 218652 3621 218653
rect 3555 218588 3556 218652
rect 3620 218588 3621 218652
rect 3555 218587 3621 218588
rect 3371 188868 3437 188869
rect 3371 188804 3372 188868
rect 3436 188804 3437 188868
rect 3371 188803 3437 188804
rect 3374 185605 3434 188803
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 3371 185604 3437 185605
rect 3371 185540 3372 185604
rect 3436 185540 3437 185604
rect 3371 185539 3437 185540
rect 3371 184516 3437 184517
rect 3371 184452 3372 184516
rect 3436 184452 3437 184516
rect 3371 184451 3437 184452
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 3374 136781 3434 184451
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 3371 136780 3437 136781
rect 3371 136716 3372 136780
rect 3436 136716 3437 136780
rect 3371 136715 3437 136716
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 3371 113252 3437 113253
rect 3371 113188 3372 113252
rect 3436 113188 3437 113252
rect 3371 113187 3437 113188
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 3374 19413 3434 113187
rect 3555 86324 3621 86325
rect 3555 86260 3556 86324
rect 3620 86260 3621 86324
rect 3555 86259 3621 86260
rect 3558 84693 3618 86259
rect 3555 84692 3621 84693
rect 3555 84628 3556 84692
rect 3620 84628 3621 84692
rect 3555 84627 3621 84628
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 3371 19412 3437 19413
rect 3371 19348 3372 19412
rect 3436 19348 3437 19412
rect 3371 19347 3437 19348
rect 4107 7716 4173 7717
rect 4107 7652 4108 7716
rect 4172 7652 4173 7716
rect 4107 7651 4173 7652
rect 4110 6493 4170 7651
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 4107 6492 4173 6493
rect 4107 6428 4108 6492
rect 4172 6428 4173 6492
rect 4107 6427 4173 6428
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 1794 -7654 2414 -902
rect 5514 -1306 6134 6618
rect 5514 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 6134 -1306
rect 5514 -1626 6134 -1542
rect 5514 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 6134 -1626
rect 5514 -7654 6134 -1862
rect 9234 706758 9854 711590
rect 9234 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 9854 706758
rect 9234 706438 9854 706522
rect 9234 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 9854 706438
rect 9234 694894 9854 706202
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 -2266 9854 10338
rect 9234 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 9854 -2266
rect 9234 -2586 9854 -2502
rect 9234 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 9854 -2586
rect 9234 -7654 9854 -2822
rect 12954 707718 13574 711590
rect 12954 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 13574 707718
rect 12954 707398 13574 707482
rect 12954 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 13574 707398
rect 12954 698614 13574 707162
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 16674 708678 17294 711590
rect 16674 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 17294 708678
rect 16674 708358 17294 708442
rect 16674 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 17294 708358
rect 16674 666334 17294 708122
rect 16674 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 17294 666334
rect 16674 666014 17294 666098
rect 16674 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 17294 666014
rect 15699 658204 15765 658205
rect 15699 658140 15700 658204
rect 15764 658140 15765 658204
rect 15699 658139 15765 658140
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 15702 192541 15762 658139
rect 16674 630334 17294 665778
rect 16674 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 17294 630334
rect 16674 630014 17294 630098
rect 16674 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 17294 630014
rect 16674 594334 17294 629778
rect 16674 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 17294 594334
rect 16674 594014 17294 594098
rect 16674 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 17294 594014
rect 16674 558334 17294 593778
rect 16674 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 17294 558334
rect 16674 558014 17294 558098
rect 16674 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 17294 558014
rect 16674 522334 17294 557778
rect 20394 709638 21014 711590
rect 20394 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 21014 709638
rect 20394 709318 21014 709402
rect 20394 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 21014 709318
rect 20394 670054 21014 709082
rect 20394 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 21014 670054
rect 20394 669734 21014 669818
rect 20394 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 21014 669734
rect 20394 634054 21014 669498
rect 20394 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 21014 634054
rect 20394 633734 21014 633818
rect 20394 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 21014 633734
rect 20394 598054 21014 633498
rect 20394 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 21014 598054
rect 20394 597734 21014 597818
rect 20394 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 21014 597734
rect 20394 562054 21014 597498
rect 20394 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 21014 562054
rect 20394 561734 21014 561818
rect 20394 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 21014 561734
rect 18459 553892 18525 553893
rect 18459 553828 18460 553892
rect 18524 553828 18525 553892
rect 18459 553827 18525 553828
rect 16674 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 17294 522334
rect 16674 522014 17294 522098
rect 16674 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 17294 522014
rect 16674 486334 17294 521778
rect 16674 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 17294 486334
rect 16674 486014 17294 486098
rect 16674 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 17294 486014
rect 16674 450334 17294 485778
rect 16674 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 17294 450334
rect 16674 450014 17294 450098
rect 16674 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 17294 450014
rect 16674 414334 17294 449778
rect 16674 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 17294 414334
rect 16674 414014 17294 414098
rect 16674 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 17294 414014
rect 16674 378334 17294 413778
rect 16674 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 17294 378334
rect 16674 378014 17294 378098
rect 16674 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 17294 378014
rect 16674 342334 17294 377778
rect 16674 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 17294 342334
rect 16674 342014 17294 342098
rect 16674 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 17294 342014
rect 16674 306334 17294 341778
rect 16674 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 17294 306334
rect 16674 306014 17294 306098
rect 16674 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 17294 306014
rect 16674 270334 17294 305778
rect 16674 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 17294 270334
rect 16674 270014 17294 270098
rect 16674 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 17294 270014
rect 16674 234334 17294 269778
rect 16674 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 17294 234334
rect 16674 234014 17294 234098
rect 16674 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 17294 234014
rect 16674 198334 17294 233778
rect 16674 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 17294 198334
rect 16674 198014 17294 198098
rect 16674 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 17294 198014
rect 15699 192540 15765 192541
rect 15699 192476 15700 192540
rect 15764 192476 15765 192540
rect 15699 192475 15765 192476
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 -3226 13574 14058
rect 12954 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 13574 -3226
rect 12954 -3546 13574 -3462
rect 12954 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 13574 -3546
rect 12954 -7654 13574 -3782
rect 16674 162334 17294 197778
rect 18462 193901 18522 553827
rect 20394 526054 21014 561498
rect 20394 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 21014 526054
rect 20394 525734 21014 525818
rect 20394 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 21014 525734
rect 20394 490054 21014 525498
rect 24114 710598 24734 711590
rect 24114 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 24734 710598
rect 24114 710278 24734 710362
rect 24114 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 24734 710278
rect 24114 673774 24734 710042
rect 24114 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 24734 673774
rect 24114 673454 24734 673538
rect 24114 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 24734 673454
rect 24114 637774 24734 673218
rect 24114 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 24734 637774
rect 24114 637454 24734 637538
rect 24114 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 24734 637454
rect 24114 601774 24734 637218
rect 27834 711558 28454 711590
rect 27834 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 28454 711558
rect 27834 711238 28454 711322
rect 27834 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 28454 711238
rect 27834 677494 28454 711002
rect 27834 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 28454 677494
rect 27834 677174 28454 677258
rect 27834 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 28454 677174
rect 27834 641494 28454 676938
rect 37794 704838 38414 711590
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 30419 671260 30485 671261
rect 30419 671196 30420 671260
rect 30484 671196 30485 671260
rect 30419 671195 30485 671196
rect 27834 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 28454 641494
rect 27834 641174 28454 641258
rect 27834 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 28454 641174
rect 26739 606116 26805 606117
rect 26739 606052 26740 606116
rect 26804 606052 26805 606116
rect 26739 606051 26805 606052
rect 24114 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 24734 601774
rect 24114 601454 24734 601538
rect 24114 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 24734 601454
rect 24114 565774 24734 601218
rect 24114 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 24734 565774
rect 24114 565454 24734 565538
rect 24114 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 24734 565454
rect 24114 529774 24734 565218
rect 24114 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 24734 529774
rect 24114 529454 24734 529538
rect 24114 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 24734 529454
rect 22691 501804 22757 501805
rect 22691 501740 22692 501804
rect 22756 501740 22757 501804
rect 22691 501739 22757 501740
rect 20394 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 21014 490054
rect 20394 489734 21014 489818
rect 20394 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 21014 489734
rect 20394 454054 21014 489498
rect 20394 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 21014 454054
rect 20394 453734 21014 453818
rect 20394 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 21014 453734
rect 20394 418054 21014 453498
rect 20394 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 21014 418054
rect 20394 417734 21014 417818
rect 20394 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 21014 417734
rect 20394 382054 21014 417498
rect 20394 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 21014 382054
rect 20394 381734 21014 381818
rect 20394 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 21014 381734
rect 20394 346054 21014 381498
rect 20394 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 21014 346054
rect 20394 345734 21014 345818
rect 20394 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 21014 345734
rect 20394 310054 21014 345498
rect 20394 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 21014 310054
rect 20394 309734 21014 309818
rect 20394 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 21014 309734
rect 20394 274054 21014 309498
rect 20394 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 21014 274054
rect 20394 273734 21014 273818
rect 20394 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 21014 273734
rect 20394 238054 21014 273498
rect 20394 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 21014 238054
rect 20394 237734 21014 237818
rect 20394 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 21014 237734
rect 20394 202054 21014 237498
rect 20394 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 21014 202054
rect 20394 201734 21014 201818
rect 20394 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 21014 201734
rect 18459 193900 18525 193901
rect 18459 193836 18460 193900
rect 18524 193836 18525 193900
rect 18459 193835 18525 193836
rect 16674 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 17294 162334
rect 16674 162014 17294 162098
rect 16674 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 17294 162014
rect 16674 126334 17294 161778
rect 16674 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 17294 126334
rect 16674 126014 17294 126098
rect 16674 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 17294 126014
rect 16674 90334 17294 125778
rect 16674 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 17294 90334
rect 16674 90014 17294 90098
rect 16674 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 17294 90014
rect 16674 54334 17294 89778
rect 16674 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 17294 54334
rect 16674 54014 17294 54098
rect 16674 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 17294 54014
rect 16674 18334 17294 53778
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 -4186 17294 17778
rect 16674 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 17294 -4186
rect 16674 -4506 17294 -4422
rect 16674 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 17294 -4506
rect 16674 -7654 17294 -4742
rect 20394 166054 21014 201498
rect 22694 188325 22754 501739
rect 24114 493774 24734 529218
rect 26003 528188 26069 528189
rect 26003 528124 26004 528188
rect 26068 528124 26069 528188
rect 26003 528123 26069 528124
rect 24114 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 24734 493774
rect 24114 493454 24734 493538
rect 24114 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 24734 493454
rect 24114 457774 24734 493218
rect 24114 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 24734 457774
rect 24114 457454 24734 457538
rect 24114 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 24734 457454
rect 24114 421774 24734 457218
rect 26006 452437 26066 528123
rect 26003 452436 26069 452437
rect 26003 452372 26004 452436
rect 26068 452372 26069 452436
rect 26003 452371 26069 452372
rect 24114 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 24734 421774
rect 24114 421454 24734 421538
rect 24114 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 24734 421454
rect 24114 385774 24734 421218
rect 24114 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 24734 385774
rect 24114 385454 24734 385538
rect 24114 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 24734 385454
rect 24114 349774 24734 385218
rect 24114 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 24734 349774
rect 24114 349454 24734 349538
rect 24114 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 24734 349454
rect 24114 313774 24734 349218
rect 24114 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 24734 313774
rect 24114 313454 24734 313538
rect 24114 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 24734 313454
rect 24114 277774 24734 313218
rect 24114 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 24734 277774
rect 24114 277454 24734 277538
rect 24114 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 24734 277454
rect 24114 241774 24734 277218
rect 24114 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 24734 241774
rect 24114 241454 24734 241538
rect 24114 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 24734 241454
rect 24114 205774 24734 241218
rect 24114 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 24734 205774
rect 24114 205454 24734 205538
rect 24114 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 24734 205454
rect 22691 188324 22757 188325
rect 22691 188260 22692 188324
rect 22756 188260 22757 188324
rect 22691 188259 22757 188260
rect 20394 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 21014 166054
rect 20394 165734 21014 165818
rect 20394 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 21014 165734
rect 20394 130054 21014 165498
rect 20394 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 21014 130054
rect 20394 129734 21014 129818
rect 20394 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 21014 129734
rect 20394 94054 21014 129498
rect 20394 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 21014 94054
rect 20394 93734 21014 93818
rect 20394 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 21014 93734
rect 20394 58054 21014 93498
rect 20394 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 21014 58054
rect 20394 57734 21014 57818
rect 20394 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 21014 57734
rect 20394 22054 21014 57498
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 -5146 21014 21498
rect 20394 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 21014 -5146
rect 20394 -5466 21014 -5382
rect 20394 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 21014 -5466
rect 20394 -7654 21014 -5702
rect 24114 169774 24734 205218
rect 26742 191045 26802 606051
rect 27834 605494 28454 640938
rect 29131 619172 29197 619173
rect 29131 619108 29132 619172
rect 29196 619108 29197 619172
rect 29131 619107 29197 619108
rect 27834 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 28454 605494
rect 27834 605174 28454 605258
rect 27834 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 28454 605174
rect 27834 569494 28454 604938
rect 27834 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 28454 569494
rect 27834 569174 28454 569258
rect 27834 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 28454 569174
rect 27475 545732 27541 545733
rect 27475 545668 27476 545732
rect 27540 545668 27541 545732
rect 27475 545667 27541 545668
rect 27478 487253 27538 545667
rect 27834 533494 28454 568938
rect 28763 543828 28829 543829
rect 28763 543764 28764 543828
rect 28828 543764 28829 543828
rect 28763 543763 28829 543764
rect 27834 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 28454 533494
rect 27834 533174 28454 533258
rect 27834 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 28454 533174
rect 27834 497494 28454 532938
rect 27834 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 28454 497494
rect 27834 497174 28454 497258
rect 27834 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 28454 497174
rect 27475 487252 27541 487253
rect 27475 487188 27476 487252
rect 27540 487188 27541 487252
rect 27475 487187 27541 487188
rect 27834 461494 28454 496938
rect 27834 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 28454 461494
rect 27834 461174 28454 461258
rect 27834 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 28454 461174
rect 27834 425494 28454 460938
rect 28766 451893 28826 543763
rect 29134 542333 29194 619107
rect 30051 552260 30117 552261
rect 30051 552196 30052 552260
rect 30116 552196 30117 552260
rect 30051 552195 30117 552196
rect 29867 546548 29933 546549
rect 29867 546484 29868 546548
rect 29932 546484 29933 546548
rect 29867 546483 29933 546484
rect 29131 542332 29197 542333
rect 29131 542268 29132 542332
rect 29196 542268 29197 542332
rect 29131 542267 29197 542268
rect 29683 541108 29749 541109
rect 29683 541044 29684 541108
rect 29748 541044 29749 541108
rect 29683 541043 29749 541044
rect 29686 486165 29746 541043
rect 29683 486164 29749 486165
rect 29683 486100 29684 486164
rect 29748 486100 29749 486164
rect 29683 486099 29749 486100
rect 29870 485621 29930 546483
rect 29867 485620 29933 485621
rect 29867 485556 29868 485620
rect 29932 485556 29933 485620
rect 29867 485555 29933 485556
rect 30054 485077 30114 552195
rect 30235 548452 30301 548453
rect 30235 548388 30236 548452
rect 30300 548388 30301 548452
rect 30235 548387 30301 548388
rect 30051 485076 30117 485077
rect 30051 485012 30052 485076
rect 30116 485012 30117 485076
rect 30051 485011 30117 485012
rect 28763 451892 28829 451893
rect 28763 451828 28764 451892
rect 28828 451828 28829 451892
rect 28763 451827 28829 451828
rect 27834 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 28454 425494
rect 27834 425174 28454 425258
rect 27834 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 28454 425174
rect 27834 389494 28454 424938
rect 30238 414901 30298 548387
rect 30422 514861 30482 671195
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 31523 639436 31589 639437
rect 31523 639372 31524 639436
rect 31588 639372 31589 639436
rect 31523 639371 31589 639372
rect 30971 554844 31037 554845
rect 30971 554780 30972 554844
rect 31036 554780 31037 554844
rect 30971 554779 31037 554780
rect 30419 514860 30485 514861
rect 30419 514796 30420 514860
rect 30484 514796 30485 514860
rect 30419 514795 30485 514796
rect 30974 488341 31034 554779
rect 31339 537708 31405 537709
rect 31339 537644 31340 537708
rect 31404 537644 31405 537708
rect 31339 537643 31405 537644
rect 31155 514996 31221 514997
rect 31155 514932 31156 514996
rect 31220 514932 31221 514996
rect 31155 514931 31221 514932
rect 30971 488340 31037 488341
rect 30971 488276 30972 488340
rect 31036 488276 31037 488340
rect 30971 488275 31037 488276
rect 30235 414900 30301 414901
rect 30235 414836 30236 414900
rect 30300 414836 30301 414900
rect 30235 414835 30301 414836
rect 27834 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 28454 389494
rect 27834 389174 28454 389258
rect 27834 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 28454 389174
rect 27834 353494 28454 388938
rect 31158 354653 31218 514931
rect 31342 448085 31402 537643
rect 31526 450805 31586 639371
rect 34283 637940 34349 637941
rect 34283 637876 34284 637940
rect 34348 637876 34349 637940
rect 34283 637875 34349 637876
rect 32995 637260 33061 637261
rect 32995 637196 32996 637260
rect 33060 637196 33061 637260
rect 32995 637195 33061 637196
rect 32811 557564 32877 557565
rect 32811 557500 32812 557564
rect 32876 557500 32877 557564
rect 32811 557499 32877 557500
rect 32443 550764 32509 550765
rect 32443 550700 32444 550764
rect 32508 550700 32509 550764
rect 32443 550699 32509 550700
rect 32446 495957 32506 550699
rect 32627 541924 32693 541925
rect 32627 541860 32628 541924
rect 32692 541860 32693 541924
rect 32627 541859 32693 541860
rect 32443 495956 32509 495957
rect 32443 495892 32444 495956
rect 32508 495892 32509 495956
rect 32443 495891 32509 495892
rect 31523 450804 31589 450805
rect 31523 450740 31524 450804
rect 31588 450740 31589 450804
rect 31523 450739 31589 450740
rect 31339 448084 31405 448085
rect 31339 448020 31340 448084
rect 31404 448020 31405 448084
rect 31339 448019 31405 448020
rect 32630 440469 32690 541859
rect 32814 441557 32874 557499
rect 32998 449173 33058 637195
rect 33915 554300 33981 554301
rect 33915 554236 33916 554300
rect 33980 554236 33981 554300
rect 33915 554235 33981 554236
rect 33731 539612 33797 539613
rect 33731 539548 33732 539612
rect 33796 539548 33797 539612
rect 33731 539547 33797 539548
rect 33734 484533 33794 539547
rect 33731 484532 33797 484533
rect 33731 484468 33732 484532
rect 33796 484468 33797 484532
rect 33731 484467 33797 484468
rect 33918 454069 33978 554235
rect 34099 546140 34165 546141
rect 34099 546076 34100 546140
rect 34164 546076 34165 546140
rect 34099 546075 34165 546076
rect 33915 454068 33981 454069
rect 33915 454004 33916 454068
rect 33980 454004 33981 454068
rect 33915 454003 33981 454004
rect 32995 449172 33061 449173
rect 32995 449108 32996 449172
rect 33060 449108 33061 449172
rect 32995 449107 33061 449108
rect 32811 441556 32877 441557
rect 32811 441492 32812 441556
rect 32876 441492 32877 441556
rect 32811 441491 32877 441492
rect 34102 441013 34162 546075
rect 34286 450261 34346 637875
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 35755 554980 35821 554981
rect 35755 554916 35756 554980
rect 35820 554916 35821 554980
rect 35755 554915 35821 554916
rect 35571 553892 35637 553893
rect 35571 553828 35572 553892
rect 35636 553828 35637 553892
rect 35571 553827 35637 553828
rect 35387 537436 35453 537437
rect 35387 537372 35388 537436
rect 35452 537372 35453 537436
rect 35387 537371 35453 537372
rect 35203 526012 35269 526013
rect 35203 525948 35204 526012
rect 35268 525948 35269 526012
rect 35203 525947 35269 525948
rect 35206 495413 35266 525947
rect 35203 495412 35269 495413
rect 35203 495348 35204 495412
rect 35268 495348 35269 495412
rect 35203 495347 35269 495348
rect 35390 489429 35450 537371
rect 35574 505205 35634 553827
rect 35571 505204 35637 505205
rect 35571 505140 35572 505204
rect 35636 505140 35637 505204
rect 35571 505139 35637 505140
rect 35758 492149 35818 554915
rect 36859 549404 36925 549405
rect 36859 549340 36860 549404
rect 36924 549340 36925 549404
rect 36859 549339 36925 549340
rect 36675 529956 36741 529957
rect 36675 529892 36676 529956
rect 36740 529892 36741 529956
rect 36675 529891 36741 529892
rect 36491 524924 36557 524925
rect 36491 524860 36492 524924
rect 36556 524860 36557 524924
rect 36491 524859 36557 524860
rect 36494 497589 36554 524859
rect 36678 501941 36738 529891
rect 36675 501940 36741 501941
rect 36675 501876 36676 501940
rect 36740 501876 36741 501940
rect 36675 501875 36741 501876
rect 36491 497588 36557 497589
rect 36491 497524 36492 497588
rect 36556 497524 36557 497588
rect 36491 497523 36557 497524
rect 35755 492148 35821 492149
rect 35755 492084 35756 492148
rect 35820 492084 35821 492148
rect 35755 492083 35821 492084
rect 35387 489428 35453 489429
rect 35387 489364 35388 489428
rect 35452 489364 35453 489428
rect 35387 489363 35453 489364
rect 36862 483989 36922 549339
rect 37043 547500 37109 547501
rect 37043 547436 37044 547500
rect 37108 547436 37109 547500
rect 37043 547435 37109 547436
rect 36859 483988 36925 483989
rect 36859 483924 36860 483988
rect 36924 483924 36925 483988
rect 36859 483923 36925 483924
rect 34283 450260 34349 450261
rect 34283 450196 34284 450260
rect 34348 450196 34349 450260
rect 34283 450195 34349 450196
rect 37046 442101 37106 547435
rect 37794 543454 38414 578898
rect 41514 705798 42134 711590
rect 41514 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 42134 705798
rect 41514 705478 42134 705562
rect 41514 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 42134 705478
rect 41514 691174 42134 705242
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 45234 706758 45854 711590
rect 45234 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 45854 706758
rect 45234 706438 45854 706522
rect 45234 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 45854 706438
rect 45234 694894 45854 706202
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 44035 648276 44101 648277
rect 44035 648212 44036 648276
rect 44100 648212 44101 648276
rect 44035 648211 44101 648212
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 40723 553620 40789 553621
rect 40723 553556 40724 553620
rect 40788 553556 40789 553620
rect 40723 553555 40789 553556
rect 39803 553484 39869 553485
rect 39803 553420 39804 553484
rect 39868 553420 39869 553484
rect 39803 553419 39869 553420
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37411 524108 37477 524109
rect 37411 524044 37412 524108
rect 37476 524044 37477 524108
rect 37411 524043 37477 524044
rect 37227 522748 37293 522749
rect 37227 522684 37228 522748
rect 37292 522684 37293 522748
rect 37227 522683 37293 522684
rect 37230 483445 37290 522683
rect 37227 483444 37293 483445
rect 37227 483380 37228 483444
rect 37292 483380 37293 483444
rect 37227 483379 37293 483380
rect 37414 442645 37474 524043
rect 37794 507454 38414 542898
rect 39435 524516 39501 524517
rect 39435 524452 39436 524516
rect 39500 524452 39501 524516
rect 39435 524451 39501 524452
rect 39251 523292 39317 523293
rect 39251 523228 39252 523292
rect 39316 523228 39317 523292
rect 39251 523227 39317 523228
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 38883 502348 38949 502349
rect 38883 502284 38884 502348
rect 38948 502284 38949 502348
rect 38883 502283 38949 502284
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37411 442644 37477 442645
rect 37411 442580 37412 442644
rect 37476 442580 37477 442644
rect 37411 442579 37477 442580
rect 37043 442100 37109 442101
rect 37043 442036 37044 442100
rect 37108 442036 37109 442100
rect 37043 442035 37109 442036
rect 34099 441012 34165 441013
rect 34099 440948 34100 441012
rect 34164 440948 34165 441012
rect 34099 440947 34165 440948
rect 32627 440468 32693 440469
rect 32627 440404 32628 440468
rect 32692 440404 32693 440468
rect 32627 440403 32693 440404
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 38886 414357 38946 502283
rect 39067 494732 39133 494733
rect 39067 494668 39068 494732
rect 39132 494668 39133 494732
rect 39067 494667 39133 494668
rect 39070 415989 39130 494667
rect 39254 494325 39314 523227
rect 39251 494324 39317 494325
rect 39251 494260 39252 494324
rect 39316 494260 39317 494324
rect 39251 494259 39317 494260
rect 39251 491196 39317 491197
rect 39251 491132 39252 491196
rect 39316 491132 39317 491196
rect 39251 491131 39317 491132
rect 39254 416533 39314 491131
rect 39438 490517 39498 524451
rect 39619 522340 39685 522341
rect 39619 522276 39620 522340
rect 39684 522276 39685 522340
rect 39619 522275 39685 522276
rect 39435 490516 39501 490517
rect 39435 490452 39436 490516
rect 39500 490452 39501 490516
rect 39435 490451 39501 490452
rect 39622 443733 39682 522275
rect 39806 501397 39866 553419
rect 40726 502485 40786 553555
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41091 525876 41157 525877
rect 41091 525812 41092 525876
rect 41156 525812 41157 525876
rect 41091 525811 41157 525812
rect 40907 520572 40973 520573
rect 40907 520508 40908 520572
rect 40972 520508 40973 520572
rect 40907 520507 40973 520508
rect 40723 502484 40789 502485
rect 40723 502420 40724 502484
rect 40788 502420 40789 502484
rect 40723 502419 40789 502420
rect 39803 501396 39869 501397
rect 39803 501332 39804 501396
rect 39868 501332 39869 501396
rect 39803 501331 39869 501332
rect 40910 494869 40970 520507
rect 40907 494868 40973 494869
rect 40907 494804 40908 494868
rect 40972 494804 40973 494868
rect 40907 494803 40973 494804
rect 41094 444821 41154 525811
rect 41275 525060 41341 525061
rect 41275 524996 41276 525060
rect 41340 524996 41341 525060
rect 41275 524995 41341 524996
rect 41278 507381 41338 524995
rect 41514 511174 42134 546618
rect 43851 530228 43917 530229
rect 43851 530164 43852 530228
rect 43916 530164 43917 530228
rect 43851 530163 43917 530164
rect 42563 528596 42629 528597
rect 42563 528532 42564 528596
rect 42628 528532 42629 528596
rect 42563 528531 42629 528532
rect 42379 524788 42445 524789
rect 42379 524724 42380 524788
rect 42444 524724 42445 524788
rect 42379 524723 42445 524724
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41275 507380 41341 507381
rect 41275 507316 41276 507380
rect 41340 507316 41341 507380
rect 41275 507315 41341 507316
rect 41275 506564 41341 506565
rect 41275 506500 41276 506564
rect 41340 506500 41341 506564
rect 41275 506499 41341 506500
rect 41091 444820 41157 444821
rect 41091 444756 41092 444820
rect 41156 444756 41157 444820
rect 41091 444755 41157 444756
rect 39619 443732 39685 443733
rect 39619 443668 39620 443732
rect 39684 443668 39685 443732
rect 39619 443667 39685 443668
rect 41278 417077 41338 506499
rect 41514 475174 42134 510618
rect 42382 502210 42442 524723
rect 42566 502350 42626 528531
rect 43483 521932 43549 521933
rect 43483 521868 43484 521932
rect 43548 521868 43549 521932
rect 43483 521867 43549 521868
rect 42566 502290 42994 502350
rect 42382 502150 42810 502210
rect 42379 498132 42445 498133
rect 42379 498068 42380 498132
rect 42444 498068 42445 498132
rect 42379 498067 42445 498068
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41275 417076 41341 417077
rect 41275 417012 41276 417076
rect 41340 417012 41341 417076
rect 41275 417011 41341 417012
rect 39251 416532 39317 416533
rect 39251 416468 39252 416532
rect 39316 416468 39317 416532
rect 39251 416467 39317 416468
rect 39067 415988 39133 415989
rect 39067 415924 39068 415988
rect 39132 415924 39133 415988
rect 39067 415923 39133 415924
rect 38883 414356 38949 414357
rect 38883 414292 38884 414356
rect 38948 414292 38949 414356
rect 38883 414291 38949 414292
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 31155 354652 31221 354653
rect 31155 354588 31156 354652
rect 31220 354588 31221 354652
rect 31155 354587 31221 354588
rect 27834 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 28454 353494
rect 27834 353174 28454 353258
rect 27834 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 28454 353174
rect 27834 317494 28454 352938
rect 27834 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 28454 317494
rect 27834 317174 28454 317258
rect 27834 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 28454 317174
rect 27834 281494 28454 316938
rect 27834 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 28454 281494
rect 27834 281174 28454 281258
rect 27834 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 28454 281174
rect 27834 245494 28454 280938
rect 27834 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 28454 245494
rect 27834 245174 28454 245258
rect 27834 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 28454 245174
rect 27834 209494 28454 244938
rect 27834 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 28454 209494
rect 27834 209174 28454 209258
rect 27834 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 28454 209174
rect 26739 191044 26805 191045
rect 26739 190980 26740 191044
rect 26804 190980 26805 191044
rect 26739 190979 26805 190980
rect 24114 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 24734 169774
rect 24114 169454 24734 169538
rect 24114 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 24734 169454
rect 24114 133774 24734 169218
rect 24114 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 24734 133774
rect 24114 133454 24734 133538
rect 24114 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 24734 133454
rect 24114 97774 24734 133218
rect 24114 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 24734 97774
rect 24114 97454 24734 97538
rect 24114 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 24734 97454
rect 24114 61774 24734 97218
rect 24114 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 24734 61774
rect 24114 61454 24734 61538
rect 24114 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 24734 61454
rect 24114 25774 24734 61218
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 -6106 24734 25218
rect 24114 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 24734 -6106
rect 24114 -6426 24734 -6342
rect 24114 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 24734 -6426
rect 24114 -7654 24734 -6662
rect 27834 173494 28454 208938
rect 27834 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 28454 173494
rect 27834 173174 28454 173258
rect 27834 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 28454 173174
rect 27834 137494 28454 172938
rect 27834 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 28454 137494
rect 27834 137174 28454 137258
rect 27834 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 28454 137174
rect 27834 101494 28454 136938
rect 27834 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 28454 101494
rect 27834 101174 28454 101258
rect 27834 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 28454 101174
rect 27834 65494 28454 100938
rect 27834 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 28454 65494
rect 27834 65174 28454 65258
rect 27834 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 28454 65174
rect 27834 29494 28454 64938
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 -7066 28454 28938
rect 27834 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 28454 -7066
rect 27834 -7386 28454 -7302
rect 27834 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 28454 -7386
rect 27834 -7654 28454 -7622
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -7654 38414 -902
rect 41514 403174 42134 438618
rect 42382 415445 42442 498067
rect 42750 497045 42810 502150
rect 42747 497044 42813 497045
rect 42747 496980 42748 497044
rect 42812 496980 42813 497044
rect 42747 496979 42813 496980
rect 42934 492690 42994 502290
rect 43486 496773 43546 521867
rect 43667 521796 43733 521797
rect 43667 521732 43668 521796
rect 43732 521732 43733 521796
rect 43667 521731 43733 521732
rect 43483 496772 43549 496773
rect 43483 496708 43484 496772
rect 43548 496708 43549 496772
rect 43483 496707 43549 496708
rect 42566 492630 42994 492690
rect 42566 491605 42626 492630
rect 42563 491604 42629 491605
rect 42563 491540 42564 491604
rect 42628 491540 42629 491604
rect 42563 491539 42629 491540
rect 42379 415444 42445 415445
rect 42379 415380 42380 415444
rect 42444 415380 42445 415444
rect 42379 415379 42445 415380
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 43670 360909 43730 521731
rect 43854 509557 43914 530163
rect 44038 518805 44098 648211
rect 45234 622894 45854 658338
rect 48954 707718 49574 711590
rect 48954 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 49574 707718
rect 48954 707398 49574 707482
rect 48954 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 49574 707398
rect 48954 698614 49574 707162
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48635 643652 48701 643653
rect 48635 643588 48636 643652
rect 48700 643588 48701 643652
rect 48635 643587 48701 643588
rect 46795 643380 46861 643381
rect 46795 643316 46796 643380
rect 46860 643316 46861 643380
rect 46795 643315 46861 643316
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 44955 526828 45021 526829
rect 44955 526764 44956 526828
rect 45020 526764 45021 526828
rect 44955 526763 45021 526764
rect 44771 525468 44837 525469
rect 44771 525404 44772 525468
rect 44836 525404 44837 525468
rect 44771 525403 44837 525404
rect 44587 523836 44653 523837
rect 44587 523772 44588 523836
rect 44652 523772 44653 523836
rect 44587 523771 44653 523772
rect 44035 518804 44101 518805
rect 44035 518740 44036 518804
rect 44100 518740 44101 518804
rect 44035 518739 44101 518740
rect 43851 509556 43917 509557
rect 43851 509492 43852 509556
rect 43916 509492 43917 509556
rect 43851 509491 43917 509492
rect 44403 494052 44469 494053
rect 44403 493988 44404 494052
rect 44468 493988 44469 494052
rect 44403 493987 44469 493988
rect 44406 413813 44466 493987
rect 44590 493237 44650 523771
rect 44587 493236 44653 493237
rect 44587 493172 44588 493236
rect 44652 493172 44653 493236
rect 44587 493171 44653 493172
rect 44774 443189 44834 525403
rect 44771 443188 44837 443189
rect 44771 443124 44772 443188
rect 44836 443124 44837 443188
rect 44771 443123 44837 443124
rect 44958 438837 45018 526763
rect 45234 514894 45854 550338
rect 46427 525196 46493 525197
rect 46427 525132 46428 525196
rect 46492 525132 46493 525196
rect 46427 525131 46493 525132
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 46430 494733 46490 525131
rect 46611 523564 46677 523565
rect 46611 523500 46612 523564
rect 46676 523500 46677 523564
rect 46611 523499 46677 523500
rect 46427 494732 46493 494733
rect 46427 494668 46428 494732
rect 46492 494668 46493 494732
rect 46427 494667 46493 494668
rect 46059 491876 46125 491877
rect 46059 491812 46060 491876
rect 46124 491812 46125 491876
rect 46059 491811 46125 491812
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 46062 475421 46122 491811
rect 46059 475420 46125 475421
rect 46059 475356 46060 475420
rect 46124 475356 46125 475420
rect 46059 475355 46125 475356
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 44955 438836 45021 438837
rect 44955 438772 44956 438836
rect 45020 438772 45021 438836
rect 44955 438771 45021 438772
rect 44403 413812 44469 413813
rect 44403 413748 44404 413812
rect 44468 413748 44469 413812
rect 44403 413747 44469 413748
rect 45234 406894 45854 442338
rect 46614 439381 46674 523499
rect 46798 458421 46858 643315
rect 47899 639708 47965 639709
rect 47899 639644 47900 639708
rect 47964 639644 47965 639708
rect 47899 639643 47965 639644
rect 47715 635356 47781 635357
rect 47715 635292 47716 635356
rect 47780 635292 47781 635356
rect 47715 635291 47781 635292
rect 47531 556204 47597 556205
rect 47531 556140 47532 556204
rect 47596 556140 47597 556204
rect 47531 556139 47597 556140
rect 46795 458420 46861 458421
rect 46795 458356 46796 458420
rect 46860 458356 46861 458420
rect 46795 458355 46861 458356
rect 47534 439925 47594 556139
rect 47718 455157 47778 635291
rect 47902 455701 47962 639643
rect 48083 636716 48149 636717
rect 48083 636652 48084 636716
rect 48148 636652 48149 636716
rect 48083 636651 48149 636652
rect 47899 455700 47965 455701
rect 47899 455636 47900 455700
rect 47964 455636 47965 455700
rect 47899 455635 47965 455636
rect 47715 455156 47781 455157
rect 47715 455092 47716 455156
rect 47780 455092 47781 455156
rect 47715 455091 47781 455092
rect 48086 451349 48146 636651
rect 48451 636580 48517 636581
rect 48451 636516 48452 636580
rect 48516 636516 48517 636580
rect 48451 636515 48517 636516
rect 48454 454613 48514 636515
rect 48638 457877 48698 643587
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 52674 708678 53294 711590
rect 52674 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 53294 708678
rect 52674 708358 53294 708442
rect 52674 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 53294 708358
rect 52674 666334 53294 708122
rect 52674 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 53294 666334
rect 52674 666014 53294 666098
rect 52674 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 53294 666014
rect 52674 630334 53294 665778
rect 56394 709638 57014 711590
rect 56394 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 57014 709638
rect 56394 709318 57014 709402
rect 56394 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 57014 709318
rect 56394 670054 57014 709082
rect 56394 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 57014 670054
rect 56394 669734 57014 669818
rect 56394 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 57014 669734
rect 54891 645420 54957 645421
rect 54891 645356 54892 645420
rect 54956 645356 54957 645420
rect 54891 645355 54957 645356
rect 52674 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 53294 630334
rect 52674 630014 53294 630098
rect 52674 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 53294 630014
rect 52674 594334 53294 629778
rect 52674 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 53294 594334
rect 52674 594014 53294 594098
rect 52674 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 53294 594014
rect 52674 558334 53294 593778
rect 52674 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 53294 558334
rect 52674 558014 53294 558098
rect 52674 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 53294 558014
rect 52315 531860 52381 531861
rect 52315 531796 52316 531860
rect 52380 531796 52381 531860
rect 52315 531795 52381 531796
rect 50843 530364 50909 530365
rect 50843 530300 50844 530364
rect 50908 530300 50909 530364
rect 50843 530299 50909 530300
rect 49739 527236 49805 527237
rect 49739 527172 49740 527236
rect 49804 527172 49805 527236
rect 49739 527171 49805 527172
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 49742 506565 49802 527171
rect 50291 520300 50357 520301
rect 50291 520236 50292 520300
rect 50356 520236 50357 520300
rect 50291 520235 50357 520236
rect 49739 506564 49805 506565
rect 49739 506500 49740 506564
rect 49804 506500 49805 506564
rect 49739 506499 49805 506500
rect 50294 482901 50354 520235
rect 50659 519620 50725 519621
rect 50659 519556 50660 519620
rect 50724 519556 50725 519620
rect 50659 519555 50725 519556
rect 50662 510645 50722 519555
rect 50659 510644 50725 510645
rect 50659 510580 50660 510644
rect 50724 510580 50725 510644
rect 50659 510579 50725 510580
rect 50291 482900 50357 482901
rect 50291 482836 50292 482900
rect 50356 482836 50357 482900
rect 50291 482835 50357 482836
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48635 457876 48701 457877
rect 48635 457812 48636 457876
rect 48700 457812 48701 457876
rect 48635 457811 48701 457812
rect 48451 454612 48517 454613
rect 48451 454548 48452 454612
rect 48516 454548 48517 454612
rect 48451 454547 48517 454548
rect 48083 451348 48149 451349
rect 48083 451284 48084 451348
rect 48148 451284 48149 451348
rect 48083 451283 48149 451284
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 47531 439924 47597 439925
rect 47531 439860 47532 439924
rect 47596 439860 47597 439924
rect 47531 439859 47597 439860
rect 46611 439380 46677 439381
rect 46611 439316 46612 439380
rect 46676 439316 46677 439380
rect 46611 439315 46677 439316
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 43667 360908 43733 360909
rect 43667 360844 43668 360908
rect 43732 360844 43733 360908
rect 43667 360843 43733 360844
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -1306 42134 6618
rect 41514 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 42134 -1306
rect 41514 -1626 42134 -1542
rect 41514 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 42134 -1626
rect 41514 -7654 42134 -1862
rect 45234 334894 45854 370338
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48083 346492 48149 346493
rect 48083 346428 48084 346492
rect 48148 346428 48149 346492
rect 48083 346427 48149 346428
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 48086 285021 48146 346427
rect 48954 338614 49574 374058
rect 50846 352613 50906 530299
rect 51211 520300 51277 520301
rect 51211 520236 51212 520300
rect 51276 520236 51277 520300
rect 51211 520235 51277 520236
rect 52131 520300 52197 520301
rect 52131 520236 52132 520300
rect 52196 520236 52197 520300
rect 52131 520235 52197 520236
rect 51214 509250 51274 520235
rect 51579 519348 51645 519349
rect 51579 519284 51580 519348
rect 51644 519284 51645 519348
rect 51579 519283 51645 519284
rect 51030 509190 51274 509250
rect 51030 503709 51090 509190
rect 51027 503708 51093 503709
rect 51027 503644 51028 503708
rect 51092 503644 51093 503708
rect 51027 503643 51093 503644
rect 51582 476237 51642 519283
rect 52134 499901 52194 520235
rect 52131 499900 52197 499901
rect 52131 499836 52132 499900
rect 52196 499836 52197 499900
rect 52131 499835 52197 499836
rect 51579 476236 51645 476237
rect 51579 476172 51580 476236
rect 51644 476172 51645 476236
rect 51579 476171 51645 476172
rect 52318 445365 52378 531795
rect 52674 522334 53294 557778
rect 53603 557700 53669 557701
rect 53603 557636 53604 557700
rect 53668 557636 53669 557700
rect 53603 557635 53669 557636
rect 52674 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 53294 522334
rect 52674 522014 53294 522098
rect 52674 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 53294 522014
rect 52674 486334 53294 521778
rect 52674 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 53294 486334
rect 52674 486014 53294 486098
rect 52674 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 53294 486014
rect 52674 450334 53294 485778
rect 52674 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 53294 450334
rect 52674 450014 53294 450098
rect 52674 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 53294 450014
rect 52315 445364 52381 445365
rect 52315 445300 52316 445364
rect 52380 445300 52381 445364
rect 52315 445299 52381 445300
rect 52674 414334 53294 449778
rect 53606 447541 53666 557635
rect 54523 554164 54589 554165
rect 54523 554100 54524 554164
rect 54588 554100 54589 554164
rect 54523 554099 54589 554100
rect 53787 529820 53853 529821
rect 53787 529756 53788 529820
rect 53852 529756 53853 529820
rect 53787 529755 53853 529756
rect 53790 513365 53850 529755
rect 53787 513364 53853 513365
rect 53787 513300 53788 513364
rect 53852 513300 53853 513364
rect 53787 513299 53853 513300
rect 54526 503573 54586 554099
rect 54707 524380 54773 524381
rect 54707 524316 54708 524380
rect 54772 524316 54773 524380
rect 54707 524315 54773 524316
rect 54523 503572 54589 503573
rect 54523 503508 54524 503572
rect 54588 503508 54589 503572
rect 54523 503507 54589 503508
rect 54339 475420 54405 475421
rect 54339 475356 54340 475420
rect 54404 475356 54405 475420
rect 54339 475355 54405 475356
rect 54342 452981 54402 475355
rect 54339 452980 54405 452981
rect 54339 452916 54340 452980
rect 54404 452916 54405 452980
rect 54339 452915 54405 452916
rect 54710 449717 54770 524315
rect 54894 456245 54954 645355
rect 55995 635900 56061 635901
rect 55995 635836 55996 635900
rect 56060 635836 56061 635900
rect 55995 635835 56061 635836
rect 55811 554980 55877 554981
rect 55811 554916 55812 554980
rect 55876 554916 55877 554980
rect 55811 554915 55877 554916
rect 55075 527236 55141 527237
rect 55075 527172 55076 527236
rect 55140 527172 55141 527236
rect 55075 527171 55141 527172
rect 54891 456244 54957 456245
rect 54891 456180 54892 456244
rect 54956 456180 54957 456244
rect 54891 456179 54957 456180
rect 54707 449716 54773 449717
rect 54707 449652 54708 449716
rect 54772 449652 54773 449716
rect 54707 449651 54773 449652
rect 53603 447540 53669 447541
rect 53603 447476 53604 447540
rect 53668 447476 53669 447540
rect 53603 447475 53669 447476
rect 52674 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 53294 414334
rect 52674 414014 53294 414098
rect 52674 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 53294 414014
rect 52674 378334 53294 413778
rect 52674 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 53294 378334
rect 52674 378014 53294 378098
rect 52674 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 53294 378014
rect 50843 352612 50909 352613
rect 50843 352548 50844 352612
rect 50908 352548 50909 352612
rect 50843 352547 50909 352548
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48083 285020 48149 285021
rect 48083 284956 48084 285020
rect 48148 284956 48149 285020
rect 48083 284955 48149 284956
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48635 254148 48701 254149
rect 48635 254084 48636 254148
rect 48700 254084 48701 254148
rect 48635 254083 48701 254084
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 48638 119373 48698 254083
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48635 119372 48701 119373
rect 48635 119308 48636 119372
rect 48700 119308 48701 119372
rect 48635 119307 48701 119308
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 46059 112436 46125 112437
rect 46059 112372 46060 112436
rect 46124 112372 46125 112436
rect 46059 112371 46125 112372
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 46062 58581 46122 112371
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 46059 58580 46125 58581
rect 46059 58516 46060 58580
rect 46124 58516 46125 58580
rect 46059 58515 46125 58516
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -2266 45854 10338
rect 45234 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 45854 -2266
rect 45234 -2586 45854 -2502
rect 45234 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 45854 -2586
rect 45234 -7654 45854 -2822
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 48954 -3226 49574 14058
rect 48954 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 49574 -3226
rect 48954 -3546 49574 -3462
rect 48954 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 49574 -3546
rect 48954 -7654 49574 -3782
rect 52674 342334 53294 377778
rect 52674 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 53294 342334
rect 52674 342014 53294 342098
rect 52674 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 53294 342014
rect 52674 306334 53294 341778
rect 52674 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 53294 306334
rect 52674 306014 53294 306098
rect 52674 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 53294 306014
rect 52674 270334 53294 305778
rect 55078 301477 55138 527171
rect 55443 520028 55509 520029
rect 55443 519964 55444 520028
rect 55508 519964 55509 520028
rect 55443 519963 55509 519964
rect 55446 503709 55506 519963
rect 55627 514044 55693 514045
rect 55627 513980 55628 514044
rect 55692 513980 55693 514044
rect 55627 513979 55693 513980
rect 55443 503708 55509 503709
rect 55443 503644 55444 503708
rect 55508 503644 55509 503708
rect 55443 503643 55509 503644
rect 55630 500717 55690 513979
rect 55627 500716 55693 500717
rect 55627 500652 55628 500716
rect 55692 500652 55693 500716
rect 55627 500651 55693 500652
rect 55814 487797 55874 554915
rect 55998 514453 56058 635835
rect 56394 634054 57014 669498
rect 56394 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 57014 634054
rect 56394 633734 57014 633818
rect 56394 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 57014 633734
rect 56394 598054 57014 633498
rect 60114 710598 60734 711590
rect 60114 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 60734 710598
rect 60114 710278 60734 710362
rect 60114 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 60734 710278
rect 60114 673774 60734 710042
rect 60114 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 60734 673774
rect 60114 673454 60734 673538
rect 60114 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 60734 673454
rect 60114 637774 60734 673218
rect 60114 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 60734 637774
rect 60114 637454 60734 637538
rect 60114 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 60734 637454
rect 60114 633233 60734 637218
rect 63834 711558 64454 711590
rect 63834 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 64454 711558
rect 63834 711238 64454 711322
rect 63834 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 64454 711238
rect 63834 677494 64454 711002
rect 63834 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 64454 677494
rect 63834 677174 64454 677258
rect 63834 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 64454 677174
rect 63834 641494 64454 676938
rect 63834 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 64454 641494
rect 63834 641174 64454 641258
rect 63834 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 64454 641174
rect 63834 634540 64454 640938
rect 73794 704838 74414 711590
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 633233 74414 650898
rect 77514 705798 78134 711590
rect 77514 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 78134 705798
rect 77514 705478 78134 705562
rect 77514 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 78134 705478
rect 77514 691174 78134 705242
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 633233 78134 654618
rect 81234 706758 81854 711590
rect 81234 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 81854 706758
rect 81234 706438 81854 706522
rect 81234 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 81854 706438
rect 81234 694894 81854 706202
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 633233 81854 658338
rect 84954 707718 85574 711590
rect 84954 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 85574 707718
rect 84954 707398 85574 707482
rect 84954 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 85574 707398
rect 84954 698614 85574 707162
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 633233 85574 662058
rect 88674 708678 89294 711590
rect 88674 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 89294 708678
rect 88674 708358 89294 708442
rect 88674 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 89294 708358
rect 88674 666334 89294 708122
rect 88674 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 89294 666334
rect 88674 666014 89294 666098
rect 88674 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 89294 666014
rect 88674 633233 89294 665778
rect 92394 709638 93014 711590
rect 92394 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 93014 709638
rect 92394 709318 93014 709402
rect 92394 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 93014 709318
rect 92394 670054 93014 709082
rect 92394 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 93014 670054
rect 92394 669734 93014 669818
rect 92394 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 93014 669734
rect 92394 634054 93014 669498
rect 92394 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 93014 634054
rect 92394 633734 93014 633818
rect 92394 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 93014 633734
rect 92394 633233 93014 633498
rect 96114 710598 96734 711590
rect 96114 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 96734 710598
rect 96114 710278 96734 710362
rect 96114 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 96734 710278
rect 96114 673774 96734 710042
rect 96114 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 96734 673774
rect 96114 673454 96734 673538
rect 96114 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 96734 673454
rect 96114 637774 96734 673218
rect 96114 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 96734 637774
rect 96114 637454 96734 637538
rect 96114 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 96734 637454
rect 96114 633233 96734 637218
rect 99834 711558 100454 711590
rect 99834 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 100454 711558
rect 99834 711238 100454 711322
rect 99834 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 100454 711238
rect 99834 677494 100454 711002
rect 99834 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 100454 677494
rect 99834 677174 100454 677258
rect 99834 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 100454 677174
rect 99834 641494 100454 676938
rect 99834 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 100454 641494
rect 99834 641174 100454 641258
rect 99834 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 100454 641174
rect 99834 633233 100454 640938
rect 109794 704838 110414 711590
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 634540 110414 650898
rect 113514 705798 114134 711590
rect 113514 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 114134 705798
rect 113514 705478 114134 705562
rect 113514 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 114134 705478
rect 113514 691174 114134 705242
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 633233 114134 654618
rect 117234 706758 117854 711590
rect 117234 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 117854 706758
rect 117234 706438 117854 706522
rect 117234 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 117854 706438
rect 117234 694894 117854 706202
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 633233 117854 658338
rect 120954 707718 121574 711590
rect 120954 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 121574 707718
rect 120954 707398 121574 707482
rect 120954 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 121574 707398
rect 120954 698614 121574 707162
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 633233 121574 662058
rect 124674 708678 125294 711590
rect 124674 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 125294 708678
rect 124674 708358 125294 708442
rect 124674 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 125294 708358
rect 124674 666334 125294 708122
rect 124674 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 125294 666334
rect 124674 666014 125294 666098
rect 124674 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 125294 666014
rect 124674 633233 125294 665778
rect 128394 709638 129014 711590
rect 128394 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 129014 709638
rect 128394 709318 129014 709402
rect 128394 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 129014 709318
rect 128394 670054 129014 709082
rect 128394 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 129014 670054
rect 128394 669734 129014 669818
rect 128394 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 129014 669734
rect 127571 634132 127637 634133
rect 127571 634068 127572 634132
rect 127636 634068 127637 634132
rect 127571 634067 127637 634068
rect 127574 633725 127634 634067
rect 128394 634054 129014 669498
rect 128394 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 129014 634054
rect 128394 633734 129014 633818
rect 127571 633724 127637 633725
rect 127571 633660 127572 633724
rect 127636 633660 127637 633724
rect 127571 633659 127637 633660
rect 128394 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 129014 633734
rect 128394 633233 129014 633498
rect 132114 710598 132734 711590
rect 132114 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 132734 710598
rect 132114 710278 132734 710362
rect 132114 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 132734 710278
rect 132114 673774 132734 710042
rect 132114 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 132734 673774
rect 132114 673454 132734 673538
rect 132114 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 132734 673454
rect 132114 637774 132734 673218
rect 132114 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 132734 637774
rect 132114 637454 132734 637538
rect 132114 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 132734 637454
rect 132114 633233 132734 637218
rect 135834 711558 136454 711590
rect 135834 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 136454 711558
rect 135834 711238 136454 711322
rect 135834 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 136454 711238
rect 135834 677494 136454 711002
rect 135834 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 136454 677494
rect 135834 677174 136454 677258
rect 135834 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 136454 677174
rect 135834 641494 136454 676938
rect 135834 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 136454 641494
rect 135834 641174 136454 641258
rect 135834 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 136454 641174
rect 57651 628828 57717 628829
rect 57651 628764 57652 628828
rect 57716 628764 57717 628828
rect 57651 628763 57717 628764
rect 56394 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 57014 598054
rect 56394 597734 57014 597818
rect 56394 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 57014 597734
rect 56394 562054 57014 597498
rect 56394 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 57014 562054
rect 56394 561734 57014 561818
rect 56394 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 57014 561734
rect 56394 526054 57014 561498
rect 57654 560285 57714 628763
rect 57835 627740 57901 627741
rect 57835 627676 57836 627740
rect 57900 627676 57901 627740
rect 57835 627675 57901 627676
rect 57651 560284 57717 560285
rect 57651 560220 57652 560284
rect 57716 560220 57717 560284
rect 57651 560219 57717 560220
rect 57838 534853 57898 627675
rect 58939 626652 59005 626653
rect 58939 626588 58940 626652
rect 59004 626588 59005 626652
rect 58939 626587 59005 626588
rect 58755 619172 58821 619173
rect 58755 619108 58756 619172
rect 58820 619108 58821 619172
rect 58755 619107 58821 619108
rect 58758 559469 58818 619107
rect 58755 559468 58821 559469
rect 58755 559404 58756 559468
rect 58820 559404 58821 559468
rect 58755 559403 58821 559404
rect 58571 554436 58637 554437
rect 58571 554372 58572 554436
rect 58636 554372 58637 554436
rect 58571 554371 58637 554372
rect 58387 542196 58453 542197
rect 58387 542132 58388 542196
rect 58452 542132 58453 542196
rect 58387 542131 58453 542132
rect 57835 534852 57901 534853
rect 57835 534788 57836 534852
rect 57900 534788 57901 534852
rect 57835 534787 57901 534788
rect 56394 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 57014 526054
rect 56394 525734 57014 525818
rect 56394 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 57014 525734
rect 55995 514452 56061 514453
rect 55995 514388 55996 514452
rect 56060 514388 56061 514452
rect 55995 514387 56061 514388
rect 55995 497180 56061 497181
rect 55995 497116 55996 497180
rect 56060 497116 56061 497180
rect 55995 497115 56061 497116
rect 55811 487796 55877 487797
rect 55811 487732 55812 487796
rect 55876 487732 55877 487796
rect 55811 487731 55877 487732
rect 55998 478957 56058 497115
rect 56394 490054 57014 525498
rect 57651 523156 57717 523157
rect 57651 523092 57652 523156
rect 57716 523092 57717 523156
rect 57651 523091 57717 523092
rect 57654 510645 57714 523091
rect 57835 520980 57901 520981
rect 57835 520916 57836 520980
rect 57900 520916 57901 520980
rect 57835 520915 57901 520916
rect 57651 510644 57717 510645
rect 57651 510580 57652 510644
rect 57716 510580 57717 510644
rect 57651 510579 57717 510580
rect 57651 508604 57717 508605
rect 57651 508540 57652 508604
rect 57716 508540 57717 508604
rect 57651 508539 57717 508540
rect 57654 505749 57714 508539
rect 57651 505748 57717 505749
rect 57651 505684 57652 505748
rect 57716 505684 57717 505748
rect 57651 505683 57717 505684
rect 57467 505340 57533 505341
rect 57467 505276 57468 505340
rect 57532 505276 57533 505340
rect 57467 505275 57533 505276
rect 57470 499221 57530 505275
rect 57467 499220 57533 499221
rect 57467 499156 57468 499220
rect 57532 499156 57533 499220
rect 57467 499155 57533 499156
rect 57651 498948 57717 498949
rect 57651 498884 57652 498948
rect 57716 498884 57717 498948
rect 57651 498883 57717 498884
rect 57654 496501 57714 498883
rect 57651 496500 57717 496501
rect 57651 496436 57652 496500
rect 57716 496436 57717 496500
rect 57651 496435 57717 496436
rect 57283 494732 57349 494733
rect 57283 494668 57284 494732
rect 57348 494668 57349 494732
rect 57283 494667 57349 494668
rect 56394 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 57014 490054
rect 56394 489734 57014 489818
rect 56394 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 57014 489734
rect 55995 478956 56061 478957
rect 55995 478892 55996 478956
rect 56060 478892 56061 478956
rect 55995 478891 56061 478892
rect 56394 454054 57014 489498
rect 56394 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 57014 454054
rect 56394 453734 57014 453818
rect 56394 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 57014 453734
rect 56394 418054 57014 453498
rect 57286 448629 57346 494667
rect 57283 448628 57349 448629
rect 57283 448564 57284 448628
rect 57348 448564 57349 448628
rect 57283 448563 57349 448564
rect 57838 444277 57898 520915
rect 58390 446453 58450 542131
rect 58574 503029 58634 554371
rect 58942 538117 59002 626587
rect 59123 620260 59189 620261
rect 59123 620196 59124 620260
rect 59188 620196 59189 620260
rect 59123 620195 59189 620196
rect 59126 560285 59186 620195
rect 79568 619174 79888 619206
rect 79568 618938 79610 619174
rect 79846 618938 79888 619174
rect 79568 618854 79888 618938
rect 79568 618618 79610 618854
rect 79846 618618 79888 618854
rect 79568 618586 79888 618618
rect 110288 619174 110608 619206
rect 110288 618938 110330 619174
rect 110566 618938 110608 619174
rect 110288 618854 110608 618938
rect 110288 618618 110330 618854
rect 110566 618618 110608 618854
rect 110288 618586 110608 618618
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 125648 615454 125968 615486
rect 125648 615218 125690 615454
rect 125926 615218 125968 615454
rect 125648 615134 125968 615218
rect 125648 614898 125690 615134
rect 125926 614898 125968 615134
rect 125648 614866 125968 614898
rect 59675 610468 59741 610469
rect 59675 610404 59676 610468
rect 59740 610404 59741 610468
rect 59675 610403 59741 610404
rect 59123 560284 59189 560285
rect 59123 560220 59124 560284
rect 59188 560220 59189 560284
rect 59123 560219 59189 560220
rect 59678 551581 59738 610403
rect 135834 605494 136454 640938
rect 135834 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 136454 605494
rect 135834 605174 136454 605258
rect 135834 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 136454 605174
rect 79568 583174 79888 583206
rect 79568 582938 79610 583174
rect 79846 582938 79888 583174
rect 79568 582854 79888 582938
rect 79568 582618 79610 582854
rect 79846 582618 79888 582854
rect 79568 582586 79888 582618
rect 110288 583174 110608 583206
rect 110288 582938 110330 583174
rect 110566 582938 110608 583174
rect 110288 582854 110608 582938
rect 110288 582618 110330 582854
rect 110566 582618 110608 582854
rect 110288 582586 110608 582618
rect 64208 579454 64528 579486
rect 64208 579218 64250 579454
rect 64486 579218 64528 579454
rect 64208 579134 64528 579218
rect 64208 578898 64250 579134
rect 64486 578898 64528 579134
rect 64208 578866 64528 578898
rect 94928 579454 95248 579486
rect 94928 579218 94970 579454
rect 95206 579218 95248 579454
rect 94928 579134 95248 579218
rect 94928 578898 94970 579134
rect 95206 578898 95248 579134
rect 94928 578866 95248 578898
rect 125648 579454 125968 579486
rect 125648 579218 125690 579454
rect 125926 579218 125968 579454
rect 125648 579134 125968 579218
rect 125648 578898 125690 579134
rect 125926 578898 125968 579134
rect 125648 578866 125968 578898
rect 135834 569494 136454 604938
rect 135834 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 136454 569494
rect 135834 569174 136454 569258
rect 135834 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 136454 569174
rect 59859 559060 59925 559061
rect 59859 558996 59860 559060
rect 59924 558996 59925 559060
rect 59859 558995 59925 558996
rect 59675 551580 59741 551581
rect 59675 551516 59676 551580
rect 59740 551516 59741 551580
rect 59675 551515 59741 551516
rect 59123 550900 59189 550901
rect 59123 550836 59124 550900
rect 59188 550836 59189 550900
rect 59123 550835 59189 550836
rect 58939 538116 59005 538117
rect 58939 538052 58940 538116
rect 59004 538052 59005 538116
rect 58939 538051 59005 538052
rect 58755 535804 58821 535805
rect 58755 535740 58756 535804
rect 58820 535740 58821 535804
rect 58755 535739 58821 535740
rect 58571 503028 58637 503029
rect 58571 502964 58572 503028
rect 58636 502964 58637 503028
rect 58571 502963 58637 502964
rect 58758 453525 58818 535739
rect 58755 453524 58821 453525
rect 58755 453460 58756 453524
rect 58820 453460 58821 453524
rect 58755 453459 58821 453460
rect 59126 446997 59186 550835
rect 59675 520300 59741 520301
rect 59675 520236 59676 520300
rect 59740 520236 59741 520300
rect 59675 520235 59741 520236
rect 59678 493781 59738 520235
rect 59675 493780 59741 493781
rect 59675 493716 59676 493780
rect 59740 493716 59741 493780
rect 59675 493715 59741 493716
rect 59123 446996 59189 446997
rect 59123 446932 59124 446996
rect 59188 446932 59189 446996
rect 59123 446931 59189 446932
rect 58387 446452 58453 446453
rect 58387 446388 58388 446452
rect 58452 446388 58453 446452
rect 58387 446387 58453 446388
rect 59862 445909 59922 558995
rect 60114 529774 60734 558575
rect 73794 543454 74414 558575
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 61883 530500 61949 530501
rect 61883 530436 61884 530500
rect 61948 530436 61949 530500
rect 61883 530435 61949 530436
rect 60114 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 60734 529774
rect 60114 529454 60734 529538
rect 60114 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 60734 529454
rect 61331 529412 61397 529413
rect 61331 529348 61332 529412
rect 61396 529348 61397 529412
rect 61331 529347 61397 529348
rect 60114 493774 60734 529218
rect 61334 520301 61394 529347
rect 61886 520301 61946 530435
rect 61331 520300 61397 520301
rect 61331 520236 61332 520300
rect 61396 520236 61397 520300
rect 61331 520235 61397 520236
rect 61883 520300 61949 520301
rect 61883 520236 61884 520300
rect 61948 520236 61949 520300
rect 61883 520235 61949 520236
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 60114 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 60734 493774
rect 60114 493454 60734 493538
rect 60114 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 60734 493454
rect 60114 457774 60734 493218
rect 64208 471454 64528 471486
rect 64208 471218 64250 471454
rect 64486 471218 64528 471454
rect 64208 471134 64528 471218
rect 64208 470898 64250 471134
rect 64486 470898 64528 471134
rect 64208 470866 64528 470898
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 60114 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 60734 457774
rect 60114 457454 60734 457538
rect 60114 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 60734 457454
rect 59859 445908 59925 445909
rect 59859 445844 59860 445908
rect 59924 445844 59925 445908
rect 59859 445843 59925 445844
rect 57835 444276 57901 444277
rect 57835 444212 57836 444276
rect 57900 444212 57901 444276
rect 57835 444211 57901 444212
rect 56394 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 57014 418054
rect 56394 417734 57014 417818
rect 56394 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 57014 417734
rect 56394 382054 57014 417498
rect 56394 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 57014 382054
rect 56394 381734 57014 381818
rect 56394 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 57014 381734
rect 56394 346054 57014 381498
rect 56394 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 57014 346054
rect 56394 345734 57014 345818
rect 56394 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 57014 345734
rect 56394 310054 57014 345498
rect 56394 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 57014 310054
rect 56394 309734 57014 309818
rect 56394 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 57014 309734
rect 55075 301476 55141 301477
rect 55075 301412 55076 301476
rect 55140 301412 55141 301476
rect 55075 301411 55141 301412
rect 54208 291454 54528 291486
rect 54208 291218 54250 291454
rect 54486 291218 54528 291454
rect 54208 291134 54528 291218
rect 54208 290898 54250 291134
rect 54486 290898 54528 291134
rect 54208 290866 54528 290898
rect 52674 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 53294 270334
rect 52674 270014 53294 270098
rect 52674 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 53294 270014
rect 52674 234334 53294 269778
rect 56394 274054 57014 309498
rect 60114 421774 60734 457218
rect 64208 435454 64528 435486
rect 64208 435218 64250 435454
rect 64486 435218 64528 435454
rect 64208 435134 64528 435218
rect 64208 434898 64250 435134
rect 64486 434898 64528 435134
rect 64208 434866 64528 434898
rect 73794 435454 74414 470898
rect 73794 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 74414 435454
rect 73794 435134 74414 435218
rect 73794 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 74414 435134
rect 60114 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 60734 421774
rect 60114 421454 60734 421538
rect 60114 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 60734 421454
rect 60114 385774 60734 421218
rect 64208 399454 64528 399486
rect 64208 399218 64250 399454
rect 64486 399218 64528 399454
rect 64208 399134 64528 399218
rect 64208 398898 64250 399134
rect 64486 398898 64528 399134
rect 64208 398866 64528 398898
rect 73794 399454 74414 434898
rect 73794 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 74414 399454
rect 73794 399134 74414 399218
rect 73794 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 74414 399134
rect 60114 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 60734 385774
rect 60114 385454 60734 385538
rect 60114 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 60734 385454
rect 60114 349774 60734 385218
rect 60114 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 60734 349774
rect 60114 349454 60734 349538
rect 60114 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 60734 349454
rect 60114 313774 60734 349218
rect 60114 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 60734 313774
rect 60114 313454 60734 313538
rect 60114 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 60734 313454
rect 60114 300449 60734 313218
rect 63834 389494 64454 389988
rect 63834 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 64454 389494
rect 63834 389174 64454 389258
rect 63834 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 64454 389174
rect 63834 353494 64454 388938
rect 63834 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 64454 353494
rect 63834 353174 64454 353258
rect 63834 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 64454 353174
rect 63834 317494 64454 352938
rect 63834 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 64454 317494
rect 63834 317174 64454 317258
rect 63834 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 64454 317174
rect 63834 300449 64454 316938
rect 73794 363454 74414 398898
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 300449 74414 326898
rect 77514 547174 78134 558575
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 81234 550894 81854 558575
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 79568 511174 79888 511206
rect 79568 510938 79610 511174
rect 79846 510938 79888 511174
rect 79568 510854 79888 510938
rect 79568 510618 79610 510854
rect 79846 510618 79888 510854
rect 79568 510586 79888 510618
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 439174 78134 474618
rect 79568 475174 79888 475206
rect 79568 474938 79610 475174
rect 79846 474938 79888 475174
rect 79568 474854 79888 474938
rect 79568 474618 79610 474854
rect 79846 474618 79888 474854
rect 79568 474586 79888 474618
rect 81234 442894 81854 478338
rect 81234 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 81854 442894
rect 81234 442574 81854 442658
rect 81234 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 81854 442574
rect 77514 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 78134 439174
rect 77514 438854 78134 438938
rect 77514 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 78134 438854
rect 77514 403174 78134 438618
rect 79568 439174 79888 439206
rect 79568 438938 79610 439174
rect 79846 438938 79888 439174
rect 79568 438854 79888 438938
rect 79568 438618 79610 438854
rect 79846 438618 79888 438854
rect 79568 438586 79888 438618
rect 81234 406894 81854 442338
rect 81234 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 81854 406894
rect 81234 406574 81854 406658
rect 81234 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 81854 406574
rect 77514 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 78134 403174
rect 77514 402854 78134 402938
rect 77514 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 78134 402854
rect 77514 367174 78134 402618
rect 79568 403174 79888 403206
rect 79568 402938 79610 403174
rect 79846 402938 79888 403174
rect 79568 402854 79888 402938
rect 79568 402618 79610 402854
rect 79846 402618 79888 402854
rect 79568 402586 79888 402618
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 300449 78134 330618
rect 81234 370894 81854 406338
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 300449 81854 334338
rect 84954 554614 85574 558575
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446614 85574 482058
rect 84954 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 85574 446614
rect 84954 446294 85574 446378
rect 84954 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 85574 446294
rect 84954 410614 85574 446058
rect 84954 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 85574 410614
rect 84954 410294 85574 410378
rect 84954 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 85574 410294
rect 84954 374614 85574 410058
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 300449 85574 302058
rect 88674 558334 89294 558575
rect 88674 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 89294 558334
rect 88674 558014 89294 558098
rect 88674 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 89294 558014
rect 88674 522334 89294 557778
rect 88674 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 89294 522334
rect 88674 522014 89294 522098
rect 88674 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 89294 522014
rect 88674 486334 89294 521778
rect 88674 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 89294 486334
rect 88674 486014 89294 486098
rect 88674 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 89294 486014
rect 88674 450334 89294 485778
rect 88674 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 89294 450334
rect 88674 450014 89294 450098
rect 88674 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 89294 450014
rect 88674 414334 89294 449778
rect 88674 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 89294 414334
rect 88674 414014 89294 414098
rect 88674 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 89294 414014
rect 88674 378334 89294 413778
rect 88674 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 89294 378334
rect 88674 378014 89294 378098
rect 88674 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 89294 378014
rect 88674 342334 89294 377778
rect 88674 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 89294 342334
rect 88674 342014 89294 342098
rect 88674 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 89294 342014
rect 88674 306334 89294 341778
rect 88674 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 89294 306334
rect 88674 306014 89294 306098
rect 88674 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 89294 306014
rect 88674 300449 89294 305778
rect 92394 526054 93014 558575
rect 92394 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 93014 526054
rect 92394 525734 93014 525818
rect 92394 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 93014 525734
rect 92394 490054 93014 525498
rect 96114 529774 96734 558575
rect 96114 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 96734 529774
rect 96114 529454 96734 529538
rect 96114 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 96734 529454
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 92394 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 93014 490054
rect 92394 489734 93014 489818
rect 92394 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 93014 489734
rect 92394 454054 93014 489498
rect 96114 493774 96734 529218
rect 96114 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 96734 493774
rect 96114 493454 96734 493538
rect 96114 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 96734 493454
rect 94928 471454 95248 471486
rect 94928 471218 94970 471454
rect 95206 471218 95248 471454
rect 94928 471134 95248 471218
rect 94928 470898 94970 471134
rect 95206 470898 95248 471134
rect 94928 470866 95248 470898
rect 92394 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 93014 454054
rect 92394 453734 93014 453818
rect 92394 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 93014 453734
rect 92394 418054 93014 453498
rect 96114 457774 96734 493218
rect 96114 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 96734 457774
rect 96114 457454 96734 457538
rect 96114 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 96734 457454
rect 94928 435454 95248 435486
rect 94928 435218 94970 435454
rect 95206 435218 95248 435454
rect 94928 435134 95248 435218
rect 94928 434898 94970 435134
rect 95206 434898 95248 435134
rect 94928 434866 95248 434898
rect 92394 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 93014 418054
rect 92394 417734 93014 417818
rect 92394 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 93014 417734
rect 92394 382054 93014 417498
rect 96114 421774 96734 457218
rect 96114 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 96734 421774
rect 96114 421454 96734 421538
rect 96114 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 96734 421454
rect 94928 399454 95248 399486
rect 94928 399218 94970 399454
rect 95206 399218 95248 399454
rect 94928 399134 95248 399218
rect 94928 398898 94970 399134
rect 95206 398898 95248 399134
rect 94928 398866 95248 398898
rect 92394 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 93014 382054
rect 92394 381734 93014 381818
rect 92394 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 93014 381734
rect 92394 346054 93014 381498
rect 92394 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 93014 346054
rect 92394 345734 93014 345818
rect 92394 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 93014 345734
rect 92394 310054 93014 345498
rect 92394 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 93014 310054
rect 92394 309734 93014 309818
rect 92394 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 93014 309734
rect 92394 300449 93014 309498
rect 96114 385774 96734 421218
rect 96114 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 96734 385774
rect 96114 385454 96734 385538
rect 96114 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 96734 385454
rect 96114 349774 96734 385218
rect 96114 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 96734 349774
rect 96114 349454 96734 349538
rect 96114 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 96734 349454
rect 96114 313774 96734 349218
rect 96114 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 96734 313774
rect 96114 313454 96734 313538
rect 96114 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 96734 313454
rect 96114 300449 96734 313218
rect 99834 533494 100454 558575
rect 99834 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 100454 533494
rect 99834 533174 100454 533258
rect 99834 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 100454 533174
rect 99834 497494 100454 532938
rect 113514 547174 114134 558575
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 110288 511174 110608 511206
rect 110288 510938 110330 511174
rect 110566 510938 110608 511174
rect 110288 510854 110608 510938
rect 110288 510618 110330 510854
rect 110566 510618 110608 510854
rect 110288 510586 110608 510618
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 99834 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 100454 497494
rect 99834 497174 100454 497258
rect 99834 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 100454 497174
rect 99834 461494 100454 496938
rect 110288 475174 110608 475206
rect 110288 474938 110330 475174
rect 110566 474938 110608 475174
rect 110288 474854 110608 474938
rect 110288 474618 110330 474854
rect 110566 474618 110608 474854
rect 110288 474586 110608 474618
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 99834 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 100454 461494
rect 99834 461174 100454 461258
rect 99834 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 100454 461174
rect 99834 425494 100454 460938
rect 110288 439174 110608 439206
rect 110288 438938 110330 439174
rect 110566 438938 110608 439174
rect 110288 438854 110608 438938
rect 110288 438618 110330 438854
rect 110566 438618 110608 438854
rect 110288 438586 110608 438618
rect 113514 439174 114134 474618
rect 113514 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 114134 439174
rect 113514 438854 114134 438938
rect 113514 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 114134 438854
rect 99834 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 100454 425494
rect 99834 425174 100454 425258
rect 99834 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 100454 425174
rect 99834 389494 100454 424938
rect 110288 403174 110608 403206
rect 110288 402938 110330 403174
rect 110566 402938 110608 403174
rect 110288 402854 110608 402938
rect 110288 402618 110330 402854
rect 110566 402618 110608 402854
rect 110288 402586 110608 402618
rect 113514 403174 114134 438618
rect 113514 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 114134 403174
rect 113514 402854 114134 402938
rect 113514 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 114134 402854
rect 99834 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 100454 389494
rect 99834 389174 100454 389258
rect 99834 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 100454 389174
rect 99834 353494 100454 388938
rect 99834 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 100454 353494
rect 99834 353174 100454 353258
rect 99834 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 100454 353174
rect 99834 317494 100454 352938
rect 99834 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 100454 317494
rect 99834 317174 100454 317258
rect 99834 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 100454 317174
rect 99834 300449 100454 316938
rect 109794 363454 110414 389988
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 300449 110414 326898
rect 113514 367174 114134 402618
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 69568 295174 69888 295206
rect 69568 294938 69610 295174
rect 69846 294938 69888 295174
rect 69568 294854 69888 294938
rect 69568 294618 69610 294854
rect 69846 294618 69888 294854
rect 69568 294586 69888 294618
rect 100288 295174 100608 295206
rect 100288 294938 100330 295174
rect 100566 294938 100608 295174
rect 100288 294854 100608 294938
rect 100288 294618 100330 294854
rect 100566 294618 100608 294854
rect 100288 294586 100608 294618
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 84928 291454 85248 291486
rect 84928 291218 84970 291454
rect 85206 291218 85248 291454
rect 84928 291134 85248 291218
rect 84928 290898 84970 291134
rect 85206 290898 85248 291134
rect 84928 290866 85248 290898
rect 56394 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 57014 274054
rect 56394 273734 57014 273818
rect 56394 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 57014 273734
rect 54208 255454 54528 255486
rect 54208 255218 54250 255454
rect 54486 255218 54528 255454
rect 54208 255134 54528 255218
rect 54208 254898 54250 255134
rect 54486 254898 54528 255134
rect 54208 254866 54528 254898
rect 52674 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 53294 234334
rect 52674 234014 53294 234098
rect 52674 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 53294 234014
rect 52674 198334 53294 233778
rect 52674 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 53294 198334
rect 52674 198014 53294 198098
rect 52674 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 53294 198014
rect 52674 162334 53294 197778
rect 52674 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 53294 162334
rect 52674 162014 53294 162098
rect 52674 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 53294 162014
rect 52674 126334 53294 161778
rect 56394 238054 57014 273498
rect 69568 259174 69888 259206
rect 69568 258938 69610 259174
rect 69846 258938 69888 259174
rect 69568 258854 69888 258938
rect 69568 258618 69610 258854
rect 69846 258618 69888 258854
rect 69568 258586 69888 258618
rect 100288 259174 100608 259206
rect 100288 258938 100330 259174
rect 100566 258938 100608 259174
rect 100288 258854 100608 258938
rect 100288 258618 100330 258854
rect 100566 258618 100608 258854
rect 100288 258586 100608 258618
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 84928 255454 85248 255486
rect 84928 255218 84970 255454
rect 85206 255218 85248 255454
rect 84928 255134 85248 255218
rect 84928 254898 84970 255134
rect 85206 254898 85248 255134
rect 84928 254866 85248 254898
rect 56394 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 57014 238054
rect 56394 237734 57014 237818
rect 56394 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 57014 237734
rect 56394 202054 57014 237498
rect 59123 235924 59189 235925
rect 59123 235860 59124 235924
rect 59188 235860 59189 235924
rect 59123 235859 59189 235860
rect 58571 233748 58637 233749
rect 58571 233684 58572 233748
rect 58636 233684 58637 233748
rect 58571 233683 58637 233684
rect 56394 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 57014 202054
rect 56394 201734 57014 201818
rect 56394 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 57014 201734
rect 56394 166054 57014 201498
rect 57467 189684 57533 189685
rect 57467 189620 57468 189684
rect 57532 189620 57533 189684
rect 57467 189619 57533 189620
rect 57470 174181 57530 189619
rect 57651 186964 57717 186965
rect 57651 186900 57652 186964
rect 57716 186900 57717 186964
rect 57651 186899 57717 186900
rect 57654 179893 57714 186899
rect 57651 179892 57717 179893
rect 57651 179828 57652 179892
rect 57716 179828 57717 179892
rect 57651 179827 57717 179828
rect 57835 179484 57901 179485
rect 57835 179420 57836 179484
rect 57900 179420 57901 179484
rect 57835 179419 57901 179420
rect 57651 176492 57717 176493
rect 57651 176428 57652 176492
rect 57716 176428 57717 176492
rect 57651 176427 57717 176428
rect 57467 174180 57533 174181
rect 57467 174116 57468 174180
rect 57532 174116 57533 174180
rect 57467 174115 57533 174116
rect 57283 172412 57349 172413
rect 57283 172348 57284 172412
rect 57348 172348 57349 172412
rect 57283 172347 57349 172348
rect 56394 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 57014 166054
rect 56394 165734 57014 165818
rect 56394 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 57014 165734
rect 54339 149836 54405 149837
rect 54339 149772 54340 149836
rect 54404 149772 54405 149836
rect 54339 149771 54405 149772
rect 52674 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 53294 126334
rect 52674 126014 53294 126098
rect 52674 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 53294 126014
rect 52674 90334 53294 125778
rect 54342 116109 54402 149771
rect 56394 130054 57014 165498
rect 57286 153237 57346 172347
rect 57654 172277 57714 176427
rect 57838 176085 57898 179419
rect 57835 176084 57901 176085
rect 57835 176020 57836 176084
rect 57900 176020 57901 176084
rect 57835 176019 57901 176020
rect 57835 175268 57901 175269
rect 57835 175204 57836 175268
rect 57900 175204 57901 175268
rect 57835 175203 57901 175204
rect 57651 172276 57717 172277
rect 57651 172212 57652 172276
rect 57716 172212 57717 172276
rect 57651 172211 57717 172212
rect 57838 170373 57898 175203
rect 58574 171150 58634 233683
rect 58939 226948 59005 226949
rect 58939 226884 58940 226948
rect 59004 226884 59005 226948
rect 58939 226883 59005 226884
rect 58755 207636 58821 207637
rect 58755 207572 58756 207636
rect 58820 207572 58821 207636
rect 58755 207571 58821 207572
rect 58022 171090 58634 171150
rect 57835 170372 57901 170373
rect 57835 170308 57836 170372
rect 57900 170308 57901 170372
rect 57835 170307 57901 170308
rect 58022 167650 58082 171090
rect 57654 167590 58082 167650
rect 57654 158949 57714 167590
rect 58571 167108 58637 167109
rect 58571 167044 58572 167108
rect 58636 167044 58637 167108
rect 58571 167043 58637 167044
rect 57651 158948 57717 158949
rect 57651 158884 57652 158948
rect 57716 158884 57717 158948
rect 57651 158883 57717 158884
rect 57835 158812 57901 158813
rect 57835 158748 57836 158812
rect 57900 158748 57901 158812
rect 57835 158747 57901 158748
rect 57467 154460 57533 154461
rect 57467 154396 57468 154460
rect 57532 154396 57533 154460
rect 57467 154395 57533 154396
rect 57283 153236 57349 153237
rect 57283 153172 57284 153236
rect 57348 153172 57349 153236
rect 57283 153171 57349 153172
rect 57470 139909 57530 154395
rect 57651 144804 57717 144805
rect 57651 144740 57652 144804
rect 57716 144740 57717 144804
rect 57651 144739 57717 144740
rect 57654 141813 57714 144739
rect 57838 143717 57898 158747
rect 58574 157045 58634 167043
rect 58758 160853 58818 207571
rect 58755 160852 58821 160853
rect 58755 160788 58756 160852
rect 58820 160788 58821 160852
rect 58755 160787 58821 160788
rect 58755 160172 58821 160173
rect 58755 160108 58756 160172
rect 58820 160108 58821 160172
rect 58755 160107 58821 160108
rect 58571 157044 58637 157045
rect 58571 156980 58572 157044
rect 58636 156980 58637 157044
rect 58571 156979 58637 156980
rect 58387 156636 58453 156637
rect 58387 156572 58388 156636
rect 58452 156572 58453 156636
rect 58387 156571 58453 156572
rect 58390 145621 58450 156571
rect 58571 155956 58637 155957
rect 58571 155892 58572 155956
rect 58636 155892 58637 155956
rect 58571 155891 58637 155892
rect 58574 147525 58634 155891
rect 58758 151333 58818 160107
rect 58942 155141 59002 226883
rect 59126 171150 59186 235859
rect 60411 235244 60477 235245
rect 60411 235180 60412 235244
rect 60476 235180 60477 235244
rect 60411 235179 60477 235180
rect 60043 231164 60109 231165
rect 60043 231100 60044 231164
rect 60108 231100 60109 231164
rect 60043 231099 60109 231100
rect 59675 182068 59741 182069
rect 59675 182004 59676 182068
rect 59740 182004 59741 182068
rect 59675 182003 59741 182004
rect 59126 171090 59370 171150
rect 59310 162757 59370 171090
rect 59123 162756 59189 162757
rect 59123 162692 59124 162756
rect 59188 162692 59189 162756
rect 59123 162691 59189 162692
rect 59307 162756 59373 162757
rect 59307 162692 59308 162756
rect 59372 162692 59373 162756
rect 59307 162691 59373 162692
rect 58939 155140 59005 155141
rect 58939 155076 58940 155140
rect 59004 155076 59005 155140
rect 58939 155075 59005 155076
rect 58755 151332 58821 151333
rect 58755 151268 58756 151332
rect 58820 151268 58821 151332
rect 58755 151267 58821 151268
rect 59126 149429 59186 162691
rect 59123 149428 59189 149429
rect 59123 149364 59124 149428
rect 59188 149364 59189 149428
rect 59123 149363 59189 149364
rect 58571 147524 58637 147525
rect 58571 147460 58572 147524
rect 58636 147460 58637 147524
rect 58571 147459 58637 147460
rect 58387 145620 58453 145621
rect 58387 145556 58388 145620
rect 58452 145556 58453 145620
rect 58387 145555 58453 145556
rect 57835 143716 57901 143717
rect 57835 143652 57836 143716
rect 57900 143652 57901 143716
rect 57835 143651 57901 143652
rect 57651 141812 57717 141813
rect 57651 141748 57652 141812
rect 57716 141748 57717 141812
rect 57651 141747 57717 141748
rect 57467 139908 57533 139909
rect 57467 139844 57468 139908
rect 57532 139844 57533 139908
rect 57467 139843 57533 139844
rect 59678 136101 59738 182003
rect 59859 168740 59925 168741
rect 59859 168676 59860 168740
rect 59924 168676 59925 168740
rect 59859 168675 59925 168676
rect 59862 138549 59922 168675
rect 60046 166565 60106 231099
rect 60227 225588 60293 225589
rect 60227 225524 60228 225588
rect 60292 225524 60293 225588
rect 60227 225523 60293 225524
rect 60230 168469 60290 225523
rect 60414 181797 60474 235179
rect 73794 219454 74414 238167
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 60595 195260 60661 195261
rect 60595 195196 60596 195260
rect 60660 195196 60661 195260
rect 60595 195195 60661 195196
rect 60411 181796 60477 181797
rect 60411 181732 60412 181796
rect 60476 181732 60477 181796
rect 60411 181731 60477 181732
rect 60227 168468 60293 168469
rect 60227 168404 60228 168468
rect 60292 168404 60293 168468
rect 60227 168403 60293 168404
rect 60043 166564 60109 166565
rect 60043 166500 60044 166564
rect 60108 166500 60109 166564
rect 60043 166499 60109 166500
rect 60598 164661 60658 195195
rect 73794 183305 74414 218898
rect 77514 223174 78134 238167
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 183305 78134 186618
rect 81234 226894 81854 238167
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 183305 81854 190338
rect 84954 230614 85574 238167
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 183305 85574 194058
rect 88674 234334 89294 238167
rect 88674 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 89294 234334
rect 88674 234014 89294 234098
rect 88674 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 89294 234014
rect 88674 198334 89294 233778
rect 88674 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 89294 198334
rect 88674 198014 89294 198098
rect 88674 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 89294 198014
rect 88674 183305 89294 197778
rect 92394 238054 93014 238167
rect 92394 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 93014 238054
rect 92394 237734 93014 237818
rect 92394 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 93014 237734
rect 92394 202054 93014 237498
rect 92394 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 93014 202054
rect 92394 201734 93014 201818
rect 92394 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 93014 201734
rect 92394 183305 93014 201498
rect 113514 223174 114134 258618
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113514 183305 114134 186618
rect 117234 550894 117854 558575
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 442894 117854 478338
rect 117234 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 117854 442894
rect 117234 442574 117854 442658
rect 117234 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 117854 442574
rect 117234 406894 117854 442338
rect 117234 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 117854 406894
rect 117234 406574 117854 406658
rect 117234 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 117854 406574
rect 117234 370894 117854 406338
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 226894 117854 262338
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 60595 164660 60661 164661
rect 60595 164596 60596 164660
rect 60660 164596 60661 164660
rect 60595 164595 60661 164596
rect 117234 154894 117854 190338
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 79568 151174 79888 151206
rect 79568 150938 79610 151174
rect 79846 150938 79888 151174
rect 79568 150854 79888 150938
rect 79568 150618 79610 150854
rect 79846 150618 79888 150854
rect 79568 150586 79888 150618
rect 110288 151174 110608 151206
rect 110288 150938 110330 151174
rect 110566 150938 110608 151174
rect 110288 150854 110608 150938
rect 110288 150618 110330 150854
rect 110566 150618 110608 150854
rect 110288 150586 110608 150618
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 59859 138548 59925 138549
rect 59859 138484 59860 138548
rect 59924 138484 59925 138548
rect 59859 138483 59925 138484
rect 59675 136100 59741 136101
rect 59675 136036 59676 136100
rect 59740 136036 59741 136100
rect 59675 136035 59741 136036
rect 56394 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 57014 130054
rect 56394 129734 57014 129818
rect 56394 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 57014 129734
rect 54339 116108 54405 116109
rect 54339 116044 54340 116108
rect 54404 116044 54405 116108
rect 54339 116043 54405 116044
rect 52674 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 53294 90334
rect 52674 90014 53294 90098
rect 52674 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 53294 90014
rect 52674 54334 53294 89778
rect 56394 94054 57014 129498
rect 57835 121548 57901 121549
rect 57835 121484 57836 121548
rect 57900 121484 57901 121548
rect 57835 121483 57901 121484
rect 56394 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 57014 94054
rect 56394 93734 57014 93818
rect 56394 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 57014 93734
rect 55038 75454 55358 75486
rect 55038 75218 55080 75454
rect 55316 75218 55358 75454
rect 55038 75134 55358 75218
rect 55038 74898 55080 75134
rect 55316 74898 55358 75134
rect 55038 74866 55358 74898
rect 52674 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 53294 54334
rect 52674 54014 53294 54098
rect 52674 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 53294 54014
rect 52674 18334 53294 53778
rect 52674 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 53294 18334
rect 52674 18014 53294 18098
rect 52674 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 53294 18014
rect 52674 -4186 53294 17778
rect 52674 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 53294 -4186
rect 52674 -4506 53294 -4422
rect 52674 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 53294 -4506
rect 52674 -7654 53294 -4742
rect 56394 58054 57014 93498
rect 56394 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 57014 58054
rect 56394 57734 57014 57818
rect 56394 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 57014 57734
rect 56394 22054 57014 57498
rect 57838 51509 57898 121483
rect 60114 97774 60734 120207
rect 60114 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 60734 97774
rect 60114 97454 60734 97538
rect 60114 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 60734 97454
rect 59132 79174 59452 79206
rect 59132 78938 59174 79174
rect 59410 78938 59452 79174
rect 59132 78854 59452 78938
rect 59132 78618 59174 78854
rect 59410 78618 59452 78854
rect 59132 78586 59452 78618
rect 60114 61774 60734 97218
rect 63834 101494 64454 119988
rect 63834 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 64454 101494
rect 63834 101174 64454 101258
rect 63834 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 64454 101174
rect 63226 75454 63546 75486
rect 63226 75218 63268 75454
rect 63504 75218 63546 75454
rect 63226 75134 63546 75218
rect 63226 74898 63268 75134
rect 63504 74898 63546 75134
rect 63226 74866 63546 74898
rect 60114 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 60734 61774
rect 60114 61454 60734 61538
rect 60114 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 60734 61454
rect 57835 51508 57901 51509
rect 57835 51444 57836 51508
rect 57900 51444 57901 51508
rect 57835 51443 57901 51444
rect 57838 46205 57898 51443
rect 57835 46204 57901 46205
rect 57835 46140 57836 46204
rect 57900 46140 57901 46204
rect 57835 46139 57901 46140
rect 56394 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 57014 22054
rect 56394 21734 57014 21818
rect 56394 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 57014 21734
rect 56394 -5146 57014 21498
rect 56394 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 57014 -5146
rect 56394 -5466 57014 -5382
rect 56394 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 57014 -5466
rect 56394 -7654 57014 -5702
rect 60114 25774 60734 61218
rect 60114 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 60734 25774
rect 60114 25454 60734 25538
rect 60114 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 60734 25454
rect 60114 -6106 60734 25218
rect 60114 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 60734 -6106
rect 60114 -6426 60734 -6342
rect 60114 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 60734 -6426
rect 60114 -7654 60734 -6662
rect 63834 65494 64454 100938
rect 73794 111454 74414 120207
rect 73794 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 74414 111454
rect 73794 111134 74414 111218
rect 73794 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 74414 111134
rect 67320 79174 67640 79206
rect 67320 78938 67362 79174
rect 67598 78938 67640 79174
rect 67320 78854 67640 78938
rect 67320 78618 67362 78854
rect 67598 78618 67640 78854
rect 67320 78586 67640 78618
rect 71414 75454 71734 75486
rect 71414 75218 71456 75454
rect 71692 75218 71734 75454
rect 71414 75134 71734 75218
rect 71414 74898 71456 75134
rect 71692 74898 71734 75134
rect 71414 74866 71734 74898
rect 73794 75454 74414 110898
rect 77514 115174 78134 120207
rect 77514 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 78134 115174
rect 77514 114854 78134 114938
rect 77514 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 78134 114854
rect 75508 79174 75828 79206
rect 75508 78938 75550 79174
rect 75786 78938 75828 79174
rect 75508 78854 75828 78938
rect 75508 78618 75550 78854
rect 75786 78618 75828 78854
rect 75508 78586 75828 78618
rect 77514 79174 78134 114618
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 63834 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 64454 65494
rect 63834 65174 64454 65258
rect 63834 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 64454 65174
rect 63834 29494 64454 64938
rect 63834 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 64454 29494
rect 63834 29174 64454 29258
rect 63834 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 64454 29174
rect 63834 -7066 64454 28938
rect 63834 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 64454 -7066
rect 63834 -7386 64454 -7302
rect 63834 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 64454 -7386
rect 63834 -7654 64454 -7622
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -7654 74414 -902
rect 77514 43174 78134 78618
rect 81234 118894 81854 120207
rect 81234 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 81854 118894
rect 81234 118574 81854 118658
rect 81234 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 81854 118574
rect 81234 82894 81854 118338
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 79602 75454 79922 75486
rect 79602 75218 79644 75454
rect 79880 75218 79922 75454
rect 79602 75134 79922 75218
rect 79602 74898 79644 75134
rect 79880 74898 79922 75134
rect 79602 74866 79922 74898
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -1306 78134 6618
rect 77514 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 78134 -1306
rect 77514 -1626 78134 -1542
rect 77514 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 78134 -1626
rect 77514 -7654 78134 -1862
rect 81234 46894 81854 82338
rect 84954 86614 85574 120207
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 83696 79174 84016 79206
rect 83696 78938 83738 79174
rect 83974 78938 84016 79174
rect 83696 78854 84016 78938
rect 83696 78618 83738 78854
rect 83974 78618 84016 78854
rect 83696 78586 84016 78618
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -2266 81854 10338
rect 81234 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 81854 -2266
rect 81234 -2586 81854 -2502
rect 81234 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 81854 -2586
rect 81234 -7654 81854 -2822
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 84954 -3226 85574 14058
rect 84954 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 85574 -3226
rect 84954 -3546 85574 -3462
rect 84954 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 85574 -3546
rect 84954 -7654 85574 -3782
rect 88674 90334 89294 120207
rect 88674 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 89294 90334
rect 88674 90014 89294 90098
rect 88674 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 89294 90014
rect 88674 54334 89294 89778
rect 88674 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 89294 54334
rect 88674 54014 89294 54098
rect 88674 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 89294 54014
rect 88674 18334 89294 53778
rect 88674 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 89294 18334
rect 88674 18014 89294 18098
rect 88674 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 89294 18014
rect 88674 -4186 89294 17778
rect 88674 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 89294 -4186
rect 88674 -4506 89294 -4422
rect 88674 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 89294 -4506
rect 88674 -7654 89294 -4742
rect 92394 94054 93014 120207
rect 92394 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 93014 94054
rect 92394 93734 93014 93818
rect 92394 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 93014 93734
rect 92394 58054 93014 93498
rect 92394 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 93014 58054
rect 92394 57734 93014 57818
rect 92394 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 93014 57734
rect 92394 22054 93014 57498
rect 92394 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 93014 22054
rect 92394 21734 93014 21818
rect 92394 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 93014 21734
rect 92394 -5146 93014 21498
rect 92394 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 93014 -5146
rect 92394 -5466 93014 -5382
rect 92394 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 93014 -5466
rect 92394 -7654 93014 -5702
rect 96114 97774 96734 120207
rect 96114 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 96734 97774
rect 96114 97454 96734 97538
rect 96114 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 96734 97454
rect 96114 61774 96734 97218
rect 96114 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 96734 61774
rect 96114 61454 96734 61538
rect 96114 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 96734 61454
rect 96114 25774 96734 61218
rect 96114 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 96734 25774
rect 96114 25454 96734 25538
rect 96114 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 96734 25454
rect 96114 -6106 96734 25218
rect 96114 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 96734 -6106
rect 96114 -6426 96734 -6342
rect 96114 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 96734 -6426
rect 96114 -7654 96734 -6662
rect 99834 101494 100454 120207
rect 99834 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 100454 101494
rect 99834 101174 100454 101258
rect 99834 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 100454 101174
rect 99834 65494 100454 100938
rect 99834 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 100454 65494
rect 99834 65174 100454 65258
rect 99834 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 100454 65174
rect 99834 29494 100454 64938
rect 99834 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 100454 29494
rect 99834 29174 100454 29258
rect 99834 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 100454 29174
rect 99834 -7066 100454 28938
rect 99834 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 100454 -7066
rect 99834 -7386 100454 -7302
rect 99834 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 100454 -7386
rect 99834 -7654 100454 -7622
rect 109794 111454 110414 119988
rect 109794 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 110414 111454
rect 109794 111134 110414 111218
rect 109794 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 110414 111134
rect 109794 75454 110414 110898
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -7654 110414 -902
rect 113514 115174 114134 120207
rect 113514 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 114134 115174
rect 113514 114854 114134 114938
rect 113514 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 114134 114854
rect 113514 79174 114134 114618
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -1306 114134 6618
rect 113514 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 114134 -1306
rect 113514 -1626 114134 -1542
rect 113514 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 114134 -1626
rect 113514 -7654 114134 -1862
rect 117234 118894 117854 154338
rect 117234 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 117854 118894
rect 117234 118574 117854 118658
rect 117234 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 117854 118574
rect 117234 82894 117854 118338
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -2266 117854 10338
rect 117234 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 117854 -2266
rect 117234 -2586 117854 -2502
rect 117234 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 117854 -2586
rect 117234 -7654 117854 -2822
rect 120954 554614 121574 558575
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 446614 121574 482058
rect 120954 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 121574 446614
rect 120954 446294 121574 446378
rect 120954 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 121574 446294
rect 120954 410614 121574 446058
rect 120954 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 121574 410614
rect 120954 410294 121574 410378
rect 120954 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 121574 410294
rect 120954 374614 121574 410058
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120954 158614 121574 194058
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 122614 121574 158058
rect 120954 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 121574 122614
rect 120954 122294 121574 122378
rect 120954 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 121574 122294
rect 120954 86614 121574 122058
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 120954 -3226 121574 14058
rect 120954 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 121574 -3226
rect 120954 -3546 121574 -3462
rect 120954 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 121574 -3546
rect 120954 -7654 121574 -3782
rect 124674 558334 125294 558575
rect 124674 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 125294 558334
rect 124674 558014 125294 558098
rect 124674 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 125294 558014
rect 124674 522334 125294 557778
rect 124674 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 125294 522334
rect 124674 522014 125294 522098
rect 124674 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 125294 522014
rect 124674 486334 125294 521778
rect 128394 526054 129014 558575
rect 128394 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 129014 526054
rect 128394 525734 129014 525818
rect 128394 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 129014 525734
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 124674 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 125294 486334
rect 124674 486014 125294 486098
rect 124674 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 125294 486014
rect 124674 450334 125294 485778
rect 128394 490054 129014 525498
rect 128394 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 129014 490054
rect 128394 489734 129014 489818
rect 128394 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 129014 489734
rect 125648 471454 125968 471486
rect 125648 471218 125690 471454
rect 125926 471218 125968 471454
rect 125648 471134 125968 471218
rect 125648 470898 125690 471134
rect 125926 470898 125968 471134
rect 125648 470866 125968 470898
rect 124674 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 125294 450334
rect 124674 450014 125294 450098
rect 124674 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 125294 450014
rect 124674 414334 125294 449778
rect 128394 454054 129014 489498
rect 128394 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 129014 454054
rect 128394 453734 129014 453818
rect 128394 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 129014 453734
rect 125648 435454 125968 435486
rect 125648 435218 125690 435454
rect 125926 435218 125968 435454
rect 125648 435134 125968 435218
rect 125648 434898 125690 435134
rect 125926 434898 125968 435134
rect 125648 434866 125968 434898
rect 124674 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 125294 414334
rect 124674 414014 125294 414098
rect 124674 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 125294 414014
rect 124674 378334 125294 413778
rect 128394 418054 129014 453498
rect 128394 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 129014 418054
rect 128394 417734 129014 417818
rect 128394 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 129014 417734
rect 125648 399454 125968 399486
rect 125648 399218 125690 399454
rect 125926 399218 125968 399454
rect 125648 399134 125968 399218
rect 125648 398898 125690 399134
rect 125926 398898 125968 399134
rect 125648 398866 125968 398898
rect 124674 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 125294 378334
rect 124674 378014 125294 378098
rect 124674 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 125294 378014
rect 124674 342334 125294 377778
rect 124674 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 125294 342334
rect 124674 342014 125294 342098
rect 124674 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 125294 342014
rect 124674 306334 125294 341778
rect 124674 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 125294 306334
rect 124674 306014 125294 306098
rect 124674 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 125294 306014
rect 124674 270334 125294 305778
rect 124674 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 125294 270334
rect 124674 270014 125294 270098
rect 124674 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 125294 270014
rect 124674 234334 125294 269778
rect 124674 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 125294 234334
rect 124674 234014 125294 234098
rect 124674 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 125294 234014
rect 124674 198334 125294 233778
rect 124674 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 125294 198334
rect 124674 198014 125294 198098
rect 124674 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 125294 198014
rect 124674 162334 125294 197778
rect 124674 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 125294 162334
rect 124674 162014 125294 162098
rect 124674 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 125294 162014
rect 124674 126334 125294 161778
rect 128394 382054 129014 417498
rect 128394 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 129014 382054
rect 128394 381734 129014 381818
rect 128394 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 129014 381734
rect 128394 346054 129014 381498
rect 128394 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 129014 346054
rect 128394 345734 129014 345818
rect 128394 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 129014 345734
rect 128394 310054 129014 345498
rect 128394 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 129014 310054
rect 128394 309734 129014 309818
rect 128394 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 129014 309734
rect 128394 274054 129014 309498
rect 128394 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 129014 274054
rect 128394 273734 129014 273818
rect 128394 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 129014 273734
rect 128394 238054 129014 273498
rect 128394 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 129014 238054
rect 128394 237734 129014 237818
rect 128394 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 129014 237734
rect 128394 202054 129014 237498
rect 128394 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 129014 202054
rect 128394 201734 129014 201818
rect 128394 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 129014 201734
rect 128394 166054 129014 201498
rect 128394 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 129014 166054
rect 128394 165734 129014 165818
rect 128394 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 129014 165734
rect 127571 148340 127637 148341
rect 127571 148276 127572 148340
rect 127636 148276 127637 148340
rect 127571 148275 127637 148276
rect 124674 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 125294 126334
rect 124674 126014 125294 126098
rect 124674 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 125294 126014
rect 124674 90334 125294 125778
rect 127574 121413 127634 148275
rect 127755 146708 127821 146709
rect 127755 146644 127756 146708
rect 127820 146644 127821 146708
rect 127755 146643 127821 146644
rect 127571 121412 127637 121413
rect 127571 121348 127572 121412
rect 127636 121348 127637 121412
rect 127571 121347 127637 121348
rect 127758 119917 127818 146643
rect 127939 145076 128005 145077
rect 127939 145012 127940 145076
rect 128004 145012 128005 145076
rect 127939 145011 128005 145012
rect 127755 119916 127821 119917
rect 127755 119852 127756 119916
rect 127820 119852 127821 119916
rect 127755 119851 127821 119852
rect 127942 119781 128002 145011
rect 128123 143444 128189 143445
rect 128123 143380 128124 143444
rect 128188 143380 128189 143444
rect 128123 143379 128189 143380
rect 128126 121277 128186 143379
rect 128394 130054 129014 165498
rect 128394 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 129014 130054
rect 128394 129734 129014 129818
rect 128394 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 129014 129734
rect 128123 121276 128189 121277
rect 128123 121212 128124 121276
rect 128188 121212 128189 121276
rect 128123 121211 128189 121212
rect 127939 119780 128005 119781
rect 127939 119716 127940 119780
rect 128004 119716 128005 119780
rect 127939 119715 128005 119716
rect 124674 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 125294 90334
rect 124674 90014 125294 90098
rect 124674 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 125294 90014
rect 124674 54334 125294 89778
rect 124674 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 125294 54334
rect 124674 54014 125294 54098
rect 124674 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 125294 54014
rect 124674 18334 125294 53778
rect 124674 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 125294 18334
rect 124674 18014 125294 18098
rect 124674 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 125294 18014
rect 124674 -4186 125294 17778
rect 124674 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 125294 -4186
rect 124674 -4506 125294 -4422
rect 124674 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 125294 -4506
rect 124674 -7654 125294 -4742
rect 128394 94054 129014 129498
rect 128394 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 129014 94054
rect 128394 93734 129014 93818
rect 128394 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 129014 93734
rect 128394 58054 129014 93498
rect 128394 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 129014 58054
rect 128394 57734 129014 57818
rect 128394 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 129014 57734
rect 128394 22054 129014 57498
rect 128394 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 129014 22054
rect 128394 21734 129014 21818
rect 128394 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 129014 21734
rect 128394 -5146 129014 21498
rect 128394 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 129014 -5146
rect 128394 -5466 129014 -5382
rect 128394 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 129014 -5466
rect 128394 -7654 129014 -5702
rect 132114 529774 132734 558575
rect 132114 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 132734 529774
rect 132114 529454 132734 529538
rect 132114 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 132734 529454
rect 132114 493774 132734 529218
rect 132114 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 132734 493774
rect 132114 493454 132734 493538
rect 132114 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 132734 493454
rect 132114 457774 132734 493218
rect 132114 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 132734 457774
rect 132114 457454 132734 457538
rect 132114 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 132734 457454
rect 132114 421774 132734 457218
rect 132114 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 132734 421774
rect 132114 421454 132734 421538
rect 132114 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 132734 421454
rect 132114 385774 132734 421218
rect 132114 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 132734 385774
rect 132114 385454 132734 385538
rect 132114 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 132734 385454
rect 132114 349774 132734 385218
rect 132114 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 132734 349774
rect 132114 349454 132734 349538
rect 132114 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 132734 349454
rect 132114 313774 132734 349218
rect 132114 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 132734 313774
rect 132114 313454 132734 313538
rect 132114 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 132734 313454
rect 132114 277774 132734 313218
rect 132114 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 132734 277774
rect 132114 277454 132734 277538
rect 132114 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 132734 277454
rect 132114 241774 132734 277218
rect 132114 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 132734 241774
rect 132114 241454 132734 241538
rect 132114 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 132734 241454
rect 132114 205774 132734 241218
rect 132114 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 132734 205774
rect 132114 205454 132734 205538
rect 132114 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 132734 205454
rect 132114 169774 132734 205218
rect 135834 533494 136454 568938
rect 135834 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 136454 533494
rect 135834 533174 136454 533258
rect 135834 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 136454 533174
rect 135834 497494 136454 532938
rect 145794 704838 146414 711590
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 141008 511174 141328 511206
rect 141008 510938 141050 511174
rect 141286 510938 141328 511174
rect 141008 510854 141328 510938
rect 141008 510618 141050 510854
rect 141286 510618 141328 510854
rect 141008 510586 141328 510618
rect 135834 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 136454 497494
rect 135834 497174 136454 497258
rect 135834 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 136454 497174
rect 135834 461494 136454 496938
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 141008 475174 141328 475206
rect 141008 474938 141050 475174
rect 141286 474938 141328 475174
rect 141008 474854 141328 474938
rect 141008 474618 141050 474854
rect 141286 474618 141328 474854
rect 141008 474586 141328 474618
rect 135834 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 136454 461494
rect 135834 461174 136454 461258
rect 135834 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 136454 461174
rect 135834 425494 136454 460938
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 141008 439174 141328 439206
rect 141008 438938 141050 439174
rect 141286 438938 141328 439174
rect 141008 438854 141328 438938
rect 141008 438618 141050 438854
rect 141286 438618 141328 438854
rect 141008 438586 141328 438618
rect 135834 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 136454 425494
rect 135834 425174 136454 425258
rect 135834 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 136454 425174
rect 135834 389494 136454 424938
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 141008 403174 141328 403206
rect 141008 402938 141050 403174
rect 141286 402938 141328 403174
rect 141008 402854 141328 402938
rect 141008 402618 141050 402854
rect 141286 402618 141328 402854
rect 141008 402586 141328 402618
rect 135834 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 136454 389494
rect 135834 389174 136454 389258
rect 135834 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 136454 389174
rect 135834 353494 136454 388938
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 137139 382940 137205 382941
rect 137139 382876 137140 382940
rect 137204 382876 137205 382940
rect 137139 382875 137205 382876
rect 135834 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 136454 353494
rect 135834 353174 136454 353258
rect 135834 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 136454 353174
rect 135834 317494 136454 352938
rect 135834 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 136454 317494
rect 135834 317174 136454 317258
rect 135834 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 136454 317174
rect 135834 281494 136454 316938
rect 135834 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 136454 281494
rect 135834 281174 136454 281258
rect 135834 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 136454 281174
rect 135834 245494 136454 280938
rect 135834 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 136454 245494
rect 135834 245174 136454 245258
rect 135834 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 136454 245174
rect 135834 209494 136454 244938
rect 135834 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 136454 209494
rect 135834 209174 136454 209258
rect 135834 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 136454 209174
rect 134379 184516 134445 184517
rect 134379 184452 134380 184516
rect 134444 184452 134445 184516
rect 134379 184451 134445 184452
rect 132114 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 132734 169774
rect 134382 169557 134442 184451
rect 135834 173494 136454 208938
rect 135834 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 136454 173494
rect 135834 173174 136454 173258
rect 135834 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 136454 173174
rect 132114 169454 132734 169538
rect 134379 169556 134445 169557
rect 134379 169492 134380 169556
rect 134444 169492 134445 169556
rect 134379 169491 134445 169492
rect 132114 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 132734 169454
rect 132114 133774 132734 169218
rect 132114 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 132734 133774
rect 132114 133454 132734 133538
rect 132114 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 132734 133454
rect 132114 97774 132734 133218
rect 132114 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 132734 97774
rect 132114 97454 132734 97538
rect 132114 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 132734 97454
rect 132114 61774 132734 97218
rect 132114 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 132734 61774
rect 132114 61454 132734 61538
rect 132114 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 132734 61454
rect 132114 25774 132734 61218
rect 132114 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 132734 25774
rect 132114 25454 132734 25538
rect 132114 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 132734 25454
rect 132114 -6106 132734 25218
rect 132114 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 132734 -6106
rect 132114 -6426 132734 -6342
rect 132114 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 132734 -6426
rect 132114 -7654 132734 -6662
rect 135834 137494 136454 172938
rect 137142 163029 137202 382875
rect 145794 363454 146414 398898
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 219454 146414 254898
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 137139 163028 137205 163029
rect 137139 162964 137140 163028
rect 137204 162964 137205 163028
rect 137139 162963 137205 162964
rect 135834 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 136454 137494
rect 135834 137174 136454 137258
rect 135834 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 136454 137174
rect 135834 101494 136454 136938
rect 135834 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 136454 101494
rect 135834 101174 136454 101258
rect 135834 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 136454 101174
rect 135834 65494 136454 100938
rect 135834 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 136454 65494
rect 135834 65174 136454 65258
rect 135834 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 136454 65174
rect 135834 29494 136454 64938
rect 135834 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 136454 29494
rect 135834 29174 136454 29258
rect 135834 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 136454 29174
rect 135834 -7066 136454 28938
rect 135834 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 136454 -7066
rect 135834 -7386 136454 -7302
rect 135834 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 136454 -7386
rect 135834 -7654 136454 -7622
rect 145794 147454 146414 182898
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 111454 146414 146898
rect 145794 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 146414 111454
rect 145794 111134 146414 111218
rect 145794 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 146414 111134
rect 145794 75454 146414 110898
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -7654 146414 -902
rect 149514 705798 150134 711590
rect 149514 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 150134 705798
rect 149514 705478 150134 705562
rect 149514 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 150134 705478
rect 149514 691174 150134 705242
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 223174 150134 258618
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 149514 151174 150134 186618
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 115174 150134 150618
rect 149514 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 150134 115174
rect 149514 114854 150134 114938
rect 149514 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 150134 114854
rect 149514 79174 150134 114618
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -1306 150134 6618
rect 149514 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 150134 -1306
rect 149514 -1626 150134 -1542
rect 149514 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 150134 -1626
rect 149514 -7654 150134 -1862
rect 153234 706758 153854 711590
rect 153234 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 153854 706758
rect 153234 706438 153854 706522
rect 153234 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 153854 706438
rect 153234 694894 153854 706202
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 156954 707718 157574 711590
rect 156954 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 157574 707718
rect 156954 707398 157574 707482
rect 156954 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 157574 707398
rect 156954 698614 157574 707162
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156368 471454 156688 471486
rect 156368 471218 156410 471454
rect 156646 471218 156688 471454
rect 156368 471134 156688 471218
rect 156368 470898 156410 471134
rect 156646 470898 156688 471134
rect 156368 470866 156688 470898
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 156954 446614 157574 482058
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156368 435454 156688 435486
rect 156368 435218 156410 435454
rect 156646 435218 156688 435454
rect 156368 435134 156688 435218
rect 156368 434898 156410 435134
rect 156646 434898 156688 435134
rect 156368 434866 156688 434898
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156368 399454 156688 399486
rect 156368 399218 156410 399454
rect 156646 399218 156688 399454
rect 156368 399134 156688 399218
rect 156368 398898 156410 399134
rect 156646 398898 156688 399134
rect 156368 398866 156688 398898
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 226894 153854 262338
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 153234 190894 153854 226338
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 154894 153854 190338
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 118894 153854 154338
rect 153234 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 153854 118894
rect 153234 118574 153854 118658
rect 153234 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 153854 118574
rect 153234 82894 153854 118338
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -2266 153854 10338
rect 153234 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 153854 -2266
rect 153234 -2586 153854 -2502
rect 153234 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 153854 -2586
rect 153234 -7654 153854 -2822
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 158614 157574 194058
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 122614 157574 158058
rect 156954 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 157574 122614
rect 156954 122294 157574 122378
rect 156954 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 157574 122294
rect 156954 86614 157574 122058
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 156954 -3226 157574 14058
rect 156954 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 157574 -3226
rect 156954 -3546 157574 -3462
rect 156954 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 157574 -3546
rect 156954 -7654 157574 -3782
rect 160674 708678 161294 711590
rect 160674 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 161294 708678
rect 160674 708358 161294 708442
rect 160674 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 161294 708358
rect 160674 666334 161294 708122
rect 160674 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 161294 666334
rect 160674 666014 161294 666098
rect 160674 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 161294 666014
rect 160674 630334 161294 665778
rect 160674 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 161294 630334
rect 160674 630014 161294 630098
rect 160674 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 161294 630014
rect 160674 594334 161294 629778
rect 160674 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 161294 594334
rect 160674 594014 161294 594098
rect 160674 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 161294 594014
rect 160674 558334 161294 593778
rect 160674 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 161294 558334
rect 160674 558014 161294 558098
rect 160674 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 161294 558014
rect 160674 522334 161294 557778
rect 160674 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 161294 522334
rect 160674 522014 161294 522098
rect 160674 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 161294 522014
rect 160674 486334 161294 521778
rect 160674 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 161294 486334
rect 160674 486014 161294 486098
rect 160674 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 161294 486014
rect 160674 450334 161294 485778
rect 160674 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 161294 450334
rect 160674 450014 161294 450098
rect 160674 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 161294 450014
rect 160674 414334 161294 449778
rect 160674 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 161294 414334
rect 160674 414014 161294 414098
rect 160674 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 161294 414014
rect 160674 378334 161294 413778
rect 160674 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 161294 378334
rect 160674 378014 161294 378098
rect 160674 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 161294 378014
rect 160674 342334 161294 377778
rect 160674 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 161294 342334
rect 160674 342014 161294 342098
rect 160674 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 161294 342014
rect 160674 306334 161294 341778
rect 160674 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 161294 306334
rect 160674 306014 161294 306098
rect 160674 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 161294 306014
rect 160674 270334 161294 305778
rect 160674 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 161294 270334
rect 160674 270014 161294 270098
rect 160674 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 161294 270014
rect 160674 234334 161294 269778
rect 160674 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 161294 234334
rect 160674 234014 161294 234098
rect 160674 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 161294 234014
rect 160674 198334 161294 233778
rect 160674 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 161294 198334
rect 160674 198014 161294 198098
rect 160674 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 161294 198014
rect 160674 162334 161294 197778
rect 160674 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 161294 162334
rect 160674 162014 161294 162098
rect 160674 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 161294 162014
rect 160674 126334 161294 161778
rect 160674 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 161294 126334
rect 160674 126014 161294 126098
rect 160674 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 161294 126014
rect 160674 90334 161294 125778
rect 160674 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 161294 90334
rect 160674 90014 161294 90098
rect 160674 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 161294 90014
rect 160674 54334 161294 89778
rect 160674 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 161294 54334
rect 160674 54014 161294 54098
rect 160674 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 161294 54014
rect 160674 18334 161294 53778
rect 160674 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 161294 18334
rect 160674 18014 161294 18098
rect 160674 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 161294 18014
rect 160674 -4186 161294 17778
rect 160674 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 161294 -4186
rect 160674 -4506 161294 -4422
rect 160674 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 161294 -4506
rect 160674 -7654 161294 -4742
rect 164394 709638 165014 711590
rect 164394 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 165014 709638
rect 164394 709318 165014 709402
rect 164394 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 165014 709318
rect 164394 670054 165014 709082
rect 164394 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 165014 670054
rect 164394 669734 165014 669818
rect 164394 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 165014 669734
rect 164394 634054 165014 669498
rect 164394 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 165014 634054
rect 164394 633734 165014 633818
rect 164394 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 165014 633734
rect 164394 598054 165014 633498
rect 168114 710598 168734 711590
rect 168114 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 168734 710598
rect 168114 710278 168734 710362
rect 168114 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 168734 710278
rect 168114 673774 168734 710042
rect 168114 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 168734 673774
rect 168114 673454 168734 673538
rect 168114 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 168734 673454
rect 168114 637774 168734 673218
rect 168114 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 168734 637774
rect 168114 637454 168734 637538
rect 168114 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 168734 637454
rect 166763 603940 166829 603941
rect 166763 603876 166764 603940
rect 166828 603876 166829 603940
rect 166763 603875 166829 603876
rect 164394 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 165014 598054
rect 164394 597734 165014 597818
rect 164394 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 165014 597734
rect 164394 562054 165014 597498
rect 166579 571300 166645 571301
rect 166579 571236 166580 571300
rect 166644 571236 166645 571300
rect 166579 571235 166645 571236
rect 164394 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 165014 562054
rect 164394 561734 165014 561818
rect 164394 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 165014 561734
rect 164394 526054 165014 561498
rect 166582 537573 166642 571235
rect 166766 560285 166826 603875
rect 168114 601774 168734 637218
rect 168114 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 168734 601774
rect 168114 601454 168734 601538
rect 168114 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 168734 601454
rect 168114 565774 168734 601218
rect 171834 711558 172454 711590
rect 171834 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 172454 711558
rect 171834 711238 172454 711322
rect 171834 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 172454 711238
rect 171834 677494 172454 711002
rect 171834 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 172454 677494
rect 171834 677174 172454 677258
rect 171834 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 172454 677174
rect 171834 641494 172454 676938
rect 181794 704838 182414 711590
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 179275 655076 179341 655077
rect 179275 655012 179276 655076
rect 179340 655012 179341 655076
rect 179275 655011 179341 655012
rect 175043 653172 175109 653173
rect 175043 653108 175044 653172
rect 175108 653108 175109 653172
rect 175043 653107 175109 653108
rect 171834 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 172454 641494
rect 171834 641174 172454 641258
rect 171834 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 172454 641174
rect 171834 605494 172454 640938
rect 175046 619173 175106 653107
rect 176515 650044 176581 650045
rect 176515 649980 176516 650044
rect 176580 649980 176581 650044
rect 176515 649979 176581 649980
rect 176331 647324 176397 647325
rect 176331 647260 176332 647324
rect 176396 647260 176397 647324
rect 176331 647259 176397 647260
rect 176147 645964 176213 645965
rect 176147 645900 176148 645964
rect 176212 645900 176213 645964
rect 176147 645899 176213 645900
rect 176150 625701 176210 645899
rect 176147 625700 176213 625701
rect 176147 625636 176148 625700
rect 176212 625636 176213 625700
rect 176147 625635 176213 625636
rect 175043 619172 175109 619173
rect 175043 619108 175044 619172
rect 175108 619108 175109 619172
rect 175043 619107 175109 619108
rect 172651 618356 172717 618357
rect 172651 618292 172652 618356
rect 172716 618292 172717 618356
rect 172651 618291 172717 618292
rect 171834 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 172454 605494
rect 171834 605174 172454 605258
rect 171834 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 172454 605174
rect 171547 570076 171613 570077
rect 171547 570012 171548 570076
rect 171612 570012 171613 570076
rect 171547 570011 171613 570012
rect 168114 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 168734 565774
rect 168114 565454 168734 565538
rect 168114 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 168734 565454
rect 166763 560284 166829 560285
rect 166763 560220 166764 560284
rect 166828 560220 166829 560284
rect 166763 560219 166829 560220
rect 166579 537572 166645 537573
rect 166579 537508 166580 537572
rect 166644 537508 166645 537572
rect 166579 537507 166645 537508
rect 164394 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 165014 526054
rect 164394 525734 165014 525818
rect 164394 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 165014 525734
rect 164394 490054 165014 525498
rect 164394 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 165014 490054
rect 164394 489734 165014 489818
rect 164394 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 165014 489734
rect 164394 454054 165014 489498
rect 164394 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 165014 454054
rect 164394 453734 165014 453818
rect 164394 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 165014 453734
rect 164394 418054 165014 453498
rect 164394 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 165014 418054
rect 164394 417734 165014 417818
rect 164394 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 165014 417734
rect 164394 382054 165014 417498
rect 164394 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 165014 382054
rect 164394 381734 165014 381818
rect 164394 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 165014 381734
rect 164394 346054 165014 381498
rect 164394 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 165014 346054
rect 164394 345734 165014 345818
rect 164394 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 165014 345734
rect 164394 310054 165014 345498
rect 164394 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 165014 310054
rect 164394 309734 165014 309818
rect 164394 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 165014 309734
rect 164394 274054 165014 309498
rect 164394 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 165014 274054
rect 164394 273734 165014 273818
rect 164394 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 165014 273734
rect 164394 238054 165014 273498
rect 164394 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 165014 238054
rect 164394 237734 165014 237818
rect 164394 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 165014 237734
rect 164394 202054 165014 237498
rect 164394 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 165014 202054
rect 164394 201734 165014 201818
rect 164394 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 165014 201734
rect 164394 166054 165014 201498
rect 164394 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 165014 166054
rect 164394 165734 165014 165818
rect 164394 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 165014 165734
rect 164394 130054 165014 165498
rect 164394 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 165014 130054
rect 164394 129734 165014 129818
rect 164394 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 165014 129734
rect 164394 94054 165014 129498
rect 164394 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 165014 94054
rect 164394 93734 165014 93818
rect 164394 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 165014 93734
rect 164394 58054 165014 93498
rect 164394 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 165014 58054
rect 164394 57734 165014 57818
rect 164394 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 165014 57734
rect 164394 22054 165014 57498
rect 164394 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 165014 22054
rect 164394 21734 165014 21818
rect 164394 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 165014 21734
rect 164394 -5146 165014 21498
rect 164394 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 165014 -5146
rect 164394 -5466 165014 -5382
rect 164394 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 165014 -5466
rect 164394 -7654 165014 -5702
rect 168114 529774 168734 565218
rect 171550 541789 171610 570011
rect 171834 569494 172454 604938
rect 171834 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 172454 569494
rect 171834 569174 172454 569258
rect 171834 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 172454 569174
rect 171547 541788 171613 541789
rect 171547 541724 171548 541788
rect 171612 541724 171613 541788
rect 171547 541723 171613 541724
rect 168114 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 168734 529774
rect 168114 529454 168734 529538
rect 168114 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 168734 529454
rect 168114 493774 168734 529218
rect 171834 533494 172454 568938
rect 172654 561645 172714 618291
rect 175227 617540 175293 617541
rect 175227 617476 175228 617540
rect 175292 617476 175293 617540
rect 175227 617475 175293 617476
rect 173939 616724 174005 616725
rect 173939 616660 173940 616724
rect 174004 616660 174005 616724
rect 173939 616659 174005 616660
rect 172651 561644 172717 561645
rect 172651 561580 172652 561644
rect 172716 561580 172717 561644
rect 172651 561579 172717 561580
rect 173942 558925 174002 616659
rect 175043 568036 175109 568037
rect 175043 567972 175044 568036
rect 175108 567972 175109 568036
rect 175043 567971 175109 567972
rect 173939 558924 174005 558925
rect 173939 558860 173940 558924
rect 174004 558860 174005 558924
rect 173939 558859 174005 558860
rect 175046 547229 175106 567971
rect 175230 560285 175290 617475
rect 176334 616997 176394 647259
rect 176331 616996 176397 616997
rect 176331 616932 176332 616996
rect 176396 616932 176397 616996
rect 176331 616931 176397 616932
rect 176518 615909 176578 649979
rect 177067 641748 177133 641749
rect 177067 641684 177068 641748
rect 177132 641684 177133 641748
rect 177067 641683 177133 641684
rect 177070 621349 177130 641683
rect 177251 640388 177317 640389
rect 177251 640324 177252 640388
rect 177316 640324 177317 640388
rect 177251 640323 177317 640324
rect 177803 640388 177869 640389
rect 177803 640324 177804 640388
rect 177868 640324 177869 640388
rect 177803 640323 177869 640324
rect 177254 624613 177314 640323
rect 177435 637668 177501 637669
rect 177435 637604 177436 637668
rect 177500 637604 177501 637668
rect 177435 637603 177501 637604
rect 177251 624612 177317 624613
rect 177251 624548 177252 624612
rect 177316 624548 177317 624612
rect 177251 624547 177317 624548
rect 177067 621348 177133 621349
rect 177067 621284 177068 621348
rect 177132 621284 177133 621348
rect 177067 621283 177133 621284
rect 177251 620260 177317 620261
rect 177251 620196 177252 620260
rect 177316 620196 177317 620260
rect 177251 620195 177317 620196
rect 176515 615908 176581 615909
rect 176515 615844 176516 615908
rect 176580 615844 176581 615908
rect 176515 615843 176581 615844
rect 177067 612644 177133 612645
rect 177067 612580 177068 612644
rect 177132 612580 177133 612644
rect 177067 612579 177133 612580
rect 176699 609380 176765 609381
rect 176699 609316 176700 609380
rect 176764 609316 176765 609380
rect 176699 609315 176765 609316
rect 176702 604485 176762 609315
rect 177070 607205 177130 612579
rect 177254 610741 177314 620195
rect 177438 618085 177498 637603
rect 177619 622436 177685 622437
rect 177619 622372 177620 622436
rect 177684 622372 177685 622436
rect 177619 622371 177685 622372
rect 177435 618084 177501 618085
rect 177435 618020 177436 618084
rect 177500 618020 177501 618084
rect 177435 618019 177501 618020
rect 177435 613732 177501 613733
rect 177435 613668 177436 613732
rect 177500 613668 177501 613732
rect 177435 613667 177501 613668
rect 177251 610740 177317 610741
rect 177251 610676 177252 610740
rect 177316 610676 177317 610740
rect 177251 610675 177317 610676
rect 177438 609789 177498 613667
rect 177622 611421 177682 622371
rect 177806 614821 177866 640323
rect 178907 637124 178973 637125
rect 178907 637060 178908 637124
rect 178972 637060 178973 637124
rect 178907 637059 178973 637060
rect 178910 628965 178970 637059
rect 179091 636444 179157 636445
rect 179091 636380 179092 636444
rect 179156 636380 179157 636444
rect 179091 636379 179157 636380
rect 179094 631141 179154 636379
rect 179278 632229 179338 655011
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 633233 182414 650898
rect 185514 705798 186134 711590
rect 185514 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 186134 705798
rect 185514 705478 186134 705562
rect 185514 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 186134 705478
rect 185514 691174 186134 705242
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 633233 186134 654618
rect 189234 706758 189854 711590
rect 189234 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 189854 706758
rect 189234 706438 189854 706522
rect 189234 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 189854 706438
rect 189234 694894 189854 706202
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 633233 189854 658338
rect 192954 707718 193574 711590
rect 192954 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 193574 707718
rect 192954 707398 193574 707482
rect 192954 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 193574 707398
rect 192954 698614 193574 707162
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 633233 193574 662058
rect 196674 708678 197294 711590
rect 196674 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 197294 708678
rect 196674 708358 197294 708442
rect 196674 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 197294 708358
rect 196674 666334 197294 708122
rect 196674 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 197294 666334
rect 196674 666014 197294 666098
rect 196674 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 197294 666014
rect 196674 633233 197294 665778
rect 200394 709638 201014 711590
rect 200394 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 201014 709638
rect 200394 709318 201014 709402
rect 200394 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 201014 709318
rect 200394 670054 201014 709082
rect 200394 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 201014 670054
rect 200394 669734 201014 669818
rect 200394 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 201014 669734
rect 200394 634054 201014 669498
rect 200394 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 201014 634054
rect 200394 633734 201014 633818
rect 200394 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 201014 633734
rect 200394 633233 201014 633498
rect 204114 710598 204734 711590
rect 204114 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 204734 710598
rect 204114 710278 204734 710362
rect 204114 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 204734 710278
rect 204114 673774 204734 710042
rect 204114 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 204734 673774
rect 204114 673454 204734 673538
rect 204114 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 204734 673454
rect 204114 637774 204734 673218
rect 204114 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 204734 637774
rect 204114 637454 204734 637538
rect 204114 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 204734 637454
rect 204114 633233 204734 637218
rect 207834 711558 208454 711590
rect 207834 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 208454 711558
rect 207834 711238 208454 711322
rect 207834 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 208454 711238
rect 207834 677494 208454 711002
rect 207834 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 208454 677494
rect 207834 677174 208454 677258
rect 207834 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 208454 677174
rect 207834 641494 208454 676938
rect 207834 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 208454 641494
rect 207834 641174 208454 641258
rect 207834 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 208454 641174
rect 207834 633233 208454 640938
rect 217794 704838 218414 711590
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 633233 218414 650898
rect 221514 705798 222134 711590
rect 221514 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 222134 705798
rect 221514 705478 222134 705562
rect 221514 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 222134 705478
rect 221514 691174 222134 705242
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 633233 222134 654618
rect 225234 706758 225854 711590
rect 225234 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 225854 706758
rect 225234 706438 225854 706522
rect 225234 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 225854 706438
rect 225234 694894 225854 706202
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 633233 225854 658338
rect 228954 707718 229574 711590
rect 228954 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 229574 707718
rect 228954 707398 229574 707482
rect 228954 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 229574 707398
rect 228954 698614 229574 707162
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 633233 229574 662058
rect 232674 708678 233294 711590
rect 232674 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 233294 708678
rect 232674 708358 233294 708442
rect 232674 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 233294 708358
rect 232674 666334 233294 708122
rect 232674 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 233294 666334
rect 232674 666014 233294 666098
rect 232674 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 233294 666014
rect 232674 633233 233294 665778
rect 236394 709638 237014 711590
rect 236394 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 237014 709638
rect 236394 709318 237014 709402
rect 236394 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 237014 709318
rect 236394 670054 237014 709082
rect 236394 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 237014 670054
rect 236394 669734 237014 669818
rect 236394 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 237014 669734
rect 236394 634054 237014 669498
rect 236394 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 237014 634054
rect 236394 633734 237014 633818
rect 236394 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 237014 633734
rect 236394 633233 237014 633498
rect 240114 710598 240734 711590
rect 240114 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 240734 710598
rect 240114 710278 240734 710362
rect 240114 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 240734 710278
rect 240114 673774 240734 710042
rect 240114 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 240734 673774
rect 240114 673454 240734 673538
rect 240114 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 240734 673454
rect 240114 637774 240734 673218
rect 240114 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 240734 637774
rect 240114 637454 240734 637538
rect 240114 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 240734 637454
rect 240114 633233 240734 637218
rect 243834 711558 244454 711590
rect 243834 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 244454 711558
rect 243834 711238 244454 711322
rect 243834 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 244454 711238
rect 243834 677494 244454 711002
rect 243834 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 244454 677494
rect 243834 677174 244454 677258
rect 243834 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 244454 677174
rect 243834 641494 244454 676938
rect 243834 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 244454 641494
rect 243834 641174 244454 641258
rect 243834 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 244454 641174
rect 243834 633233 244454 640938
rect 253794 704838 254414 711590
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 249011 634132 249077 634133
rect 249011 634068 249012 634132
rect 249076 634068 249077 634132
rect 249011 634067 249077 634068
rect 249014 633725 249074 634067
rect 249011 633724 249077 633725
rect 249011 633660 249012 633724
rect 249076 633660 249077 633724
rect 249011 633659 249077 633660
rect 253794 633233 254414 650898
rect 257514 705798 258134 711590
rect 257514 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 258134 705798
rect 257514 705478 258134 705562
rect 257514 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 258134 705478
rect 257514 691174 258134 705242
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 179275 632228 179341 632229
rect 179275 632164 179276 632228
rect 179340 632164 179341 632228
rect 179275 632163 179341 632164
rect 179091 631140 179157 631141
rect 179091 631076 179092 631140
rect 179156 631076 179157 631140
rect 179091 631075 179157 631076
rect 178907 628964 178973 628965
rect 178907 628900 178908 628964
rect 178972 628900 178973 628964
rect 178907 628899 178973 628900
rect 199568 619174 199888 619206
rect 199568 618938 199610 619174
rect 199846 618938 199888 619174
rect 199568 618854 199888 618938
rect 199568 618618 199610 618854
rect 199846 618618 199888 618854
rect 199568 618586 199888 618618
rect 230288 619174 230608 619206
rect 230288 618938 230330 619174
rect 230566 618938 230608 619174
rect 230288 618854 230608 618938
rect 230288 618618 230330 618854
rect 230566 618618 230608 618854
rect 230288 618586 230608 618618
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 184208 615454 184528 615486
rect 184208 615218 184250 615454
rect 184486 615218 184528 615454
rect 184208 615134 184528 615218
rect 184208 614898 184250 615134
rect 184486 614898 184528 615134
rect 184208 614866 184528 614898
rect 214928 615454 215248 615486
rect 214928 615218 214970 615454
rect 215206 615218 215248 615454
rect 214928 615134 215248 615218
rect 214928 614898 214970 615134
rect 215206 614898 215248 615134
rect 214928 614866 215248 614898
rect 245648 615454 245968 615486
rect 245648 615218 245690 615454
rect 245926 615218 245968 615454
rect 245648 615134 245968 615218
rect 245648 614898 245690 615134
rect 245926 614898 245968 615134
rect 245648 614866 245968 614898
rect 177803 614820 177869 614821
rect 177803 614756 177804 614820
rect 177868 614756 177869 614820
rect 177803 614755 177869 614756
rect 177803 611556 177869 611557
rect 177803 611492 177804 611556
rect 177868 611492 177869 611556
rect 177803 611491 177869 611492
rect 177619 611420 177685 611421
rect 177619 611356 177620 611420
rect 177684 611356 177685 611420
rect 177619 611355 177685 611356
rect 177435 609788 177501 609789
rect 177435 609724 177436 609788
rect 177500 609724 177501 609788
rect 177435 609723 177501 609724
rect 177806 608565 177866 611491
rect 256739 611012 256805 611013
rect 256739 610948 256740 611012
rect 256804 610948 256805 611012
rect 256739 610947 256805 610948
rect 177987 610468 178053 610469
rect 177987 610404 177988 610468
rect 178052 610404 178053 610468
rect 177987 610403 178053 610404
rect 177803 608564 177869 608565
rect 177803 608500 177804 608564
rect 177868 608500 177869 608564
rect 177803 608499 177869 608500
rect 177251 608292 177317 608293
rect 177251 608228 177252 608292
rect 177316 608228 177317 608292
rect 177251 608227 177317 608228
rect 177067 607204 177133 607205
rect 177067 607140 177068 607204
rect 177132 607140 177133 607204
rect 177067 607139 177133 607140
rect 177067 606116 177133 606117
rect 177067 606052 177068 606116
rect 177132 606052 177133 606116
rect 177067 606051 177133 606052
rect 176699 604484 176765 604485
rect 176699 604420 176700 604484
rect 176764 604420 176765 604484
rect 176699 604419 176765 604420
rect 177070 596190 177130 606051
rect 177254 601765 177314 608227
rect 177803 607204 177869 607205
rect 177803 607140 177804 607204
rect 177868 607140 177869 607204
rect 177803 607139 177869 607140
rect 177619 605028 177685 605029
rect 177619 604964 177620 605028
rect 177684 604964 177685 605028
rect 177619 604963 177685 604964
rect 177435 602852 177501 602853
rect 177435 602788 177436 602852
rect 177500 602788 177501 602852
rect 177435 602787 177501 602788
rect 177251 601764 177317 601765
rect 177251 601700 177252 601764
rect 177316 601700 177317 601764
rect 177251 601699 177317 601700
rect 177070 596130 177314 596190
rect 177254 569941 177314 596130
rect 177251 569940 177317 569941
rect 177251 569876 177252 569940
rect 177316 569876 177317 569940
rect 177251 569875 177317 569876
rect 177251 569124 177317 569125
rect 177251 569060 177252 569124
rect 177316 569060 177317 569124
rect 177251 569059 177317 569060
rect 176515 564772 176581 564773
rect 176515 564708 176516 564772
rect 176580 564708 176581 564772
rect 176515 564707 176581 564708
rect 175227 560284 175293 560285
rect 175227 560220 175228 560284
rect 175292 560220 175293 560284
rect 175227 560219 175293 560220
rect 176518 549813 176578 564707
rect 177254 554709 177314 569059
rect 177251 554708 177317 554709
rect 177251 554644 177252 554708
rect 177316 554644 177317 554708
rect 177251 554643 177317 554644
rect 176515 549812 176581 549813
rect 176515 549748 176516 549812
rect 176580 549748 176581 549812
rect 176515 549747 176581 549748
rect 175043 547228 175109 547229
rect 175043 547164 175044 547228
rect 175108 547164 175109 547228
rect 175043 547163 175109 547164
rect 171834 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 172454 533494
rect 171834 533174 172454 533258
rect 171834 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 172454 533174
rect 171834 519484 172454 532938
rect 177438 532677 177498 602787
rect 177435 532676 177501 532677
rect 177435 532612 177436 532676
rect 177500 532612 177501 532676
rect 177435 532611 177501 532612
rect 177622 525741 177682 604963
rect 177619 525740 177685 525741
rect 177619 525676 177620 525740
rect 177684 525676 177685 525740
rect 177619 525675 177685 525676
rect 177806 523429 177866 607139
rect 177990 607069 178050 610403
rect 178171 609108 178237 609109
rect 178171 609044 178172 609108
rect 178236 609044 178237 609108
rect 178171 609043 178237 609044
rect 177987 607068 178053 607069
rect 177987 607004 177988 607068
rect 178052 607004 178053 607068
rect 177987 607003 178053 607004
rect 178174 605850 178234 609043
rect 177990 605790 178234 605850
rect 177990 560421 178050 605790
rect 255267 602580 255333 602581
rect 255267 602516 255268 602580
rect 255332 602516 255333 602580
rect 255267 602515 255333 602516
rect 178539 596460 178605 596461
rect 178539 596396 178540 596460
rect 178604 596396 178605 596460
rect 178539 596395 178605 596396
rect 177987 560420 178053 560421
rect 177987 560356 177988 560420
rect 178052 560356 178053 560420
rect 177987 560355 178053 560356
rect 178542 554165 178602 596395
rect 178723 586804 178789 586805
rect 178723 586740 178724 586804
rect 178788 586740 178789 586804
rect 178723 586739 178789 586740
rect 178726 556613 178786 586739
rect 199568 583174 199888 583206
rect 199568 582938 199610 583174
rect 199846 582938 199888 583174
rect 199568 582854 199888 582938
rect 199568 582618 199610 582854
rect 199846 582618 199888 582854
rect 199568 582586 199888 582618
rect 230288 583174 230608 583206
rect 230288 582938 230330 583174
rect 230566 582938 230608 583174
rect 230288 582854 230608 582938
rect 230288 582618 230330 582854
rect 230566 582618 230608 582854
rect 230288 582586 230608 582618
rect 255270 582390 255330 602515
rect 256742 598909 256802 610947
rect 256739 598908 256805 598909
rect 256739 598844 256740 598908
rect 256804 598844 256805 598908
rect 256739 598843 256805 598844
rect 256923 598772 256989 598773
rect 256923 598708 256924 598772
rect 256988 598708 256989 598772
rect 256923 598707 256989 598708
rect 256739 597956 256805 597957
rect 256739 597892 256740 597956
rect 256804 597892 256805 597956
rect 256739 597891 256805 597892
rect 254534 582330 255330 582390
rect 184208 579454 184528 579486
rect 184208 579218 184250 579454
rect 184486 579218 184528 579454
rect 184208 579134 184528 579218
rect 184208 578898 184250 579134
rect 184486 578898 184528 579134
rect 184208 578866 184528 578898
rect 214928 579454 215248 579486
rect 214928 579218 214970 579454
rect 215206 579218 215248 579454
rect 214928 579134 215248 579218
rect 214928 578898 214970 579134
rect 215206 578898 215248 579134
rect 214928 578866 215248 578898
rect 245648 579454 245968 579486
rect 245648 579218 245690 579454
rect 245926 579218 245968 579454
rect 245648 579134 245968 579218
rect 245648 578898 245690 579134
rect 245926 578898 245968 579134
rect 245648 578866 245968 578898
rect 179827 566880 179893 566881
rect 179827 566816 179828 566880
rect 179892 566816 179893 566880
rect 179827 566815 179893 566816
rect 179459 565860 179525 565861
rect 179459 565796 179460 565860
rect 179524 565796 179525 565860
rect 179459 565795 179525 565796
rect 178723 556612 178789 556613
rect 178723 556548 178724 556612
rect 178788 556548 178789 556612
rect 178723 556547 178789 556548
rect 178539 554164 178605 554165
rect 178539 554100 178540 554164
rect 178604 554100 178605 554164
rect 178539 554099 178605 554100
rect 179462 551445 179522 565795
rect 179830 563141 179890 566815
rect 179827 563140 179893 563141
rect 179827 563076 179828 563140
rect 179892 563076 179893 563140
rect 179827 563075 179893 563076
rect 180379 562528 180445 562529
rect 180379 562464 180380 562528
rect 180444 562464 180445 562528
rect 180379 562463 180445 562464
rect 180382 558789 180442 562463
rect 180563 561440 180629 561441
rect 180563 561376 180564 561440
rect 180628 561376 180629 561440
rect 180563 561375 180629 561376
rect 180566 558925 180626 561375
rect 180563 558924 180629 558925
rect 180563 558860 180564 558924
rect 180628 558860 180629 558924
rect 180563 558859 180629 558860
rect 180379 558788 180445 558789
rect 180379 558724 180380 558788
rect 180444 558724 180445 558788
rect 180379 558723 180445 558724
rect 179459 551444 179525 551445
rect 179459 551380 179460 551444
rect 179524 551380 179525 551444
rect 179459 551379 179525 551380
rect 181794 543454 182414 558575
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 177803 523428 177869 523429
rect 177803 523364 177804 523428
rect 177868 523364 177869 523428
rect 177803 523363 177869 523364
rect 171728 511174 172048 511206
rect 171728 510938 171770 511174
rect 172006 510938 172048 511174
rect 171728 510854 172048 510938
rect 171728 510618 171770 510854
rect 172006 510618 172048 510854
rect 171728 510586 172048 510618
rect 168114 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 168734 493774
rect 168114 493454 168734 493538
rect 168114 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 168734 493454
rect 168114 457774 168734 493218
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 171728 475174 172048 475206
rect 171728 474938 171770 475174
rect 172006 474938 172048 475174
rect 171728 474854 172048 474938
rect 171728 474618 171770 474854
rect 172006 474618 172048 474854
rect 171728 474586 172048 474618
rect 168114 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 168734 457774
rect 168114 457454 168734 457538
rect 168114 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 168734 457454
rect 168114 421774 168734 457218
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 171728 439174 172048 439206
rect 171728 438938 171770 439174
rect 172006 438938 172048 439174
rect 171728 438854 172048 438938
rect 171728 438618 171770 438854
rect 172006 438618 172048 438854
rect 171728 438586 172048 438618
rect 168114 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 168734 421774
rect 168114 421454 168734 421538
rect 168114 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 168734 421454
rect 168114 385774 168734 421218
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 171728 403174 172048 403206
rect 171728 402938 171770 403174
rect 172006 402938 172048 403174
rect 171728 402854 172048 402938
rect 171728 402618 171770 402854
rect 172006 402618 172048 402854
rect 171728 402586 172048 402618
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 168114 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 168734 385774
rect 168114 385454 168734 385538
rect 168114 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 168734 385454
rect 168114 349774 168734 385218
rect 168114 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 168734 349774
rect 168114 349454 168734 349538
rect 168114 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 168734 349454
rect 168114 313774 168734 349218
rect 168114 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 168734 313774
rect 168114 313454 168734 313538
rect 168114 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 168734 313454
rect 168114 277774 168734 313218
rect 168114 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 168734 277774
rect 168114 277454 168734 277538
rect 168114 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 168734 277454
rect 168114 241774 168734 277218
rect 168114 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 168734 241774
rect 168114 241454 168734 241538
rect 168114 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 168734 241454
rect 168114 205774 168734 241218
rect 168114 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 168734 205774
rect 168114 205454 168734 205538
rect 168114 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 168734 205454
rect 168114 169774 168734 205218
rect 168114 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 168734 169774
rect 168114 169454 168734 169538
rect 168114 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 168734 169454
rect 168114 133774 168734 169218
rect 168114 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 168734 133774
rect 168114 133454 168734 133538
rect 168114 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 168734 133454
rect 168114 97774 168734 133218
rect 168114 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 168734 97774
rect 168114 97454 168734 97538
rect 168114 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 168734 97454
rect 168114 61774 168734 97218
rect 168114 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 168734 61774
rect 168114 61454 168734 61538
rect 168114 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 168734 61454
rect 168114 25774 168734 61218
rect 168114 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 168734 25774
rect 168114 25454 168734 25538
rect 168114 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 168734 25454
rect 168114 -6106 168734 25218
rect 168114 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 168734 -6106
rect 168114 -6426 168734 -6342
rect 168114 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 168734 -6426
rect 168114 -7654 168734 -6662
rect 171834 389494 172454 389988
rect 171834 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 172454 389494
rect 171834 389174 172454 389258
rect 171834 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 172454 389174
rect 171834 353494 172454 388938
rect 171834 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 172454 353494
rect 171834 353174 172454 353258
rect 171834 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 172454 353174
rect 171834 317494 172454 352938
rect 171834 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 172454 317494
rect 171834 317174 172454 317258
rect 171834 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 172454 317174
rect 171834 281494 172454 316938
rect 171834 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 172454 281494
rect 171834 281174 172454 281258
rect 171834 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 172454 281174
rect 171834 245494 172454 280938
rect 171834 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 172454 245494
rect 171834 245174 172454 245258
rect 171834 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 172454 245174
rect 171834 209494 172454 244938
rect 171834 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 172454 209494
rect 171834 209174 172454 209258
rect 171834 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 172454 209174
rect 171834 173494 172454 208938
rect 171834 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 172454 173494
rect 171834 173174 172454 173258
rect 171834 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 172454 173174
rect 171834 137494 172454 172938
rect 171834 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 172454 137494
rect 171834 137174 172454 137258
rect 171834 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 172454 137174
rect 171834 101494 172454 136938
rect 171834 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 172454 101494
rect 171834 101174 172454 101258
rect 171834 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 172454 101174
rect 171834 65494 172454 100938
rect 171834 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 172454 65494
rect 171834 65174 172454 65258
rect 171834 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 172454 65174
rect 171834 29494 172454 64938
rect 171834 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 172454 29494
rect 171834 29174 172454 29258
rect 171834 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 172454 29174
rect 171834 -7066 172454 28938
rect 171834 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 172454 -7066
rect 171834 -7386 172454 -7302
rect 171834 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 172454 -7386
rect 171834 -7654 172454 -7622
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -7654 182414 -902
rect 185514 547174 186134 558575
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 189234 550894 189854 558575
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 187088 471454 187408 471486
rect 187088 471218 187130 471454
rect 187366 471218 187408 471454
rect 187088 471134 187408 471218
rect 187088 470898 187130 471134
rect 187366 470898 187408 471134
rect 187088 470866 187408 470898
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 187088 435454 187408 435486
rect 187088 435218 187130 435454
rect 187366 435218 187408 435454
rect 187088 435134 187408 435218
rect 187088 434898 187130 435134
rect 187366 434898 187408 435134
rect 187088 434866 187408 434898
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 187088 399454 187408 399486
rect 187088 399218 187130 399454
rect 187366 399218 187408 399454
rect 187088 399134 187408 399218
rect 187088 398898 187130 399134
rect 187366 398898 187408 399134
rect 187088 398866 187408 398898
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -1306 186134 6618
rect 185514 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 186134 -1306
rect 185514 -1626 186134 -1542
rect 185514 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 186134 -1626
rect 185514 -7654 186134 -1862
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -2266 189854 10338
rect 189234 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 189854 -2266
rect 189234 -2586 189854 -2502
rect 189234 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 189854 -2586
rect 189234 -7654 189854 -2822
rect 192954 554614 193574 558575
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 192954 -3226 193574 14058
rect 192954 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 193574 -3226
rect 192954 -3546 193574 -3462
rect 192954 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 193574 -3546
rect 192954 -7654 193574 -3782
rect 196674 558334 197294 558575
rect 196674 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 197294 558334
rect 196674 558014 197294 558098
rect 196674 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 197294 558014
rect 196674 522334 197294 557778
rect 196674 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 197294 522334
rect 232674 558334 233294 558575
rect 232674 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 233294 558334
rect 232674 558014 233294 558098
rect 232674 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 233294 558014
rect 232674 522121 233294 557778
rect 196674 522014 197294 522098
rect 196674 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 197294 522014
rect 196674 486334 197294 521778
rect 254534 520981 254594 582330
rect 256742 572797 256802 597891
rect 256926 575517 256986 598707
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257107 575924 257173 575925
rect 257107 575860 257108 575924
rect 257172 575860 257173 575924
rect 257107 575859 257173 575860
rect 256923 575516 256989 575517
rect 256923 575452 256924 575516
rect 256988 575452 256989 575516
rect 256923 575451 256989 575452
rect 256739 572796 256805 572797
rect 256739 572732 256740 572796
rect 256804 572732 256805 572796
rect 256739 572731 256805 572732
rect 257110 572661 257170 575859
rect 257107 572660 257173 572661
rect 257107 572596 257108 572660
rect 257172 572596 257173 572660
rect 257107 572595 257173 572596
rect 257107 571844 257173 571845
rect 257107 571780 257108 571844
rect 257172 571780 257173 571844
rect 257107 571779 257173 571780
rect 256923 571028 256989 571029
rect 256923 570964 256924 571028
rect 256988 570964 256989 571028
rect 256923 570963 256989 570964
rect 255819 560692 255885 560693
rect 255819 560628 255820 560692
rect 255884 560628 255885 560692
rect 255819 560627 255885 560628
rect 255083 560556 255149 560557
rect 255083 560492 255084 560556
rect 255148 560492 255149 560556
rect 255083 560491 255149 560492
rect 255086 546413 255146 560491
rect 255083 546412 255149 546413
rect 255083 546348 255084 546412
rect 255148 546348 255149 546412
rect 255083 546347 255149 546348
rect 255822 534989 255882 560627
rect 256926 558245 256986 570963
rect 256923 558244 256989 558245
rect 256923 558180 256924 558244
rect 256988 558180 256989 558244
rect 256923 558179 256989 558180
rect 255819 534988 255885 534989
rect 255819 534924 255820 534988
rect 255884 534924 255885 534988
rect 255819 534923 255885 534924
rect 257110 526149 257170 571779
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257107 526148 257173 526149
rect 257107 526084 257108 526148
rect 257172 526084 257173 526148
rect 257107 526083 257173 526084
rect 257514 522121 258134 546618
rect 261234 706758 261854 711590
rect 261234 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 261854 706758
rect 261234 706438 261854 706522
rect 261234 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 261854 706438
rect 261234 694894 261854 706202
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 522121 261854 550338
rect 264954 707718 265574 711590
rect 264954 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 265574 707718
rect 264954 707398 265574 707482
rect 264954 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 265574 707398
rect 264954 698614 265574 707162
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 522121 265574 554058
rect 268674 708678 269294 711590
rect 268674 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 269294 708678
rect 268674 708358 269294 708442
rect 268674 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 269294 708358
rect 268674 666334 269294 708122
rect 268674 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 269294 666334
rect 268674 666014 269294 666098
rect 268674 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 269294 666014
rect 268674 630334 269294 665778
rect 268674 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 269294 630334
rect 268674 630014 269294 630098
rect 268674 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 269294 630014
rect 268674 594334 269294 629778
rect 268674 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 269294 594334
rect 268674 594014 269294 594098
rect 268674 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 269294 594014
rect 268674 558334 269294 593778
rect 268674 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 269294 558334
rect 268674 558014 269294 558098
rect 268674 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 269294 558014
rect 268674 522121 269294 557778
rect 272394 709638 273014 711590
rect 272394 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 273014 709638
rect 272394 709318 273014 709402
rect 272394 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 273014 709318
rect 272394 670054 273014 709082
rect 272394 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 273014 670054
rect 272394 669734 273014 669818
rect 272394 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 273014 669734
rect 272394 634054 273014 669498
rect 272394 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 273014 634054
rect 272394 633734 273014 633818
rect 272394 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 273014 633734
rect 272394 598054 273014 633498
rect 272394 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 273014 598054
rect 272394 597734 273014 597818
rect 272394 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 273014 597734
rect 272394 562054 273014 597498
rect 272394 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 273014 562054
rect 272394 561734 273014 561818
rect 272394 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 273014 561734
rect 272394 526054 273014 561498
rect 272394 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 273014 526054
rect 272394 525734 273014 525818
rect 272394 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 273014 525734
rect 272394 522121 273014 525498
rect 276114 710598 276734 711590
rect 276114 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 276734 710598
rect 276114 710278 276734 710362
rect 276114 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 276734 710278
rect 276114 673774 276734 710042
rect 276114 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 276734 673774
rect 276114 673454 276734 673538
rect 276114 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 276734 673454
rect 276114 637774 276734 673218
rect 276114 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 276734 637774
rect 276114 637454 276734 637538
rect 276114 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 276734 637454
rect 276114 601774 276734 637218
rect 276114 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 276734 601774
rect 276114 601454 276734 601538
rect 276114 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 276734 601454
rect 276114 565774 276734 601218
rect 276114 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 276734 565774
rect 276114 565454 276734 565538
rect 276114 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 276734 565454
rect 276114 529774 276734 565218
rect 276114 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 276734 529774
rect 276114 529454 276734 529538
rect 276114 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 276734 529454
rect 276114 522121 276734 529218
rect 279834 711558 280454 711590
rect 279834 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 280454 711558
rect 279834 711238 280454 711322
rect 279834 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 280454 711238
rect 279834 677494 280454 711002
rect 279834 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 280454 677494
rect 279834 677174 280454 677258
rect 279834 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 280454 677174
rect 279834 641494 280454 676938
rect 279834 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 280454 641494
rect 279834 641174 280454 641258
rect 279834 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 280454 641174
rect 279834 605494 280454 640938
rect 289794 704838 290414 711590
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 288387 622436 288453 622437
rect 288387 622372 288388 622436
rect 288452 622372 288453 622436
rect 288387 622371 288453 622372
rect 287099 617540 287165 617541
rect 287099 617476 287100 617540
rect 287164 617476 287165 617540
rect 287099 617475 287165 617476
rect 282131 615908 282197 615909
rect 282131 615844 282132 615908
rect 282196 615844 282197 615908
rect 282131 615843 282197 615844
rect 280659 613460 280725 613461
rect 280659 613396 280660 613460
rect 280724 613396 280725 613460
rect 280659 613395 280725 613396
rect 279834 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 280454 605494
rect 279834 605174 280454 605258
rect 279834 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 280454 605174
rect 279834 569494 280454 604938
rect 279834 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 280454 569494
rect 279834 569174 280454 569258
rect 279834 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 280454 569174
rect 279834 533494 280454 568938
rect 279834 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 280454 533494
rect 279834 533174 280454 533258
rect 279834 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 280454 533174
rect 279834 522121 280454 532938
rect 280662 525605 280722 613395
rect 281027 592244 281093 592245
rect 281027 592180 281028 592244
rect 281092 592180 281093 592244
rect 281027 592179 281093 592180
rect 280659 525604 280725 525605
rect 280659 525540 280660 525604
rect 280724 525540 280725 525604
rect 280659 525539 280725 525540
rect 281030 524245 281090 592179
rect 282134 539205 282194 615843
rect 284891 611828 284957 611829
rect 284891 611764 284892 611828
rect 284956 611764 284957 611828
rect 284891 611763 284957 611764
rect 283971 593876 284037 593877
rect 283971 593812 283972 593876
rect 284036 593812 284037 593876
rect 283971 593811 284037 593812
rect 283787 589660 283853 589661
rect 283787 589596 283788 589660
rect 283852 589596 283853 589660
rect 283787 589595 283853 589596
rect 283419 582452 283485 582453
rect 283419 582388 283420 582452
rect 283484 582388 283485 582452
rect 283419 582387 283485 582388
rect 282867 546548 282933 546549
rect 282867 546484 282868 546548
rect 282932 546484 282933 546548
rect 282867 546483 282933 546484
rect 282131 539204 282197 539205
rect 282131 539140 282132 539204
rect 282196 539140 282197 539204
rect 282131 539139 282197 539140
rect 282870 525197 282930 546483
rect 282867 525196 282933 525197
rect 282867 525132 282868 525196
rect 282932 525132 282933 525196
rect 282867 525131 282933 525132
rect 281027 524244 281093 524245
rect 281027 524180 281028 524244
rect 281092 524180 281093 524244
rect 281027 524179 281093 524180
rect 283422 520981 283482 582387
rect 283603 581636 283669 581637
rect 283603 581572 283604 581636
rect 283668 581572 283669 581636
rect 283603 581571 283669 581572
rect 283606 523973 283666 581571
rect 283790 537845 283850 589595
rect 283974 547637 284034 593811
rect 283971 547636 284037 547637
rect 283971 547572 283972 547636
rect 284036 547572 284037 547636
rect 283971 547571 284037 547572
rect 284894 546277 284954 611763
rect 286179 610468 286245 610469
rect 286179 610404 286180 610468
rect 286244 610404 286245 610468
rect 286179 610403 286245 610404
rect 285259 591428 285325 591429
rect 285259 591364 285260 591428
rect 285324 591364 285325 591428
rect 285259 591363 285325 591364
rect 285075 583268 285141 583269
rect 285075 583204 285076 583268
rect 285140 583204 285141 583268
rect 285075 583203 285141 583204
rect 284891 546276 284957 546277
rect 284891 546212 284892 546276
rect 284956 546212 284957 546276
rect 284891 546211 284957 546212
rect 283787 537844 283853 537845
rect 283787 537780 283788 537844
rect 283852 537780 283853 537844
rect 283787 537779 283853 537780
rect 285078 525333 285138 583203
rect 285262 542061 285322 591363
rect 285443 574292 285509 574293
rect 285443 574228 285444 574292
rect 285508 574228 285509 574292
rect 285443 574227 285509 574228
rect 285259 542060 285325 542061
rect 285259 541996 285260 542060
rect 285324 541996 285325 542060
rect 285259 541995 285325 541996
rect 285075 525332 285141 525333
rect 285075 525268 285076 525332
rect 285140 525268 285141 525332
rect 285075 525267 285141 525268
rect 285446 525197 285506 574227
rect 286182 537709 286242 610403
rect 286363 584084 286429 584085
rect 286363 584020 286364 584084
rect 286428 584020 286429 584084
rect 286363 584019 286429 584020
rect 286179 537708 286245 537709
rect 286179 537644 286180 537708
rect 286244 537644 286245 537708
rect 286179 537643 286245 537644
rect 286366 529549 286426 584019
rect 287102 578237 287162 617475
rect 287651 603668 287717 603669
rect 287651 603604 287652 603668
rect 287716 603604 287717 603668
rect 287651 603603 287717 603604
rect 287099 578236 287165 578237
rect 287099 578172 287100 578236
rect 287164 578172 287165 578236
rect 287099 578171 287165 578172
rect 286547 571300 286613 571301
rect 286547 571236 286548 571300
rect 286612 571236 286613 571300
rect 286547 571235 286613 571236
rect 286550 546141 286610 571235
rect 286547 546140 286613 546141
rect 286547 546076 286548 546140
rect 286612 546076 286613 546140
rect 286547 546075 286613 546076
rect 287654 533765 287714 603603
rect 287835 586532 287901 586533
rect 287835 586468 287836 586532
rect 287900 586468 287901 586532
rect 287835 586467 287901 586468
rect 287651 533764 287717 533765
rect 287651 533700 287652 533764
rect 287716 533700 287717 533764
rect 287651 533699 287717 533700
rect 286363 529548 286429 529549
rect 286363 529484 286364 529548
rect 286428 529484 286429 529548
rect 286363 529483 286429 529484
rect 285443 525196 285509 525197
rect 285443 525132 285444 525196
rect 285508 525132 285509 525196
rect 285443 525131 285509 525132
rect 283603 523972 283669 523973
rect 283603 523908 283604 523972
rect 283668 523908 283669 523972
rect 283603 523907 283669 523908
rect 287838 521253 287898 586467
rect 288203 584900 288269 584901
rect 288203 584836 288204 584900
rect 288268 584836 288269 584900
rect 288203 584835 288269 584836
rect 288019 577556 288085 577557
rect 288019 577492 288020 577556
rect 288084 577492 288085 577556
rect 288019 577491 288085 577492
rect 288022 526693 288082 577491
rect 288206 546141 288266 584835
rect 288390 564501 288450 622371
rect 289794 615454 290414 650898
rect 293514 705798 294134 711590
rect 293514 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 294134 705798
rect 293514 705478 294134 705562
rect 293514 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 294134 705478
rect 293514 691174 294134 705242
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 291883 639436 291949 639437
rect 291883 639372 291884 639436
rect 291948 639372 291949 639436
rect 291883 639371 291949 639372
rect 291699 637940 291765 637941
rect 291699 637876 291700 637940
rect 291764 637876 291765 637940
rect 291699 637875 291765 637876
rect 291147 626516 291213 626517
rect 291147 626452 291148 626516
rect 291212 626452 291213 626516
rect 291147 626451 291213 626452
rect 290595 619172 290661 619173
rect 290595 619108 290596 619172
rect 290660 619108 290661 619172
rect 290595 619107 290661 619108
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 288571 615092 288637 615093
rect 288571 615028 288572 615092
rect 288636 615028 288637 615092
rect 288571 615027 288637 615028
rect 288387 564500 288453 564501
rect 288387 564436 288388 564500
rect 288452 564436 288453 564500
rect 288387 564435 288453 564436
rect 288574 563141 288634 615027
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289307 588164 289373 588165
rect 289307 588100 289308 588164
rect 289372 588100 289373 588164
rect 289307 588099 289373 588100
rect 289123 564772 289189 564773
rect 289123 564708 289124 564772
rect 289188 564708 289189 564772
rect 289123 564707 289189 564708
rect 288939 563684 289005 563685
rect 288939 563620 288940 563684
rect 289004 563620 289005 563684
rect 288939 563619 289005 563620
rect 288571 563140 288637 563141
rect 288571 563076 288572 563140
rect 288636 563076 288637 563140
rect 288571 563075 288637 563076
rect 288387 556204 288453 556205
rect 288387 556140 288388 556204
rect 288452 556140 288453 556204
rect 288387 556139 288453 556140
rect 288203 546140 288269 546141
rect 288203 546076 288204 546140
rect 288268 546076 288269 546140
rect 288203 546075 288269 546076
rect 288019 526692 288085 526693
rect 288019 526628 288020 526692
rect 288084 526628 288085 526692
rect 288019 526627 288085 526628
rect 288390 523565 288450 556139
rect 288571 549132 288637 549133
rect 288571 549068 288572 549132
rect 288636 549068 288637 549132
rect 288571 549067 288637 549068
rect 288574 541925 288634 549067
rect 288571 541924 288637 541925
rect 288571 541860 288572 541924
rect 288636 541860 288637 541924
rect 288571 541859 288637 541860
rect 288942 524109 289002 563619
rect 289126 525469 289186 564707
rect 289310 557157 289370 588099
rect 289491 579868 289557 579869
rect 289491 579804 289492 579868
rect 289556 579804 289557 579868
rect 289491 579803 289557 579804
rect 289307 557156 289373 557157
rect 289307 557092 289308 557156
rect 289372 557092 289373 557156
rect 289307 557091 289373 557092
rect 289494 548997 289554 579803
rect 289794 579454 290414 614898
rect 290598 585173 290658 619107
rect 290779 608564 290845 608565
rect 290779 608500 290780 608564
rect 290844 608500 290845 608564
rect 290779 608499 290845 608500
rect 290595 585172 290661 585173
rect 290595 585108 290596 585172
rect 290660 585108 290661 585172
rect 290595 585107 290661 585108
rect 290782 580957 290842 608499
rect 290963 585716 291029 585717
rect 290963 585652 290964 585716
rect 291028 585652 291029 585716
rect 290963 585651 291029 585652
rect 290966 581093 291026 585651
rect 290963 581092 291029 581093
rect 290963 581028 290964 581092
rect 291028 581028 291029 581092
rect 290963 581027 291029 581028
rect 290779 580956 290845 580957
rect 290779 580892 290780 580956
rect 290844 580892 290845 580956
rect 290779 580891 290845 580892
rect 290963 580820 291029 580821
rect 290963 580756 290964 580820
rect 291028 580756 291029 580820
rect 290963 580755 291029 580756
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289491 548996 289557 548997
rect 289491 548932 289492 548996
rect 289556 548932 289557 548996
rect 289491 548931 289557 548932
rect 289794 543454 290414 578898
rect 290595 578372 290661 578373
rect 290595 578308 290596 578372
rect 290660 578308 290661 578372
rect 290595 578307 290661 578308
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289123 525468 289189 525469
rect 289123 525404 289124 525468
rect 289188 525404 289189 525468
rect 289123 525403 289189 525404
rect 288939 524108 289005 524109
rect 288939 524044 288940 524108
rect 289004 524044 289005 524108
rect 288939 524043 289005 524044
rect 288387 523564 288453 523565
rect 288387 523500 288388 523564
rect 288452 523500 288453 523564
rect 288387 523499 288453 523500
rect 289794 522121 290414 542898
rect 290598 537709 290658 578307
rect 290966 549133 291026 580755
rect 291150 562325 291210 626451
rect 291702 614821 291762 637875
rect 291886 615909 291946 639371
rect 292067 637940 292133 637941
rect 292067 637876 292068 637940
rect 292132 637876 292133 637940
rect 292067 637875 292133 637876
rect 292070 621621 292130 637875
rect 292067 621620 292133 621621
rect 292067 621556 292068 621620
rect 292132 621556 292133 621620
rect 292067 621555 292133 621556
rect 293514 619174 294134 654618
rect 297234 706758 297854 711590
rect 297234 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 297854 706758
rect 297234 706438 297854 706522
rect 297234 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 297854 706438
rect 297234 694894 297854 706202
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 296851 645420 296917 645421
rect 296851 645356 296852 645420
rect 296916 645356 296917 645420
rect 296851 645355 296917 645356
rect 294827 641204 294893 641205
rect 294827 641140 294828 641204
rect 294892 641140 294893 641204
rect 294827 641139 294893 641140
rect 294643 639436 294709 639437
rect 294643 639372 294644 639436
rect 294708 639372 294709 639436
rect 294643 639371 294709 639372
rect 294459 638076 294525 638077
rect 294459 638012 294460 638076
rect 294524 638012 294525 638076
rect 294459 638011 294525 638012
rect 294462 620805 294522 638011
rect 294646 623253 294706 639371
rect 294830 624069 294890 641139
rect 296854 640250 296914 645355
rect 297035 643652 297101 643653
rect 297035 643588 297036 643652
rect 297100 643588 297101 643652
rect 297035 643587 297101 643588
rect 297038 640253 297098 643587
rect 296486 640190 296914 640250
rect 297035 640252 297101 640253
rect 296486 635490 296546 640190
rect 297035 640188 297036 640252
rect 297100 640188 297101 640252
rect 297035 640187 297101 640188
rect 296851 639708 296917 639709
rect 296851 639644 296852 639708
rect 296916 639644 296917 639708
rect 296851 639643 296917 639644
rect 296667 635492 296733 635493
rect 296667 635490 296668 635492
rect 296486 635430 296668 635490
rect 296667 635428 296668 635430
rect 296732 635428 296733 635492
rect 296667 635427 296733 635428
rect 296483 635356 296549 635357
rect 296483 635292 296484 635356
rect 296548 635292 296549 635356
rect 296483 635291 296549 635292
rect 296486 625170 296546 635291
rect 296854 625701 296914 639643
rect 296851 625700 296917 625701
rect 296851 625636 296852 625700
rect 296916 625636 296917 625700
rect 296851 625635 296917 625636
rect 296486 625110 297098 625170
rect 297038 624613 297098 625110
rect 297035 624612 297101 624613
rect 297035 624548 297036 624612
rect 297100 624548 297101 624612
rect 297035 624547 297101 624548
rect 294827 624068 294893 624069
rect 294827 624004 294828 624068
rect 294892 624004 294893 624068
rect 294827 624003 294893 624004
rect 294643 623252 294709 623253
rect 294643 623188 294644 623252
rect 294708 623188 294709 623252
rect 294643 623187 294709 623188
rect 297234 622894 297854 658338
rect 300954 707718 301574 711590
rect 300954 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 301574 707718
rect 300954 707398 301574 707482
rect 300954 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 301574 707398
rect 300954 698614 301574 707162
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 633233 301574 662058
rect 304674 708678 305294 711590
rect 304674 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 305294 708678
rect 304674 708358 305294 708442
rect 304674 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 305294 708358
rect 304674 666334 305294 708122
rect 304674 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 305294 666334
rect 304674 666014 305294 666098
rect 304674 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 305294 666014
rect 304674 633233 305294 665778
rect 308394 709638 309014 711590
rect 308394 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 309014 709638
rect 308394 709318 309014 709402
rect 308394 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 309014 709318
rect 308394 670054 309014 709082
rect 308394 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 309014 670054
rect 308394 669734 309014 669818
rect 308394 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 309014 669734
rect 308394 634054 309014 669498
rect 308394 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 309014 634054
rect 308394 633734 309014 633818
rect 308394 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 309014 633734
rect 308394 633233 309014 633498
rect 312114 710598 312734 711590
rect 312114 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 312734 710598
rect 312114 710278 312734 710362
rect 312114 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 312734 710278
rect 312114 673774 312734 710042
rect 312114 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 312734 673774
rect 312114 673454 312734 673538
rect 312114 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 312734 673454
rect 312114 637774 312734 673218
rect 312114 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 312734 637774
rect 312114 637454 312734 637538
rect 312114 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 312734 637454
rect 312114 633233 312734 637218
rect 315834 711558 316454 711590
rect 315834 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 316454 711558
rect 315834 711238 316454 711322
rect 315834 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 316454 711238
rect 315834 677494 316454 711002
rect 315834 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 316454 677494
rect 315834 677174 316454 677258
rect 315834 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 316454 677174
rect 315834 641494 316454 676938
rect 315834 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 316454 641494
rect 315834 641174 316454 641258
rect 315834 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 316454 641174
rect 315834 633233 316454 640938
rect 325794 704838 326414 711590
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 633233 326414 650898
rect 329514 705798 330134 711590
rect 329514 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 330134 705798
rect 329514 705478 330134 705562
rect 329514 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 330134 705478
rect 329514 691174 330134 705242
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 633233 330134 654618
rect 333234 706758 333854 711590
rect 333234 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 333854 706758
rect 333234 706438 333854 706522
rect 333234 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 333854 706438
rect 333234 694894 333854 706202
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 633233 333854 658338
rect 336954 707718 337574 711590
rect 336954 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 337574 707718
rect 336954 707398 337574 707482
rect 336954 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 337574 707398
rect 336954 698614 337574 707162
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 633233 337574 662058
rect 340674 708678 341294 711590
rect 340674 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 341294 708678
rect 340674 708358 341294 708442
rect 340674 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 341294 708358
rect 340674 666334 341294 708122
rect 340674 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 341294 666334
rect 340674 666014 341294 666098
rect 340674 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 341294 666014
rect 340674 633233 341294 665778
rect 344394 709638 345014 711590
rect 344394 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 345014 709638
rect 344394 709318 345014 709402
rect 344394 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 345014 709318
rect 344394 670054 345014 709082
rect 344394 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 345014 670054
rect 344394 669734 345014 669818
rect 344394 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 345014 669734
rect 344394 634054 345014 669498
rect 344394 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 345014 634054
rect 344394 633734 345014 633818
rect 344394 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 345014 633734
rect 344394 633233 345014 633498
rect 348114 710598 348734 711590
rect 348114 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 348734 710598
rect 348114 710278 348734 710362
rect 348114 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 348734 710278
rect 348114 673774 348734 710042
rect 348114 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 348734 673774
rect 348114 673454 348734 673538
rect 348114 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 348734 673454
rect 348114 637774 348734 673218
rect 348114 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 348734 637774
rect 348114 637454 348734 637538
rect 348114 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 348734 637454
rect 348114 633233 348734 637218
rect 351834 711558 352454 711590
rect 351834 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 352454 711558
rect 351834 711238 352454 711322
rect 351834 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 352454 711238
rect 351834 677494 352454 711002
rect 351834 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 352454 677494
rect 351834 677174 352454 677258
rect 351834 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 352454 677174
rect 351834 641494 352454 676938
rect 351834 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 352454 641494
rect 351834 641174 352454 641258
rect 351834 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 352454 641174
rect 351834 633233 352454 640938
rect 361794 704838 362414 711590
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 633233 362414 650898
rect 365514 705798 366134 711590
rect 365514 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 366134 705798
rect 365514 705478 366134 705562
rect 365514 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 366134 705478
rect 365514 691174 366134 705242
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 634540 366134 654618
rect 369234 706758 369854 711590
rect 369234 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 369854 706758
rect 369234 706438 369854 706522
rect 369234 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 369854 706438
rect 369234 694894 369854 706202
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 633233 369854 658338
rect 372954 707718 373574 711590
rect 372954 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 373574 707718
rect 372954 707398 373574 707482
rect 372954 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 373574 707398
rect 372954 698614 373574 707162
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 633233 373574 662058
rect 376674 708678 377294 711590
rect 376674 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 377294 708678
rect 376674 708358 377294 708442
rect 376674 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 377294 708358
rect 376674 666334 377294 708122
rect 376674 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 377294 666334
rect 376674 666014 377294 666098
rect 376674 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 377294 666014
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 294459 620804 294525 620805
rect 294459 620740 294460 620804
rect 294524 620740 294525 620804
rect 294459 620739 294525 620740
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 291883 615908 291949 615909
rect 291883 615844 291884 615908
rect 291948 615844 291949 615908
rect 291883 615843 291949 615844
rect 291699 614820 291765 614821
rect 291699 614756 291700 614820
rect 291764 614756 291765 614820
rect 291699 614755 291765 614756
rect 292619 606116 292685 606117
rect 292619 606052 292620 606116
rect 292684 606052 292685 606116
rect 292619 606051 292685 606052
rect 291699 594692 291765 594693
rect 291699 594628 291700 594692
rect 291764 594628 291765 594692
rect 291699 594627 291765 594628
rect 291147 562324 291213 562325
rect 291147 562260 291148 562324
rect 291212 562260 291213 562324
rect 291147 562259 291213 562260
rect 291147 551716 291213 551717
rect 291147 551652 291148 551716
rect 291212 551652 291213 551716
rect 291147 551651 291213 551652
rect 290963 549132 291029 549133
rect 290963 549068 290964 549132
rect 291028 549068 291029 549132
rect 290963 549067 291029 549068
rect 290595 537708 290661 537709
rect 290595 537644 290596 537708
rect 290660 537644 290661 537708
rect 290595 537643 290661 537644
rect 291150 526829 291210 551651
rect 291702 536349 291762 594627
rect 292067 576740 292133 576741
rect 292067 576676 292068 576740
rect 292132 576676 292133 576740
rect 292067 576675 292133 576676
rect 291883 575108 291949 575109
rect 291883 575044 291884 575108
rect 291948 575044 291949 575108
rect 291883 575043 291949 575044
rect 291699 536348 291765 536349
rect 291699 536284 291700 536348
rect 291764 536284 291765 536348
rect 291699 536283 291765 536284
rect 291147 526828 291213 526829
rect 291147 526764 291148 526828
rect 291212 526764 291213 526828
rect 291147 526763 291213 526764
rect 287835 521252 287901 521253
rect 287835 521188 287836 521252
rect 287900 521188 287901 521252
rect 287835 521187 287901 521188
rect 254531 520980 254597 520981
rect 254531 520916 254532 520980
rect 254596 520916 254597 520980
rect 254531 520915 254597 520916
rect 283419 520980 283485 520981
rect 283419 520916 283420 520980
rect 283484 520916 283485 520980
rect 283419 520915 283485 520916
rect 291886 520437 291946 575043
rect 292070 551581 292130 576675
rect 292622 568581 292682 606051
rect 293514 583174 294134 618618
rect 295379 618356 295445 618357
rect 295379 618292 295380 618356
rect 295444 618292 295445 618356
rect 295379 618291 295445 618292
rect 294827 614276 294893 614277
rect 294827 614212 294828 614276
rect 294892 614212 294893 614276
rect 294827 614211 294893 614212
rect 294459 612644 294525 612645
rect 294459 612580 294460 612644
rect 294524 612580 294525 612644
rect 294459 612579 294525 612580
rect 294462 590613 294522 612579
rect 294643 609380 294709 609381
rect 294643 609316 294644 609380
rect 294708 609316 294709 609380
rect 294643 609315 294709 609316
rect 294459 590612 294525 590613
rect 294459 590548 294460 590612
rect 294524 590548 294525 590612
rect 294459 590547 294525 590548
rect 294646 589253 294706 609315
rect 294830 601085 294890 614211
rect 295011 601220 295077 601221
rect 295011 601156 295012 601220
rect 295076 601156 295077 601220
rect 295011 601155 295077 601156
rect 294827 601084 294893 601085
rect 294827 601020 294828 601084
rect 294892 601020 294893 601084
rect 294827 601019 294893 601020
rect 294827 590340 294893 590341
rect 294827 590276 294828 590340
rect 294892 590276 294893 590340
rect 294827 590275 294893 590276
rect 294643 589252 294709 589253
rect 294643 589188 294644 589252
rect 294708 589188 294709 589252
rect 294643 589187 294709 589188
rect 294459 588980 294525 588981
rect 294459 588916 294460 588980
rect 294524 588916 294525 588980
rect 294459 588915 294525 588916
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293171 579188 293237 579189
rect 293171 579124 293172 579188
rect 293236 579124 293237 579188
rect 293171 579123 293237 579124
rect 292619 568580 292685 568581
rect 292619 568516 292620 568580
rect 292684 568516 292685 568580
rect 292619 568515 292685 568516
rect 292987 568308 293053 568309
rect 292987 568244 292988 568308
rect 293052 568244 293053 568308
rect 292987 568243 293053 568244
rect 292251 562596 292317 562597
rect 292251 562532 292252 562596
rect 292316 562532 292317 562596
rect 292251 562531 292317 562532
rect 292067 551580 292133 551581
rect 292067 551516 292068 551580
rect 292132 551516 292133 551580
rect 292067 551515 292133 551516
rect 292254 547501 292314 562531
rect 292251 547500 292317 547501
rect 292251 547436 292252 547500
rect 292316 547436 292317 547500
rect 292251 547435 292317 547436
rect 292619 546548 292685 546549
rect 292619 546484 292620 546548
rect 292684 546484 292685 546548
rect 292619 546483 292685 546484
rect 292622 522341 292682 546483
rect 292990 543421 293050 568243
rect 293174 547501 293234 579123
rect 293171 547500 293237 547501
rect 293171 547436 293172 547500
rect 293236 547436 293237 547500
rect 293171 547435 293237 547436
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 292987 543420 293053 543421
rect 292987 543356 292988 543420
rect 293052 543356 293053 543420
rect 292987 543355 293053 543356
rect 292619 522340 292685 522341
rect 292619 522276 292620 522340
rect 292684 522276 292685 522340
rect 292619 522275 292685 522276
rect 293514 522121 294134 546618
rect 294462 541925 294522 588915
rect 294643 587348 294709 587349
rect 294643 587284 294644 587348
rect 294708 587284 294709 587348
rect 294643 587283 294709 587284
rect 294646 557429 294706 587283
rect 294830 569941 294890 590275
rect 295014 586533 295074 601155
rect 295382 597549 295442 618291
rect 295931 616724 295997 616725
rect 295931 616660 295932 616724
rect 295996 616660 295997 616724
rect 295931 616659 295997 616660
rect 295747 600404 295813 600405
rect 295747 600340 295748 600404
rect 295812 600340 295813 600404
rect 295747 600339 295813 600340
rect 295379 597548 295445 597549
rect 295379 597484 295380 597548
rect 295444 597484 295445 597548
rect 295379 597483 295445 597484
rect 295750 596325 295810 600339
rect 295747 596324 295813 596325
rect 295747 596260 295748 596324
rect 295812 596260 295813 596324
rect 295747 596259 295813 596260
rect 295011 586532 295077 586533
rect 295011 586468 295012 586532
rect 295076 586468 295077 586532
rect 295011 586467 295077 586468
rect 294827 569940 294893 569941
rect 294827 569876 294828 569940
rect 294892 569876 294893 569940
rect 294827 569875 294893 569876
rect 295011 569396 295077 569397
rect 295011 569332 295012 569396
rect 295076 569332 295077 569396
rect 295011 569331 295077 569332
rect 295014 558517 295074 569331
rect 295011 558516 295077 558517
rect 295011 558452 295012 558516
rect 295076 558452 295077 558516
rect 295011 558451 295077 558452
rect 294643 557428 294709 557429
rect 294643 557364 294644 557428
rect 294708 557364 294709 557428
rect 294643 557363 294709 557364
rect 294459 541924 294525 541925
rect 294459 541860 294460 541924
rect 294524 541860 294525 541924
rect 294459 541859 294525 541860
rect 295934 540973 295994 616659
rect 296667 607204 296733 607205
rect 296667 607140 296668 607204
rect 296732 607140 296733 607204
rect 296667 607139 296733 607140
rect 296670 606930 296730 607139
rect 296486 606870 296730 606930
rect 296299 599452 296365 599453
rect 296299 599388 296300 599452
rect 296364 599388 296365 599452
rect 296299 599387 296365 599388
rect 296115 597140 296181 597141
rect 296115 597076 296116 597140
rect 296180 597076 296181 597140
rect 296115 597075 296181 597076
rect 295931 540972 295997 540973
rect 295931 540908 295932 540972
rect 295996 540908 295997 540972
rect 295931 540907 295997 540908
rect 296118 526829 296178 597075
rect 296302 596730 296362 599387
rect 296486 597410 296546 606870
rect 297035 605028 297101 605029
rect 297035 604964 297036 605028
rect 297100 604964 297101 605028
rect 297035 604963 297101 604964
rect 296486 597350 296914 597410
rect 296302 596670 296546 596730
rect 296299 596324 296365 596325
rect 296299 596260 296300 596324
rect 296364 596260 296365 596324
rect 296299 596259 296365 596260
rect 296302 545053 296362 596259
rect 296486 550629 296546 596670
rect 296854 596322 296914 597350
rect 296670 596262 296914 596322
rect 296670 596189 296730 596262
rect 296667 596188 296733 596189
rect 296667 596124 296668 596188
rect 296732 596124 296733 596188
rect 296667 596123 296733 596124
rect 297038 586530 297098 604963
rect 296854 586470 297098 586530
rect 297234 586894 297854 622338
rect 376674 630334 377294 665778
rect 380394 709638 381014 711590
rect 380394 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 381014 709638
rect 380394 709318 381014 709402
rect 380394 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 381014 709318
rect 380394 670054 381014 709082
rect 380394 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 381014 670054
rect 380394 669734 381014 669818
rect 380394 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 381014 669734
rect 377627 648276 377693 648277
rect 377627 648212 377628 648276
rect 377692 648212 377693 648276
rect 377627 648211 377693 648212
rect 376674 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 377294 630334
rect 376674 630014 377294 630098
rect 376674 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 377294 630014
rect 298139 619988 298205 619989
rect 298139 619924 298140 619988
rect 298204 619924 298205 619988
rect 298139 619923 298205 619924
rect 298142 601901 298202 619923
rect 319568 619174 319888 619206
rect 319568 618938 319610 619174
rect 319846 618938 319888 619174
rect 319568 618854 319888 618938
rect 319568 618618 319610 618854
rect 319846 618618 319888 618854
rect 319568 618586 319888 618618
rect 350288 619174 350608 619206
rect 350288 618938 350330 619174
rect 350566 618938 350608 619174
rect 350288 618854 350608 618938
rect 350288 618618 350330 618854
rect 350566 618618 350608 618854
rect 350288 618586 350608 618618
rect 304208 615454 304528 615486
rect 304208 615218 304250 615454
rect 304486 615218 304528 615454
rect 304208 615134 304528 615218
rect 304208 614898 304250 615134
rect 304486 614898 304528 615134
rect 304208 614866 304528 614898
rect 334928 615454 335248 615486
rect 334928 615218 334970 615454
rect 335206 615218 335248 615454
rect 334928 615134 335248 615218
rect 334928 614898 334970 615134
rect 335206 614898 335248 615134
rect 334928 614866 335248 614898
rect 365648 615454 365968 615486
rect 365648 615218 365690 615454
rect 365926 615218 365968 615454
rect 365648 615134 365968 615218
rect 365648 614898 365690 615134
rect 365926 614898 365968 615134
rect 365648 614866 365968 614898
rect 298323 610196 298389 610197
rect 298323 610132 298324 610196
rect 298388 610132 298389 610196
rect 298323 610131 298389 610132
rect 298139 601900 298205 601901
rect 298139 601836 298140 601900
rect 298204 601836 298205 601900
rect 298139 601835 298205 601836
rect 298326 594829 298386 610131
rect 299611 607748 299677 607749
rect 299611 607684 299612 607748
rect 299676 607684 299677 607748
rect 299611 607683 299677 607684
rect 298507 606932 298573 606933
rect 298507 606868 298508 606932
rect 298572 606868 298573 606932
rect 298507 606867 298573 606868
rect 298323 594828 298389 594829
rect 298323 594764 298324 594828
rect 298388 594764 298389 594828
rect 298323 594763 298389 594764
rect 298510 592109 298570 606867
rect 299427 605300 299493 605301
rect 299427 605236 299428 605300
rect 299492 605236 299493 605300
rect 299427 605235 299493 605236
rect 299243 604484 299309 604485
rect 299243 604420 299244 604484
rect 299308 604420 299309 604484
rect 299243 604419 299309 604420
rect 298691 602988 298757 602989
rect 298691 602924 298692 602988
rect 298756 602924 298757 602988
rect 298691 602923 298757 602924
rect 298507 592108 298573 592109
rect 298507 592044 298508 592108
rect 298572 592044 298573 592108
rect 298507 592043 298573 592044
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 296667 577420 296733 577421
rect 296667 577356 296668 577420
rect 296732 577356 296733 577420
rect 296667 577355 296733 577356
rect 296670 576741 296730 577355
rect 296667 576740 296733 576741
rect 296667 576676 296668 576740
rect 296732 576676 296733 576740
rect 296667 576675 296733 576676
rect 296667 567492 296733 567493
rect 296667 567428 296668 567492
rect 296732 567428 296733 567492
rect 296667 567427 296733 567428
rect 296670 567085 296730 567427
rect 296667 567084 296733 567085
rect 296667 567020 296668 567084
rect 296732 567020 296733 567084
rect 296667 567019 296733 567020
rect 296667 557836 296733 557837
rect 296667 557772 296668 557836
rect 296732 557772 296733 557836
rect 296667 557771 296733 557772
rect 296670 557293 296730 557771
rect 296667 557292 296733 557293
rect 296667 557228 296668 557292
rect 296732 557228 296733 557292
rect 296667 557227 296733 557228
rect 296483 550628 296549 550629
rect 296483 550564 296484 550628
rect 296548 550564 296549 550628
rect 296483 550563 296549 550564
rect 296483 550220 296549 550221
rect 296483 550156 296484 550220
rect 296548 550156 296549 550220
rect 296483 550155 296549 550156
rect 296299 545052 296365 545053
rect 296299 544988 296300 545052
rect 296364 544988 296365 545052
rect 296299 544987 296365 544988
rect 296486 543690 296546 550155
rect 296302 543630 296546 543690
rect 296302 542333 296362 543630
rect 296667 542468 296733 542469
rect 296667 542404 296668 542468
rect 296732 542404 296733 542468
rect 296667 542403 296733 542404
rect 296299 542332 296365 542333
rect 296299 542268 296300 542332
rect 296364 542268 296365 542332
rect 296670 542330 296730 542403
rect 296299 542267 296365 542268
rect 296486 542270 296730 542330
rect 296115 526828 296181 526829
rect 296115 526764 296116 526828
rect 296180 526764 296181 526828
rect 296115 526763 296181 526764
rect 296486 524381 296546 542270
rect 296854 531861 296914 586470
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 296851 531860 296917 531861
rect 296851 531796 296852 531860
rect 296916 531796 296917 531860
rect 296851 531795 296917 531796
rect 296483 524380 296549 524381
rect 296483 524316 296484 524380
rect 296548 524316 296549 524380
rect 296483 524315 296549 524316
rect 297234 522121 297854 550338
rect 298694 536621 298754 602923
rect 299059 595508 299125 595509
rect 299059 595444 299060 595508
rect 299124 595444 299125 595508
rect 299059 595443 299125 595444
rect 298875 592924 298941 592925
rect 298875 592860 298876 592924
rect 298940 592860 298941 592924
rect 298875 592859 298941 592860
rect 298878 550085 298938 592859
rect 299062 557293 299122 595443
rect 299246 571165 299306 604419
rect 299430 602989 299490 605235
rect 299614 604485 299674 607683
rect 299611 604484 299677 604485
rect 299611 604420 299612 604484
rect 299676 604420 299677 604484
rect 299611 604419 299677 604420
rect 299427 602988 299493 602989
rect 299427 602924 299428 602988
rect 299492 602924 299493 602988
rect 299427 602923 299493 602924
rect 299427 602036 299493 602037
rect 299427 601972 299428 602036
rect 299492 601972 299493 602036
rect 299427 601971 299493 601972
rect 299430 597549 299490 601971
rect 299427 597548 299493 597549
rect 299427 597484 299428 597548
rect 299492 597484 299493 597548
rect 299427 597483 299493 597484
rect 299795 596460 299861 596461
rect 299795 596396 299796 596460
rect 299860 596396 299861 596460
rect 299795 596395 299861 596396
rect 299243 571164 299309 571165
rect 299243 571100 299244 571164
rect 299308 571100 299309 571164
rect 299243 571099 299309 571100
rect 299243 570076 299309 570077
rect 299243 570012 299244 570076
rect 299308 570012 299309 570076
rect 299243 570011 299309 570012
rect 299059 557292 299125 557293
rect 299059 557228 299060 557292
rect 299124 557228 299125 557292
rect 299059 557227 299125 557228
rect 298875 550084 298941 550085
rect 298875 550020 298876 550084
rect 298940 550020 298941 550084
rect 298875 550019 298941 550020
rect 298691 536620 298757 536621
rect 298691 536556 298692 536620
rect 298756 536556 298757 536620
rect 298691 536555 298757 536556
rect 299246 536485 299306 570011
rect 299243 536484 299309 536485
rect 299243 536420 299244 536484
rect 299308 536420 299309 536484
rect 299243 536419 299309 536420
rect 299798 521389 299858 596395
rect 376674 594334 377294 629778
rect 377630 626517 377690 648211
rect 377811 635900 377877 635901
rect 377811 635836 377812 635900
rect 377876 635836 377877 635900
rect 377811 635835 377877 635836
rect 377627 626516 377693 626517
rect 377627 626452 377628 626516
rect 377692 626452 377693 626516
rect 377627 626451 377693 626452
rect 377814 615093 377874 635835
rect 380394 634054 381014 669498
rect 380394 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 381014 634054
rect 380394 633734 381014 633818
rect 380394 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 381014 633734
rect 377811 615092 377877 615093
rect 377811 615028 377812 615092
rect 377876 615028 377877 615092
rect 377811 615027 377877 615028
rect 376674 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 377294 594334
rect 376674 594014 377294 594098
rect 376674 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 377294 594014
rect 319568 583174 319888 583206
rect 319568 582938 319610 583174
rect 319846 582938 319888 583174
rect 319568 582854 319888 582938
rect 319568 582618 319610 582854
rect 319846 582618 319888 582854
rect 319568 582586 319888 582618
rect 350288 583174 350608 583206
rect 350288 582938 350330 583174
rect 350566 582938 350608 583174
rect 350288 582854 350608 582938
rect 350288 582618 350330 582854
rect 350566 582618 350608 582854
rect 350288 582586 350608 582618
rect 304208 579454 304528 579486
rect 304208 579218 304250 579454
rect 304486 579218 304528 579454
rect 304208 579134 304528 579218
rect 304208 578898 304250 579134
rect 304486 578898 304528 579134
rect 304208 578866 304528 578898
rect 334928 579454 335248 579486
rect 334928 579218 334970 579454
rect 335206 579218 335248 579454
rect 334928 579134 335248 579218
rect 334928 578898 334970 579134
rect 335206 578898 335248 579134
rect 334928 578866 335248 578898
rect 365648 579454 365968 579486
rect 365648 579218 365690 579454
rect 365926 579218 365968 579454
rect 365648 579134 365968 579218
rect 365648 578898 365690 579134
rect 365926 578898 365968 579134
rect 365648 578866 365968 578898
rect 304674 558334 305294 558575
rect 304674 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 305294 558334
rect 304674 558014 305294 558098
rect 304674 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 305294 558014
rect 304674 522121 305294 557778
rect 340674 558334 341294 558575
rect 340674 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 341294 558334
rect 340674 558014 341294 558098
rect 340674 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 341294 558014
rect 340674 522121 341294 557778
rect 376674 558334 377294 593778
rect 380394 598054 381014 633498
rect 380394 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 381014 598054
rect 380394 597734 381014 597818
rect 380394 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 381014 597734
rect 379467 577556 379533 577557
rect 379467 577492 379468 577556
rect 379532 577492 379533 577556
rect 379467 577491 379533 577492
rect 376674 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 377294 558334
rect 376674 558014 377294 558098
rect 376674 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 377294 558014
rect 376674 522121 377294 557778
rect 379470 537437 379530 577491
rect 380394 562054 381014 597498
rect 384114 710598 384734 711590
rect 384114 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 384734 710598
rect 384114 710278 384734 710362
rect 384114 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 384734 710278
rect 384114 673774 384734 710042
rect 384114 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 384734 673774
rect 384114 673454 384734 673538
rect 384114 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 384734 673454
rect 384114 637774 384734 673218
rect 384114 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 384734 637774
rect 384114 637454 384734 637538
rect 384114 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 384734 637454
rect 384114 601774 384734 637218
rect 384114 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 384734 601774
rect 384114 601454 384734 601538
rect 384114 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 384734 601454
rect 382227 574292 382293 574293
rect 382227 574228 382228 574292
rect 382292 574228 382293 574292
rect 382227 574227 382293 574228
rect 380394 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 381014 562054
rect 380394 561734 381014 561818
rect 380394 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 381014 561734
rect 379467 537436 379533 537437
rect 379467 537372 379468 537436
rect 379532 537372 379533 537436
rect 379467 537371 379533 537372
rect 380394 526054 381014 561498
rect 382230 545733 382290 574227
rect 384114 565774 384734 601218
rect 384114 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 384734 565774
rect 384114 565454 384734 565538
rect 384114 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 384734 565454
rect 382227 545732 382293 545733
rect 382227 545668 382228 545732
rect 382292 545668 382293 545732
rect 382227 545667 382293 545668
rect 380394 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 381014 526054
rect 380394 525734 381014 525818
rect 380394 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 381014 525734
rect 380394 522121 381014 525498
rect 384114 529774 384734 565218
rect 384114 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 384734 529774
rect 384114 529454 384734 529538
rect 384114 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 384734 529454
rect 384114 522121 384734 529218
rect 387834 711558 388454 711590
rect 387834 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 388454 711558
rect 387834 711238 388454 711322
rect 387834 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 388454 711238
rect 387834 677494 388454 711002
rect 387834 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 388454 677494
rect 387834 677174 388454 677258
rect 387834 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 388454 677174
rect 387834 641494 388454 676938
rect 387834 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 388454 641494
rect 387834 641174 388454 641258
rect 387834 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 388454 641174
rect 387834 605494 388454 640938
rect 387834 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 388454 605494
rect 387834 605174 388454 605258
rect 387834 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 388454 605174
rect 387834 569494 388454 604938
rect 387834 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 388454 569494
rect 387834 569174 388454 569258
rect 387834 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 388454 569174
rect 387834 533494 388454 568938
rect 387834 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 388454 533494
rect 387834 533174 388454 533258
rect 387834 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 388454 533174
rect 387834 522121 388454 532938
rect 397794 704838 398414 711590
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 522121 398414 542898
rect 401514 705798 402134 711590
rect 401514 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 402134 705798
rect 401514 705478 402134 705562
rect 401514 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 402134 705478
rect 401514 691174 402134 705242
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 522121 402134 546618
rect 405234 706758 405854 711590
rect 405234 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 405854 706758
rect 405234 706438 405854 706522
rect 405234 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 405854 706438
rect 405234 694894 405854 706202
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 522121 405854 550338
rect 408954 707718 409574 711590
rect 408954 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 409574 707718
rect 408954 707398 409574 707482
rect 408954 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 409574 707398
rect 408954 698614 409574 707162
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 522121 409574 554058
rect 412674 708678 413294 711590
rect 412674 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 413294 708678
rect 412674 708358 413294 708442
rect 412674 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 413294 708358
rect 412674 666334 413294 708122
rect 412674 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 413294 666334
rect 412674 666014 413294 666098
rect 412674 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 413294 666014
rect 412674 630334 413294 665778
rect 412674 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 413294 630334
rect 412674 630014 413294 630098
rect 412674 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 413294 630014
rect 412674 594334 413294 629778
rect 412674 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 413294 594334
rect 412674 594014 413294 594098
rect 412674 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 413294 594014
rect 412674 558334 413294 593778
rect 412674 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 413294 558334
rect 412674 558014 413294 558098
rect 412674 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 413294 558014
rect 412674 522121 413294 557778
rect 416394 709638 417014 711590
rect 416394 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 417014 709638
rect 416394 709318 417014 709402
rect 416394 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 417014 709318
rect 416394 670054 417014 709082
rect 416394 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 417014 670054
rect 416394 669734 417014 669818
rect 416394 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 417014 669734
rect 416394 634054 417014 669498
rect 416394 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 417014 634054
rect 416394 633734 417014 633818
rect 416394 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 417014 633734
rect 416394 598054 417014 633498
rect 416394 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 417014 598054
rect 416394 597734 417014 597818
rect 416394 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 417014 597734
rect 416394 562054 417014 597498
rect 416394 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 417014 562054
rect 416394 561734 417014 561818
rect 416394 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 417014 561734
rect 416394 526054 417014 561498
rect 416394 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 417014 526054
rect 416394 525734 417014 525818
rect 416394 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 417014 525734
rect 416394 522121 417014 525498
rect 420114 710598 420734 711590
rect 420114 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 420734 710598
rect 420114 710278 420734 710362
rect 420114 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 420734 710278
rect 420114 673774 420734 710042
rect 420114 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 420734 673774
rect 420114 673454 420734 673538
rect 420114 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 420734 673454
rect 420114 637774 420734 673218
rect 420114 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 420734 637774
rect 420114 637454 420734 637538
rect 420114 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 420734 637454
rect 420114 601774 420734 637218
rect 420114 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 420734 601774
rect 420114 601454 420734 601538
rect 420114 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 420734 601454
rect 420114 565774 420734 601218
rect 420114 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 420734 565774
rect 420114 565454 420734 565538
rect 420114 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 420734 565454
rect 420114 529774 420734 565218
rect 420114 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 420734 529774
rect 420114 529454 420734 529538
rect 420114 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 420734 529454
rect 420114 522121 420734 529218
rect 423834 711558 424454 711590
rect 423834 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 424454 711558
rect 423834 711238 424454 711322
rect 423834 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 424454 711238
rect 423834 677494 424454 711002
rect 423834 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 424454 677494
rect 423834 677174 424454 677258
rect 423834 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 424454 677174
rect 423834 641494 424454 676938
rect 423834 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 424454 641494
rect 423834 641174 424454 641258
rect 423834 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 424454 641174
rect 423834 605494 424454 640938
rect 423834 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 424454 605494
rect 423834 605174 424454 605258
rect 423834 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 424454 605174
rect 423834 569494 424454 604938
rect 423834 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 424454 569494
rect 423834 569174 424454 569258
rect 423834 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 424454 569174
rect 423834 533494 424454 568938
rect 423834 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 424454 533494
rect 423834 533174 424454 533258
rect 423834 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 424454 533174
rect 423834 522121 424454 532938
rect 433794 704838 434414 711590
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 522121 434414 542898
rect 437514 705798 438134 711590
rect 437514 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 438134 705798
rect 437514 705478 438134 705562
rect 437514 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 438134 705478
rect 437514 691174 438134 705242
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 522121 438134 546618
rect 441234 706758 441854 711590
rect 441234 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 441854 706758
rect 441234 706438 441854 706522
rect 441234 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 441854 706438
rect 441234 694894 441854 706202
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 522121 441854 550338
rect 444954 707718 445574 711590
rect 444954 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 445574 707718
rect 444954 707398 445574 707482
rect 444954 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 445574 707398
rect 444954 698614 445574 707162
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 522121 445574 554058
rect 448674 708678 449294 711590
rect 448674 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 449294 708678
rect 448674 708358 449294 708442
rect 448674 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 449294 708358
rect 448674 666334 449294 708122
rect 448674 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 449294 666334
rect 448674 666014 449294 666098
rect 448674 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 449294 666014
rect 448674 630334 449294 665778
rect 452394 709638 453014 711590
rect 452394 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 453014 709638
rect 452394 709318 453014 709402
rect 452394 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 453014 709318
rect 452394 670054 453014 709082
rect 452394 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 453014 670054
rect 452394 669734 453014 669818
rect 452394 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 453014 669734
rect 450491 655076 450557 655077
rect 450491 655012 450492 655076
rect 450556 655012 450557 655076
rect 450491 655011 450557 655012
rect 448674 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 449294 630334
rect 448674 630014 449294 630098
rect 448674 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 449294 630014
rect 448674 594334 449294 629778
rect 448674 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 449294 594334
rect 448674 594014 449294 594098
rect 448674 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 449294 594014
rect 448674 558334 449294 593778
rect 448674 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 449294 558334
rect 448674 558014 449294 558098
rect 448674 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 449294 558014
rect 448674 522121 449294 557778
rect 450494 529141 450554 655011
rect 452394 634054 453014 669498
rect 452394 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 453014 634054
rect 452394 633734 453014 633818
rect 452394 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 453014 633734
rect 452394 598054 453014 633498
rect 452394 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 453014 598054
rect 452394 597734 453014 597818
rect 452394 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 453014 597734
rect 452394 562054 453014 597498
rect 452394 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 453014 562054
rect 452394 561734 453014 561818
rect 452394 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 453014 561734
rect 450491 529140 450557 529141
rect 450491 529076 450492 529140
rect 450556 529076 450557 529140
rect 450491 529075 450557 529076
rect 452394 526054 453014 561498
rect 452394 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 453014 526054
rect 452394 525734 453014 525818
rect 452394 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 453014 525734
rect 452394 522121 453014 525498
rect 456114 710598 456734 711590
rect 456114 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 456734 710598
rect 456114 710278 456734 710362
rect 456114 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 456734 710278
rect 456114 673774 456734 710042
rect 456114 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 456734 673774
rect 456114 673454 456734 673538
rect 456114 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 456734 673454
rect 456114 637774 456734 673218
rect 456114 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 456734 637774
rect 456114 637454 456734 637538
rect 456114 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 456734 637454
rect 456114 601774 456734 637218
rect 456114 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 456734 601774
rect 456114 601454 456734 601538
rect 456114 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 456734 601454
rect 456114 565774 456734 601218
rect 456114 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 456734 565774
rect 456114 565454 456734 565538
rect 456114 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 456734 565454
rect 456114 529774 456734 565218
rect 456114 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 456734 529774
rect 456114 529454 456734 529538
rect 456114 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 456734 529454
rect 456114 522121 456734 529218
rect 459834 711558 460454 711590
rect 459834 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 460454 711558
rect 459834 711238 460454 711322
rect 459834 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 460454 711238
rect 459834 677494 460454 711002
rect 459834 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 460454 677494
rect 459834 677174 460454 677258
rect 459834 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 460454 677174
rect 459834 641494 460454 676938
rect 459834 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 460454 641494
rect 459834 641174 460454 641258
rect 459834 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 460454 641174
rect 459834 605494 460454 640938
rect 459834 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 460454 605494
rect 459834 605174 460454 605258
rect 459834 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 460454 605174
rect 459834 569494 460454 604938
rect 459834 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 460454 569494
rect 459834 569174 460454 569258
rect 459834 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 460454 569174
rect 459834 533494 460454 568938
rect 459834 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 460454 533494
rect 459834 533174 460454 533258
rect 459834 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 460454 533174
rect 459834 522121 460454 532938
rect 469794 704838 470414 711590
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 522121 470414 542898
rect 473514 705798 474134 711590
rect 473514 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 474134 705798
rect 473514 705478 474134 705562
rect 473514 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 474134 705478
rect 473514 691174 474134 705242
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 477234 706758 477854 711590
rect 477234 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 477854 706758
rect 477234 706438 477854 706522
rect 477234 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 477854 706438
rect 477234 694894 477854 706202
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 476619 650044 476685 650045
rect 476619 649980 476620 650044
rect 476684 649980 476685 650044
rect 476619 649979 476685 649980
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 522121 474134 546618
rect 476622 528053 476682 649979
rect 477234 622894 477854 658338
rect 480954 707718 481574 711590
rect 480954 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 481574 707718
rect 480954 707398 481574 707482
rect 480954 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 481574 707398
rect 480954 698614 481574 707162
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480299 653172 480365 653173
rect 480299 653108 480300 653172
rect 480364 653108 480365 653172
rect 480299 653107 480365 653108
rect 479379 641204 479445 641205
rect 479379 641140 479380 641204
rect 479444 641140 479445 641204
rect 479379 641139 479445 641140
rect 478091 639436 478157 639437
rect 478091 639372 478092 639436
rect 478156 639372 478157 639436
rect 478091 639371 478157 639372
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 476619 528052 476685 528053
rect 476619 527988 476620 528052
rect 476684 527988 476685 528052
rect 476619 527987 476685 527988
rect 477234 522121 477854 550338
rect 478094 522749 478154 639371
rect 478091 522748 478157 522749
rect 478091 522684 478092 522748
rect 478156 522684 478157 522748
rect 478091 522683 478157 522684
rect 479382 522613 479442 641139
rect 480302 524381 480362 653107
rect 480954 626614 481574 662058
rect 484674 708678 485294 711590
rect 484674 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 485294 708678
rect 484674 708358 485294 708442
rect 484674 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 485294 708358
rect 484674 666334 485294 708122
rect 484674 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 485294 666334
rect 484674 666014 485294 666098
rect 484674 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 485294 666014
rect 482139 638076 482205 638077
rect 482139 638012 482140 638076
rect 482204 638012 482205 638076
rect 482139 638011 482205 638012
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480299 524380 480365 524381
rect 480299 524316 480300 524380
rect 480364 524316 480365 524380
rect 480299 524315 480365 524316
rect 479379 522612 479445 522613
rect 479379 522548 479380 522612
rect 479444 522548 479445 522612
rect 479379 522547 479445 522548
rect 480954 522121 481574 554058
rect 482142 522885 482202 638011
rect 483611 637940 483677 637941
rect 483611 637876 483612 637940
rect 483676 637876 483677 637940
rect 483611 637875 483677 637876
rect 483614 523021 483674 637875
rect 484674 630334 485294 665778
rect 484674 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 485294 630334
rect 484674 630014 485294 630098
rect 484674 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 485294 630014
rect 484674 594334 485294 629778
rect 484674 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 485294 594334
rect 484674 594014 485294 594098
rect 484674 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 485294 594014
rect 484674 558334 485294 593778
rect 484674 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 485294 558334
rect 484674 558014 485294 558098
rect 484674 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 485294 558014
rect 483611 523020 483677 523021
rect 483611 522956 483612 523020
rect 483676 522956 483677 523020
rect 483611 522955 483677 522956
rect 482139 522884 482205 522885
rect 482139 522820 482140 522884
rect 482204 522820 482205 522884
rect 482139 522819 482205 522820
rect 484674 522121 485294 557778
rect 488394 709638 489014 711590
rect 488394 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 489014 709638
rect 488394 709318 489014 709402
rect 488394 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 489014 709318
rect 488394 670054 489014 709082
rect 488394 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 489014 670054
rect 488394 669734 489014 669818
rect 488394 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 489014 669734
rect 488394 634054 489014 669498
rect 488394 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 489014 634054
rect 488394 633734 489014 633818
rect 488394 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 489014 633734
rect 488394 598054 489014 633498
rect 488394 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 489014 598054
rect 488394 597734 489014 597818
rect 488394 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 489014 597734
rect 488394 562054 489014 597498
rect 488394 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 489014 562054
rect 488394 561734 489014 561818
rect 488394 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 489014 561734
rect 488394 526054 489014 561498
rect 488394 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 489014 526054
rect 488394 525734 489014 525818
rect 488394 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 489014 525734
rect 488394 522121 489014 525498
rect 492114 710598 492734 711590
rect 492114 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 492734 710598
rect 492114 710278 492734 710362
rect 492114 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 492734 710278
rect 492114 673774 492734 710042
rect 492114 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 492734 673774
rect 492114 673454 492734 673538
rect 492114 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 492734 673454
rect 492114 637774 492734 673218
rect 495834 711558 496454 711590
rect 495834 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 496454 711558
rect 495834 711238 496454 711322
rect 495834 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 496454 711238
rect 495834 677494 496454 711002
rect 495834 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 496454 677494
rect 495834 677174 496454 677258
rect 495834 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 496454 677174
rect 495834 654737 496454 676938
rect 505794 704838 506414 711590
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 654737 506414 686898
rect 509514 705798 510134 711590
rect 509514 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 510134 705798
rect 509514 705478 510134 705562
rect 509514 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 510134 705478
rect 509514 691174 510134 705242
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 654956 510134 690618
rect 513234 706758 513854 711590
rect 513234 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 513854 706758
rect 513234 706438 513854 706522
rect 513234 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 513854 706438
rect 513234 694894 513854 706202
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 654737 513854 658338
rect 516954 707718 517574 711590
rect 516954 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 517574 707718
rect 516954 707398 517574 707482
rect 516954 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 517574 707398
rect 516954 698614 517574 707162
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 654737 517574 662058
rect 520674 708678 521294 711590
rect 520674 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 521294 708678
rect 520674 708358 521294 708442
rect 520674 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 521294 708358
rect 520674 666334 521294 708122
rect 520674 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 521294 666334
rect 520674 666014 521294 666098
rect 520674 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 521294 666014
rect 520674 654737 521294 665778
rect 524394 709638 525014 711590
rect 524394 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 525014 709638
rect 524394 709318 525014 709402
rect 524394 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 525014 709318
rect 524394 670054 525014 709082
rect 524394 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 525014 670054
rect 524394 669734 525014 669818
rect 524394 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 525014 669734
rect 524394 654956 525014 669498
rect 528114 710598 528734 711590
rect 528114 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 528734 710598
rect 528114 710278 528734 710362
rect 528114 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 528734 710278
rect 528114 673774 528734 710042
rect 528114 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 528734 673774
rect 528114 673454 528734 673538
rect 528114 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 528734 673454
rect 528114 654737 528734 673218
rect 531834 711558 532454 711590
rect 531834 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 532454 711558
rect 531834 711238 532454 711322
rect 531834 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 532454 711238
rect 531834 677494 532454 711002
rect 531834 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 532454 677494
rect 531834 677174 532454 677258
rect 531834 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 532454 677174
rect 531834 654737 532454 676938
rect 541794 704838 542414 711590
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 494208 651454 494528 651486
rect 494208 651218 494250 651454
rect 494486 651218 494528 651454
rect 494208 651134 494528 651218
rect 494208 650898 494250 651134
rect 494486 650898 494528 651134
rect 494208 650866 494528 650898
rect 524928 651454 525248 651486
rect 524928 651218 524970 651454
rect 525206 651218 525248 651454
rect 524928 651134 525248 651218
rect 524928 650898 524970 651134
rect 525206 650898 525248 651134
rect 524928 650866 525248 650898
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 492114 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 492734 637774
rect 492114 637454 492734 637538
rect 492114 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 492734 637454
rect 492114 601774 492734 637218
rect 509568 619174 509888 619206
rect 509568 618938 509610 619174
rect 509846 618938 509888 619174
rect 509568 618854 509888 618938
rect 509568 618618 509610 618854
rect 509846 618618 509888 618854
rect 509568 618586 509888 618618
rect 494208 615454 494528 615486
rect 494208 615218 494250 615454
rect 494486 615218 494528 615454
rect 494208 615134 494528 615218
rect 494208 614898 494250 615134
rect 494486 614898 494528 615134
rect 494208 614866 494528 614898
rect 524928 615454 525248 615486
rect 524928 615218 524970 615454
rect 525206 615218 525248 615454
rect 524928 615134 525248 615218
rect 524928 614898 524970 615134
rect 525206 614898 525248 615134
rect 524928 614866 525248 614898
rect 541794 615454 542414 650898
rect 545514 705798 546134 711590
rect 545514 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 546134 705798
rect 545514 705478 546134 705562
rect 545514 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 546134 705478
rect 545514 691174 546134 705242
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 543779 621348 543845 621349
rect 543779 621284 543780 621348
rect 543844 621284 543845 621348
rect 543779 621283 543845 621284
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541019 614548 541085 614549
rect 541019 614484 541020 614548
rect 541084 614484 541085 614548
rect 541019 614483 541085 614484
rect 539363 605028 539429 605029
rect 539363 604964 539364 605028
rect 539428 604964 539429 605028
rect 539363 604963 539429 604964
rect 492114 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 492734 601774
rect 538259 601764 538325 601765
rect 538259 601700 538260 601764
rect 538324 601700 538325 601764
rect 538259 601699 538325 601700
rect 492114 601454 492734 601538
rect 492114 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 492734 601454
rect 492114 565774 492734 601218
rect 492114 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 492734 565774
rect 492114 565454 492734 565538
rect 492114 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 492734 565454
rect 492114 529774 492734 565218
rect 492114 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 492734 529774
rect 492114 529454 492734 529538
rect 492114 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 492734 529454
rect 492114 522121 492734 529218
rect 495834 569494 496454 600207
rect 500171 599724 500237 599725
rect 500171 599660 500172 599724
rect 500236 599660 500237 599724
rect 500171 599659 500237 599660
rect 495834 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 496454 569494
rect 495834 569174 496454 569258
rect 495834 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 496454 569174
rect 495834 533494 496454 568938
rect 499067 557428 499133 557429
rect 499067 557364 499068 557428
rect 499132 557364 499133 557428
rect 499067 557363 499133 557364
rect 498699 547636 498765 547637
rect 498699 547572 498700 547636
rect 498764 547572 498765 547636
rect 498699 547571 498765 547572
rect 497411 546140 497477 546141
rect 497411 546076 497412 546140
rect 497476 546076 497477 546140
rect 497411 546075 497477 546076
rect 495834 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 496454 533494
rect 495834 533174 496454 533258
rect 495834 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 496454 533174
rect 495834 522121 496454 532938
rect 299795 521388 299861 521389
rect 299795 521324 299796 521388
rect 299860 521324 299861 521388
rect 299795 521323 299861 521324
rect 291883 520436 291949 520437
rect 291883 520372 291884 520436
rect 291948 520372 291949 520436
rect 291883 520371 291949 520372
rect 497414 520301 497474 546075
rect 497595 529548 497661 529549
rect 497595 529484 497596 529548
rect 497660 529484 497661 529548
rect 497595 529483 497661 529484
rect 497598 520845 497658 529483
rect 498702 521661 498762 547571
rect 498883 533764 498949 533765
rect 498883 533700 498884 533764
rect 498948 533700 498949 533764
rect 498883 533699 498949 533700
rect 498699 521660 498765 521661
rect 498699 521596 498700 521660
rect 498764 521596 498765 521660
rect 498699 521595 498765 521596
rect 497595 520844 497661 520845
rect 497595 520780 497596 520844
rect 497660 520780 497661 520844
rect 497595 520779 497661 520780
rect 498886 520570 498946 533699
rect 499070 524430 499130 557363
rect 499619 534172 499685 534173
rect 499619 534108 499620 534172
rect 499684 534108 499685 534172
rect 499619 534107 499685 534108
rect 499435 525604 499501 525605
rect 499435 525540 499436 525604
rect 499500 525540 499501 525604
rect 499435 525539 499501 525540
rect 499070 524370 499314 524430
rect 499254 521797 499314 524370
rect 499251 521796 499317 521797
rect 499251 521732 499252 521796
rect 499316 521732 499317 521796
rect 499251 521731 499317 521732
rect 499438 520709 499498 525539
rect 499435 520708 499501 520709
rect 499435 520644 499436 520708
rect 499500 520644 499501 520708
rect 499435 520643 499501 520644
rect 499435 520572 499501 520573
rect 499435 520570 499436 520572
rect 498886 520510 499436 520570
rect 499435 520508 499436 520510
rect 499500 520508 499501 520572
rect 499435 520507 499501 520508
rect 497411 520300 497477 520301
rect 497411 520236 497412 520300
rect 497476 520236 497477 520300
rect 497411 520235 497477 520236
rect 499435 520164 499501 520165
rect 499435 520100 499436 520164
rect 499500 520100 499501 520164
rect 499435 520099 499501 520100
rect 202448 511174 202768 511206
rect 202448 510938 202490 511174
rect 202726 510938 202768 511174
rect 202448 510854 202768 510938
rect 202448 510618 202490 510854
rect 202726 510618 202768 510854
rect 202448 510586 202768 510618
rect 233168 511174 233488 511206
rect 233168 510938 233210 511174
rect 233446 510938 233488 511174
rect 233168 510854 233488 510938
rect 233168 510618 233210 510854
rect 233446 510618 233488 510854
rect 233168 510586 233488 510618
rect 263888 511174 264208 511206
rect 263888 510938 263930 511174
rect 264166 510938 264208 511174
rect 263888 510854 264208 510938
rect 263888 510618 263930 510854
rect 264166 510618 264208 510854
rect 263888 510586 264208 510618
rect 294608 511174 294928 511206
rect 294608 510938 294650 511174
rect 294886 510938 294928 511174
rect 294608 510854 294928 510938
rect 294608 510618 294650 510854
rect 294886 510618 294928 510854
rect 294608 510586 294928 510618
rect 325328 511174 325648 511206
rect 325328 510938 325370 511174
rect 325606 510938 325648 511174
rect 325328 510854 325648 510938
rect 325328 510618 325370 510854
rect 325606 510618 325648 510854
rect 325328 510586 325648 510618
rect 356048 511174 356368 511206
rect 356048 510938 356090 511174
rect 356326 510938 356368 511174
rect 356048 510854 356368 510938
rect 356048 510618 356090 510854
rect 356326 510618 356368 510854
rect 356048 510586 356368 510618
rect 386768 511174 387088 511206
rect 386768 510938 386810 511174
rect 387046 510938 387088 511174
rect 386768 510854 387088 510938
rect 386768 510618 386810 510854
rect 387046 510618 387088 510854
rect 386768 510586 387088 510618
rect 417488 511174 417808 511206
rect 417488 510938 417530 511174
rect 417766 510938 417808 511174
rect 417488 510854 417808 510938
rect 417488 510618 417530 510854
rect 417766 510618 417808 510854
rect 417488 510586 417808 510618
rect 448208 511174 448528 511206
rect 448208 510938 448250 511174
rect 448486 510938 448528 511174
rect 448208 510854 448528 510938
rect 448208 510618 448250 510854
rect 448486 510618 448528 510854
rect 448208 510586 448528 510618
rect 478928 511174 479248 511206
rect 478928 510938 478970 511174
rect 479206 510938 479248 511174
rect 478928 510854 479248 510938
rect 478928 510618 478970 510854
rect 479206 510618 479248 510854
rect 478928 510586 479248 510618
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 309968 507454 310288 507486
rect 309968 507218 310010 507454
rect 310246 507218 310288 507454
rect 309968 507134 310288 507218
rect 309968 506898 310010 507134
rect 310246 506898 310288 507134
rect 309968 506866 310288 506898
rect 340688 507454 341008 507486
rect 340688 507218 340730 507454
rect 340966 507218 341008 507454
rect 340688 507134 341008 507218
rect 340688 506898 340730 507134
rect 340966 506898 341008 507134
rect 340688 506866 341008 506898
rect 371408 507454 371728 507486
rect 371408 507218 371450 507454
rect 371686 507218 371728 507454
rect 371408 507134 371728 507218
rect 371408 506898 371450 507134
rect 371686 506898 371728 507134
rect 371408 506866 371728 506898
rect 402128 507454 402448 507486
rect 402128 507218 402170 507454
rect 402406 507218 402448 507454
rect 402128 507134 402448 507218
rect 402128 506898 402170 507134
rect 402406 506898 402448 507134
rect 402128 506866 402448 506898
rect 432848 507454 433168 507486
rect 432848 507218 432890 507454
rect 433126 507218 433168 507454
rect 432848 507134 433168 507218
rect 432848 506898 432890 507134
rect 433126 506898 433168 507134
rect 432848 506866 433168 506898
rect 463568 507454 463888 507486
rect 463568 507218 463610 507454
rect 463846 507218 463888 507454
rect 463568 507134 463888 507218
rect 463568 506898 463610 507134
rect 463846 506898 463888 507134
rect 463568 506866 463888 506898
rect 494288 507454 494608 507486
rect 494288 507218 494330 507454
rect 494566 507218 494608 507454
rect 494288 507134 494608 507218
rect 494288 506898 494330 507134
rect 494566 506898 494608 507134
rect 494288 506866 494608 506898
rect 499438 488341 499498 520099
rect 499435 488340 499501 488341
rect 499435 488276 499436 488340
rect 499500 488276 499501 488340
rect 499435 488275 499501 488276
rect 196674 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 197294 486334
rect 196674 486014 197294 486098
rect 196674 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 197294 486014
rect 196674 450334 197294 485778
rect 202448 475174 202768 475206
rect 202448 474938 202490 475174
rect 202726 474938 202768 475174
rect 202448 474854 202768 474938
rect 202448 474618 202490 474854
rect 202726 474618 202768 474854
rect 202448 474586 202768 474618
rect 233168 475174 233488 475206
rect 233168 474938 233210 475174
rect 233446 474938 233488 475174
rect 233168 474854 233488 474938
rect 233168 474618 233210 474854
rect 233446 474618 233488 474854
rect 233168 474586 233488 474618
rect 263888 475174 264208 475206
rect 263888 474938 263930 475174
rect 264166 474938 264208 475174
rect 263888 474854 264208 474938
rect 263888 474618 263930 474854
rect 264166 474618 264208 474854
rect 263888 474586 264208 474618
rect 294608 475174 294928 475206
rect 294608 474938 294650 475174
rect 294886 474938 294928 475174
rect 294608 474854 294928 474938
rect 294608 474618 294650 474854
rect 294886 474618 294928 474854
rect 294608 474586 294928 474618
rect 325328 475174 325648 475206
rect 325328 474938 325370 475174
rect 325606 474938 325648 475174
rect 325328 474854 325648 474938
rect 325328 474618 325370 474854
rect 325606 474618 325648 474854
rect 325328 474586 325648 474618
rect 356048 475174 356368 475206
rect 356048 474938 356090 475174
rect 356326 474938 356368 475174
rect 356048 474854 356368 474938
rect 356048 474618 356090 474854
rect 356326 474618 356368 474854
rect 356048 474586 356368 474618
rect 386768 475174 387088 475206
rect 386768 474938 386810 475174
rect 387046 474938 387088 475174
rect 386768 474854 387088 474938
rect 386768 474618 386810 474854
rect 387046 474618 387088 474854
rect 386768 474586 387088 474618
rect 417488 475174 417808 475206
rect 417488 474938 417530 475174
rect 417766 474938 417808 475174
rect 417488 474854 417808 474938
rect 417488 474618 417530 474854
rect 417766 474618 417808 474854
rect 417488 474586 417808 474618
rect 448208 475174 448528 475206
rect 448208 474938 448250 475174
rect 448486 474938 448528 475174
rect 448208 474854 448528 474938
rect 448208 474618 448250 474854
rect 448486 474618 448528 474854
rect 448208 474586 448528 474618
rect 478928 475174 479248 475206
rect 478928 474938 478970 475174
rect 479206 474938 479248 475174
rect 478928 474854 479248 474938
rect 478928 474618 478970 474854
rect 479206 474618 479248 474854
rect 478928 474586 479248 474618
rect 217808 471454 218128 471486
rect 217808 471218 217850 471454
rect 218086 471218 218128 471454
rect 217808 471134 218128 471218
rect 217808 470898 217850 471134
rect 218086 470898 218128 471134
rect 217808 470866 218128 470898
rect 248528 471454 248848 471486
rect 248528 471218 248570 471454
rect 248806 471218 248848 471454
rect 248528 471134 248848 471218
rect 248528 470898 248570 471134
rect 248806 470898 248848 471134
rect 248528 470866 248848 470898
rect 279248 471454 279568 471486
rect 279248 471218 279290 471454
rect 279526 471218 279568 471454
rect 279248 471134 279568 471218
rect 279248 470898 279290 471134
rect 279526 470898 279568 471134
rect 279248 470866 279568 470898
rect 309968 471454 310288 471486
rect 309968 471218 310010 471454
rect 310246 471218 310288 471454
rect 309968 471134 310288 471218
rect 309968 470898 310010 471134
rect 310246 470898 310288 471134
rect 309968 470866 310288 470898
rect 340688 471454 341008 471486
rect 340688 471218 340730 471454
rect 340966 471218 341008 471454
rect 340688 471134 341008 471218
rect 340688 470898 340730 471134
rect 340966 470898 341008 471134
rect 340688 470866 341008 470898
rect 371408 471454 371728 471486
rect 371408 471218 371450 471454
rect 371686 471218 371728 471454
rect 371408 471134 371728 471218
rect 371408 470898 371450 471134
rect 371686 470898 371728 471134
rect 371408 470866 371728 470898
rect 402128 471454 402448 471486
rect 402128 471218 402170 471454
rect 402406 471218 402448 471454
rect 402128 471134 402448 471218
rect 402128 470898 402170 471134
rect 402406 470898 402448 471134
rect 402128 470866 402448 470898
rect 432848 471454 433168 471486
rect 432848 471218 432890 471454
rect 433126 471218 433168 471454
rect 432848 471134 433168 471218
rect 432848 470898 432890 471134
rect 433126 470898 433168 471134
rect 432848 470866 433168 470898
rect 463568 471454 463888 471486
rect 463568 471218 463610 471454
rect 463846 471218 463888 471454
rect 463568 471134 463888 471218
rect 463568 470898 463610 471134
rect 463846 470898 463888 471134
rect 463568 470866 463888 470898
rect 494288 471454 494608 471486
rect 494288 471218 494330 471454
rect 494566 471218 494608 471454
rect 494288 471134 494608 471218
rect 494288 470898 494330 471134
rect 494566 470898 494608 471134
rect 494288 470866 494608 470898
rect 196674 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 197294 450334
rect 196674 450014 197294 450098
rect 196674 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 197294 450014
rect 196674 414334 197294 449778
rect 202448 439174 202768 439206
rect 202448 438938 202490 439174
rect 202726 438938 202768 439174
rect 202448 438854 202768 438938
rect 202448 438618 202490 438854
rect 202726 438618 202768 438854
rect 202448 438586 202768 438618
rect 233168 439174 233488 439206
rect 233168 438938 233210 439174
rect 233446 438938 233488 439174
rect 233168 438854 233488 438938
rect 233168 438618 233210 438854
rect 233446 438618 233488 438854
rect 233168 438586 233488 438618
rect 263888 439174 264208 439206
rect 263888 438938 263930 439174
rect 264166 438938 264208 439174
rect 263888 438854 264208 438938
rect 263888 438618 263930 438854
rect 264166 438618 264208 438854
rect 263888 438586 264208 438618
rect 294608 439174 294928 439206
rect 294608 438938 294650 439174
rect 294886 438938 294928 439174
rect 294608 438854 294928 438938
rect 294608 438618 294650 438854
rect 294886 438618 294928 438854
rect 294608 438586 294928 438618
rect 325328 439174 325648 439206
rect 325328 438938 325370 439174
rect 325606 438938 325648 439174
rect 325328 438854 325648 438938
rect 325328 438618 325370 438854
rect 325606 438618 325648 438854
rect 325328 438586 325648 438618
rect 356048 439174 356368 439206
rect 356048 438938 356090 439174
rect 356326 438938 356368 439174
rect 356048 438854 356368 438938
rect 356048 438618 356090 438854
rect 356326 438618 356368 438854
rect 356048 438586 356368 438618
rect 386768 439174 387088 439206
rect 386768 438938 386810 439174
rect 387046 438938 387088 439174
rect 386768 438854 387088 438938
rect 386768 438618 386810 438854
rect 387046 438618 387088 438854
rect 386768 438586 387088 438618
rect 417488 439174 417808 439206
rect 417488 438938 417530 439174
rect 417766 438938 417808 439174
rect 417488 438854 417808 438938
rect 417488 438618 417530 438854
rect 417766 438618 417808 438854
rect 417488 438586 417808 438618
rect 448208 439174 448528 439206
rect 448208 438938 448250 439174
rect 448486 438938 448528 439174
rect 448208 438854 448528 438938
rect 448208 438618 448250 438854
rect 448486 438618 448528 438854
rect 448208 438586 448528 438618
rect 478928 439174 479248 439206
rect 478928 438938 478970 439174
rect 479206 438938 479248 439174
rect 478928 438854 479248 438938
rect 478928 438618 478970 438854
rect 479206 438618 479248 438854
rect 478928 438586 479248 438618
rect 217808 435454 218128 435486
rect 217808 435218 217850 435454
rect 218086 435218 218128 435454
rect 217808 435134 218128 435218
rect 217808 434898 217850 435134
rect 218086 434898 218128 435134
rect 217808 434866 218128 434898
rect 248528 435454 248848 435486
rect 248528 435218 248570 435454
rect 248806 435218 248848 435454
rect 248528 435134 248848 435218
rect 248528 434898 248570 435134
rect 248806 434898 248848 435134
rect 248528 434866 248848 434898
rect 279248 435454 279568 435486
rect 279248 435218 279290 435454
rect 279526 435218 279568 435454
rect 279248 435134 279568 435218
rect 279248 434898 279290 435134
rect 279526 434898 279568 435134
rect 279248 434866 279568 434898
rect 309968 435454 310288 435486
rect 309968 435218 310010 435454
rect 310246 435218 310288 435454
rect 309968 435134 310288 435218
rect 309968 434898 310010 435134
rect 310246 434898 310288 435134
rect 309968 434866 310288 434898
rect 340688 435454 341008 435486
rect 340688 435218 340730 435454
rect 340966 435218 341008 435454
rect 340688 435134 341008 435218
rect 340688 434898 340730 435134
rect 340966 434898 341008 435134
rect 340688 434866 341008 434898
rect 371408 435454 371728 435486
rect 371408 435218 371450 435454
rect 371686 435218 371728 435454
rect 371408 435134 371728 435218
rect 371408 434898 371450 435134
rect 371686 434898 371728 435134
rect 371408 434866 371728 434898
rect 402128 435454 402448 435486
rect 402128 435218 402170 435454
rect 402406 435218 402448 435454
rect 402128 435134 402448 435218
rect 402128 434898 402170 435134
rect 402406 434898 402448 435134
rect 402128 434866 402448 434898
rect 432848 435454 433168 435486
rect 432848 435218 432890 435454
rect 433126 435218 433168 435454
rect 432848 435134 433168 435218
rect 432848 434898 432890 435134
rect 433126 434898 433168 435134
rect 432848 434866 433168 434898
rect 463568 435454 463888 435486
rect 463568 435218 463610 435454
rect 463846 435218 463888 435454
rect 463568 435134 463888 435218
rect 463568 434898 463610 435134
rect 463846 434898 463888 435134
rect 463568 434866 463888 434898
rect 494288 435454 494608 435486
rect 494288 435218 494330 435454
rect 494566 435218 494608 435454
rect 494288 435134 494608 435218
rect 494288 434898 494330 435134
rect 494566 434898 494608 435134
rect 494288 434866 494608 434898
rect 196674 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 197294 414334
rect 196674 414014 197294 414098
rect 196674 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 197294 414014
rect 196674 378334 197294 413778
rect 202448 403174 202768 403206
rect 202448 402938 202490 403174
rect 202726 402938 202768 403174
rect 202448 402854 202768 402938
rect 202448 402618 202490 402854
rect 202726 402618 202768 402854
rect 202448 402586 202768 402618
rect 233168 403174 233488 403206
rect 233168 402938 233210 403174
rect 233446 402938 233488 403174
rect 233168 402854 233488 402938
rect 233168 402618 233210 402854
rect 233446 402618 233488 402854
rect 233168 402586 233488 402618
rect 263888 403174 264208 403206
rect 263888 402938 263930 403174
rect 264166 402938 264208 403174
rect 263888 402854 264208 402938
rect 263888 402618 263930 402854
rect 264166 402618 264208 402854
rect 263888 402586 264208 402618
rect 294608 403174 294928 403206
rect 294608 402938 294650 403174
rect 294886 402938 294928 403174
rect 294608 402854 294928 402938
rect 294608 402618 294650 402854
rect 294886 402618 294928 402854
rect 294608 402586 294928 402618
rect 325328 403174 325648 403206
rect 325328 402938 325370 403174
rect 325606 402938 325648 403174
rect 325328 402854 325648 402938
rect 325328 402618 325370 402854
rect 325606 402618 325648 402854
rect 325328 402586 325648 402618
rect 356048 403174 356368 403206
rect 356048 402938 356090 403174
rect 356326 402938 356368 403174
rect 356048 402854 356368 402938
rect 356048 402618 356090 402854
rect 356326 402618 356368 402854
rect 356048 402586 356368 402618
rect 386768 403174 387088 403206
rect 386768 402938 386810 403174
rect 387046 402938 387088 403174
rect 386768 402854 387088 402938
rect 386768 402618 386810 402854
rect 387046 402618 387088 402854
rect 386768 402586 387088 402618
rect 417488 403174 417808 403206
rect 417488 402938 417530 403174
rect 417766 402938 417808 403174
rect 417488 402854 417808 402938
rect 417488 402618 417530 402854
rect 417766 402618 417808 402854
rect 417488 402586 417808 402618
rect 448208 403174 448528 403206
rect 448208 402938 448250 403174
rect 448486 402938 448528 403174
rect 448208 402854 448528 402938
rect 448208 402618 448250 402854
rect 448486 402618 448528 402854
rect 448208 402586 448528 402618
rect 478928 403174 479248 403206
rect 478928 402938 478970 403174
rect 479206 402938 479248 403174
rect 478928 402854 479248 402938
rect 478928 402618 478970 402854
rect 479206 402618 479248 402854
rect 478928 402586 479248 402618
rect 217808 399454 218128 399486
rect 217808 399218 217850 399454
rect 218086 399218 218128 399454
rect 217808 399134 218128 399218
rect 217808 398898 217850 399134
rect 218086 398898 218128 399134
rect 217808 398866 218128 398898
rect 248528 399454 248848 399486
rect 248528 399218 248570 399454
rect 248806 399218 248848 399454
rect 248528 399134 248848 399218
rect 248528 398898 248570 399134
rect 248806 398898 248848 399134
rect 248528 398866 248848 398898
rect 279248 399454 279568 399486
rect 279248 399218 279290 399454
rect 279526 399218 279568 399454
rect 279248 399134 279568 399218
rect 279248 398898 279290 399134
rect 279526 398898 279568 399134
rect 279248 398866 279568 398898
rect 309968 399454 310288 399486
rect 309968 399218 310010 399454
rect 310246 399218 310288 399454
rect 309968 399134 310288 399218
rect 309968 398898 310010 399134
rect 310246 398898 310288 399134
rect 309968 398866 310288 398898
rect 340688 399454 341008 399486
rect 340688 399218 340730 399454
rect 340966 399218 341008 399454
rect 340688 399134 341008 399218
rect 340688 398898 340730 399134
rect 340966 398898 341008 399134
rect 340688 398866 341008 398898
rect 371408 399454 371728 399486
rect 371408 399218 371450 399454
rect 371686 399218 371728 399454
rect 371408 399134 371728 399218
rect 371408 398898 371450 399134
rect 371686 398898 371728 399134
rect 371408 398866 371728 398898
rect 402128 399454 402448 399486
rect 402128 399218 402170 399454
rect 402406 399218 402448 399454
rect 402128 399134 402448 399218
rect 402128 398898 402170 399134
rect 402406 398898 402448 399134
rect 402128 398866 402448 398898
rect 432848 399454 433168 399486
rect 432848 399218 432890 399454
rect 433126 399218 433168 399454
rect 432848 399134 433168 399218
rect 432848 398898 432890 399134
rect 433126 398898 433168 399134
rect 432848 398866 433168 398898
rect 463568 399454 463888 399486
rect 463568 399218 463610 399454
rect 463846 399218 463888 399454
rect 463568 399134 463888 399218
rect 463568 398898 463610 399134
rect 463846 398898 463888 399134
rect 463568 398866 463888 398898
rect 494288 399454 494608 399486
rect 494288 399218 494330 399454
rect 494566 399218 494608 399454
rect 494288 399134 494608 399218
rect 494288 398898 494330 399134
rect 494566 398898 494608 399134
rect 494288 398866 494608 398898
rect 357939 390284 358005 390285
rect 357939 390220 357940 390284
rect 358004 390220 358005 390284
rect 357939 390219 358005 390220
rect 196674 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 197294 378334
rect 196674 378014 197294 378098
rect 196674 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 197294 378014
rect 196674 342334 197294 377778
rect 196674 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 197294 342334
rect 196674 342014 197294 342098
rect 196674 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 197294 342014
rect 196674 306334 197294 341778
rect 196674 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 197294 306334
rect 196674 306014 197294 306098
rect 196674 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 197294 306014
rect 196674 270334 197294 305778
rect 196674 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 197294 270334
rect 196674 270014 197294 270098
rect 196674 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 197294 270014
rect 196674 234334 197294 269778
rect 200394 382054 201014 388711
rect 200394 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 201014 382054
rect 200394 381734 201014 381818
rect 200394 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 201014 381734
rect 200394 346054 201014 381498
rect 200394 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 201014 346054
rect 200394 345734 201014 345818
rect 200394 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 201014 345734
rect 200394 310054 201014 345498
rect 200394 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 201014 310054
rect 200394 309734 201014 309818
rect 200394 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 201014 309734
rect 200394 274054 201014 309498
rect 200394 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 201014 274054
rect 200394 273734 201014 273818
rect 200394 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 201014 273734
rect 197859 245716 197925 245717
rect 197859 245652 197860 245716
rect 197924 245652 197925 245716
rect 197859 245651 197925 245652
rect 196674 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 197294 234334
rect 196674 234014 197294 234098
rect 196674 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 197294 234014
rect 196674 198334 197294 233778
rect 196674 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 197294 198334
rect 196674 198014 197294 198098
rect 196674 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 197294 198014
rect 196674 162334 197294 197778
rect 197862 186965 197922 245651
rect 200394 238054 201014 273498
rect 200394 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 201014 238054
rect 200394 237734 201014 237818
rect 200394 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 201014 237734
rect 200394 202054 201014 237498
rect 200394 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 201014 202054
rect 200394 201734 201014 201818
rect 200394 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 201014 201734
rect 197859 186964 197925 186965
rect 197859 186900 197860 186964
rect 197924 186900 197925 186964
rect 197859 186899 197925 186900
rect 196674 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 197294 162334
rect 196674 162014 197294 162098
rect 196674 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 197294 162014
rect 196674 126334 197294 161778
rect 196674 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 197294 126334
rect 196674 126014 197294 126098
rect 196674 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 197294 126014
rect 196674 90334 197294 125778
rect 196674 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 197294 90334
rect 196674 90014 197294 90098
rect 196674 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 197294 90014
rect 196674 54334 197294 89778
rect 196674 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 197294 54334
rect 196674 54014 197294 54098
rect 196674 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 197294 54014
rect 196674 18334 197294 53778
rect 196674 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 197294 18334
rect 196674 18014 197294 18098
rect 196674 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 197294 18014
rect 196674 -4186 197294 17778
rect 196674 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 197294 -4186
rect 196674 -4506 197294 -4422
rect 196674 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 197294 -4506
rect 196674 -7654 197294 -4742
rect 200394 166054 201014 201498
rect 200394 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 201014 166054
rect 200394 165734 201014 165818
rect 200394 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 201014 165734
rect 200394 130054 201014 165498
rect 200394 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 201014 130054
rect 200394 129734 201014 129818
rect 200394 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 201014 129734
rect 200394 94054 201014 129498
rect 200394 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 201014 94054
rect 200394 93734 201014 93818
rect 200394 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 201014 93734
rect 200394 58054 201014 93498
rect 200394 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 201014 58054
rect 200394 57734 201014 57818
rect 200394 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 201014 57734
rect 200394 22054 201014 57498
rect 200394 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 201014 22054
rect 200394 21734 201014 21818
rect 200394 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 201014 21734
rect 200394 -5146 201014 21498
rect 200394 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 201014 -5146
rect 200394 -5466 201014 -5382
rect 200394 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 201014 -5466
rect 200394 -7654 201014 -5702
rect 204114 385774 204734 388711
rect 204114 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 204734 385774
rect 204114 385454 204734 385538
rect 204114 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 204734 385454
rect 204114 349774 204734 385218
rect 204114 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 204734 349774
rect 204114 349454 204734 349538
rect 204114 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 204734 349454
rect 204114 313774 204734 349218
rect 204114 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 204734 313774
rect 204114 313454 204734 313538
rect 204114 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 204734 313454
rect 204114 277774 204734 313218
rect 204114 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 204734 277774
rect 204114 277454 204734 277538
rect 204114 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 204734 277454
rect 204114 241774 204734 277218
rect 204114 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 204734 241774
rect 204114 241454 204734 241538
rect 204114 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 204734 241454
rect 204114 205774 204734 241218
rect 204114 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 204734 205774
rect 204114 205454 204734 205538
rect 204114 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 204734 205454
rect 204114 169774 204734 205218
rect 204114 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 204734 169774
rect 204114 169454 204734 169538
rect 204114 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 204734 169454
rect 204114 133774 204734 169218
rect 204114 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 204734 133774
rect 204114 133454 204734 133538
rect 204114 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 204734 133454
rect 204114 97774 204734 133218
rect 204114 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 204734 97774
rect 204114 97454 204734 97538
rect 204114 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 204734 97454
rect 204114 61774 204734 97218
rect 204114 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 204734 61774
rect 204114 61454 204734 61538
rect 204114 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 204734 61454
rect 204114 25774 204734 61218
rect 204114 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 204734 25774
rect 204114 25454 204734 25538
rect 204114 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 204734 25454
rect 204114 -6106 204734 25218
rect 204114 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 204734 -6106
rect 204114 -6426 204734 -6342
rect 204114 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 204734 -6426
rect 204114 -7654 204734 -6662
rect 207834 353494 208454 388711
rect 207834 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 208454 353494
rect 207834 353174 208454 353258
rect 207834 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 208454 353174
rect 207834 317494 208454 352938
rect 217794 363454 218414 388711
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 214787 346628 214853 346629
rect 214787 346564 214788 346628
rect 214852 346564 214853 346628
rect 214787 346563 214853 346564
rect 214603 342820 214669 342821
rect 214603 342756 214604 342820
rect 214668 342756 214669 342820
rect 214603 342755 214669 342756
rect 214419 342548 214485 342549
rect 214419 342484 214420 342548
rect 214484 342484 214485 342548
rect 214419 342483 214485 342484
rect 211659 340916 211725 340917
rect 211659 340852 211660 340916
rect 211724 340852 211725 340916
rect 211659 340851 211725 340852
rect 207834 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 208454 317494
rect 207834 317174 208454 317258
rect 207834 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 208454 317174
rect 207834 281494 208454 316938
rect 207834 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 208454 281494
rect 207834 281174 208454 281258
rect 207834 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 208454 281174
rect 207834 245494 208454 280938
rect 211662 265981 211722 340851
rect 211659 265980 211725 265981
rect 211659 265916 211660 265980
rect 211724 265916 211725 265980
rect 211659 265915 211725 265916
rect 207834 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 208454 245494
rect 207834 245174 208454 245258
rect 207834 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 208454 245174
rect 207834 209494 208454 244938
rect 210555 242452 210621 242453
rect 210555 242388 210556 242452
rect 210620 242388 210621 242452
rect 210555 242387 210621 242388
rect 207834 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 208454 209494
rect 207834 209174 208454 209258
rect 207834 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 208454 209174
rect 207834 173494 208454 208938
rect 210558 189685 210618 242387
rect 213131 218652 213197 218653
rect 213131 218588 213132 218652
rect 213196 218588 213197 218652
rect 213131 218587 213197 218588
rect 210555 189684 210621 189685
rect 210555 189620 210556 189684
rect 210620 189620 210621 189684
rect 210555 189619 210621 189620
rect 207834 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 208454 173494
rect 207834 173174 208454 173258
rect 207834 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 208454 173174
rect 207834 137494 208454 172938
rect 213134 167381 213194 218587
rect 214422 179213 214482 342483
rect 214606 180981 214666 342755
rect 214790 306237 214850 346563
rect 217547 345676 217613 345677
rect 217547 345612 217548 345676
rect 217612 345612 217613 345676
rect 217547 345611 217613 345612
rect 217363 344996 217429 344997
rect 217363 344932 217364 344996
rect 217428 344932 217429 344996
rect 217363 344931 217429 344932
rect 215891 340236 215957 340237
rect 215891 340172 215892 340236
rect 215956 340172 215957 340236
rect 215891 340171 215957 340172
rect 214787 306236 214853 306237
rect 214787 306172 214788 306236
rect 214852 306172 214853 306236
rect 214787 306171 214853 306172
rect 215894 264349 215954 340171
rect 217179 339692 217245 339693
rect 217179 339628 217180 339692
rect 217244 339628 217245 339692
rect 217179 339627 217245 339628
rect 216075 338332 216141 338333
rect 216075 338268 216076 338332
rect 216140 338268 216141 338332
rect 216075 338267 216141 338268
rect 215891 264348 215957 264349
rect 215891 264284 215892 264348
rect 215956 264284 215957 264348
rect 215891 264283 215957 264284
rect 216078 262717 216138 338267
rect 216627 298076 216693 298077
rect 216627 298012 216628 298076
rect 216692 298012 216693 298076
rect 216627 298011 216693 298012
rect 216075 262716 216141 262717
rect 216075 262652 216076 262716
rect 216140 262652 216141 262716
rect 216075 262651 216141 262652
rect 214787 228308 214853 228309
rect 214787 228244 214788 228308
rect 214852 228244 214853 228308
rect 214787 228243 214853 228244
rect 214603 180980 214669 180981
rect 214603 180916 214604 180980
rect 214668 180916 214669 180980
rect 214603 180915 214669 180916
rect 214419 179212 214485 179213
rect 214419 179148 214420 179212
rect 214484 179148 214485 179212
rect 214419 179147 214485 179148
rect 213131 167380 213197 167381
rect 213131 167316 213132 167380
rect 213196 167316 213197 167380
rect 213131 167315 213197 167316
rect 214790 166429 214850 228243
rect 216630 176221 216690 298011
rect 217182 177717 217242 339627
rect 217366 295357 217426 344931
rect 217550 296989 217610 345611
rect 217794 327454 218414 362898
rect 221514 367174 222134 388711
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 218651 344860 218717 344861
rect 218651 344796 218652 344860
rect 218716 344796 218717 344860
rect 218651 344795 218717 344796
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217547 296988 217613 296989
rect 217547 296924 217548 296988
rect 217612 296924 217613 296988
rect 217547 296923 217613 296924
rect 217363 295356 217429 295357
rect 217363 295292 217364 295356
rect 217428 295292 217429 295356
rect 217363 295291 217429 295292
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 219454 218414 254898
rect 218654 241501 218714 344795
rect 220307 342004 220373 342005
rect 220307 341940 220308 342004
rect 220372 341940 220373 342004
rect 220307 341939 220373 341940
rect 219939 339556 220005 339557
rect 219939 339492 219940 339556
rect 220004 339492 220005 339556
rect 219939 339491 220005 339492
rect 218835 339012 218901 339013
rect 218835 338948 218836 339012
rect 218900 338948 218901 339012
rect 218835 338947 218901 338948
rect 218838 246397 218898 338947
rect 218835 246396 218901 246397
rect 218835 246332 218836 246396
rect 218900 246332 218901 246396
rect 218835 246331 218901 246332
rect 218651 241500 218717 241501
rect 218651 241436 218652 241500
rect 218716 241436 218717 241500
rect 218651 241435 218717 241436
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217179 177716 217245 177717
rect 217179 177652 217180 177716
rect 217244 177652 217245 177716
rect 217179 177651 217245 177652
rect 216627 176220 216693 176221
rect 216627 176156 216628 176220
rect 216692 176156 216693 176220
rect 216627 176155 216693 176156
rect 214787 166428 214853 166429
rect 214787 166364 214788 166428
rect 214852 166364 214853 166428
rect 214787 166363 214853 166364
rect 207834 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 208454 137494
rect 207834 137174 208454 137258
rect 207834 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 208454 137174
rect 207834 101494 208454 136938
rect 207834 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 208454 101494
rect 207834 101174 208454 101258
rect 207834 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 208454 101174
rect 207834 65494 208454 100938
rect 207834 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 208454 65494
rect 207834 65174 208454 65258
rect 207834 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 208454 65174
rect 207834 29494 208454 64938
rect 207834 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 208454 29494
rect 207834 29174 208454 29258
rect 207834 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 208454 29174
rect 207834 -7066 208454 28938
rect 207834 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 208454 -7066
rect 207834 -7386 208454 -7302
rect 207834 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 208454 -7386
rect 207834 -7654 208454 -7622
rect 217794 147454 218414 182898
rect 219942 172821 220002 339491
rect 220123 337788 220189 337789
rect 220123 337724 220124 337788
rect 220188 337724 220189 337788
rect 220123 337723 220189 337724
rect 220126 275773 220186 337723
rect 220310 293725 220370 341939
rect 221227 340644 221293 340645
rect 221227 340580 221228 340644
rect 221292 340580 221293 340644
rect 221227 340579 221293 340580
rect 221043 340372 221109 340373
rect 221043 340308 221044 340372
rect 221108 340308 221109 340372
rect 221043 340307 221109 340308
rect 220491 338468 220557 338469
rect 220491 338404 220492 338468
rect 220556 338404 220557 338468
rect 220491 338403 220557 338404
rect 220307 293724 220373 293725
rect 220307 293660 220308 293724
rect 220372 293660 220373 293724
rect 220307 293659 220373 293660
rect 220494 290461 220554 338403
rect 220491 290460 220557 290461
rect 220491 290396 220492 290460
rect 220556 290396 220557 290460
rect 220491 290395 220557 290396
rect 220123 275772 220189 275773
rect 220123 275708 220124 275772
rect 220188 275708 220189 275772
rect 220123 275707 220189 275708
rect 221046 256189 221106 340307
rect 221043 256188 221109 256189
rect 221043 256124 221044 256188
rect 221108 256124 221109 256188
rect 221043 256123 221109 256124
rect 220859 255372 220925 255373
rect 220859 255308 220860 255372
rect 220924 255308 220925 255372
rect 220859 255307 220925 255308
rect 219939 172820 220005 172821
rect 219939 172756 219940 172820
rect 220004 172756 220005 172820
rect 219939 172755 220005 172756
rect 220862 171189 220922 255307
rect 221230 243133 221290 340579
rect 221514 331174 222134 366618
rect 225234 370894 225854 388711
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 223435 347580 223501 347581
rect 223435 347516 223436 347580
rect 223500 347516 223501 347580
rect 223435 347515 223501 347516
rect 222699 345404 222765 345405
rect 222699 345340 222700 345404
rect 222764 345340 222765 345404
rect 222699 345339 222765 345340
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221227 243132 221293 243133
rect 221227 243068 221228 243132
rect 221292 243068 221293 243132
rect 221227 243067 221293 243068
rect 221514 223174 222134 258618
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 220859 171188 220925 171189
rect 220859 171124 220860 171188
rect 220924 171124 220925 171188
rect 220859 171123 220925 171124
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 111454 218414 146898
rect 217794 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 218414 111454
rect 217794 111134 218414 111218
rect 217794 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 218414 111134
rect 217794 75454 218414 110898
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -7654 218414 -902
rect 221514 151174 222134 186618
rect 222702 164661 222762 345339
rect 222883 341188 222949 341189
rect 222883 341124 222884 341188
rect 222948 341124 222949 341188
rect 222883 341123 222949 341124
rect 222886 280669 222946 341123
rect 223438 335370 223498 347515
rect 224355 346900 224421 346901
rect 224355 346836 224356 346900
rect 224420 346836 224421 346900
rect 224355 346835 224421 346836
rect 224171 338196 224237 338197
rect 224171 338132 224172 338196
rect 224236 338132 224237 338196
rect 224171 338131 224237 338132
rect 223070 335310 223498 335370
rect 223070 298621 223130 335310
rect 223067 298620 223133 298621
rect 223067 298556 223068 298620
rect 223132 298556 223133 298620
rect 223067 298555 223133 298556
rect 222883 280668 222949 280669
rect 222883 280604 222884 280668
rect 222948 280604 222949 280668
rect 222883 280603 222949 280604
rect 223619 256732 223685 256733
rect 223619 256668 223620 256732
rect 223684 256668 223685 256732
rect 223619 256667 223685 256668
rect 223622 167925 223682 256667
rect 223803 254012 223869 254013
rect 223803 253948 223804 254012
rect 223868 253948 223869 254012
rect 223803 253947 223869 253948
rect 223806 169693 223866 253947
rect 224174 249661 224234 338131
rect 224358 257821 224418 346835
rect 224539 343908 224605 343909
rect 224539 343844 224540 343908
rect 224604 343844 224605 343908
rect 224539 343843 224605 343844
rect 224355 257820 224421 257821
rect 224355 257756 224356 257820
rect 224420 257756 224421 257820
rect 224355 257755 224421 257756
rect 224542 254557 224602 343843
rect 224723 342548 224789 342549
rect 224723 342484 224724 342548
rect 224788 342484 224789 342548
rect 224723 342483 224789 342484
rect 224539 254556 224605 254557
rect 224539 254492 224540 254556
rect 224604 254492 224605 254556
rect 224539 254491 224605 254492
rect 224726 252925 224786 342483
rect 224907 341596 224973 341597
rect 224907 341532 224908 341596
rect 224972 341532 224973 341596
rect 224907 341531 224973 341532
rect 224910 282437 224970 341531
rect 225234 334894 225854 370338
rect 228954 374614 229574 388711
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 227483 347988 227549 347989
rect 227483 347924 227484 347988
rect 227548 347924 227549 347988
rect 227483 347923 227549 347924
rect 226931 347852 226997 347853
rect 226931 347788 226932 347852
rect 226996 347788 226997 347852
rect 226931 347787 226997 347788
rect 226195 346220 226261 346221
rect 226195 346156 226196 346220
rect 226260 346156 226261 346220
rect 226195 346155 226261 346156
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 224907 282436 224973 282437
rect 224907 282372 224908 282436
rect 224972 282372 224973 282436
rect 224907 282371 224973 282372
rect 224907 282300 224973 282301
rect 224907 282236 224908 282300
rect 224972 282236 224973 282300
rect 224907 282235 224973 282236
rect 224723 252924 224789 252925
rect 224723 252860 224724 252924
rect 224788 252860 224789 252924
rect 224723 252859 224789 252860
rect 224171 249660 224237 249661
rect 224171 249596 224172 249660
rect 224236 249596 224237 249660
rect 224171 249595 224237 249596
rect 223803 169692 223869 169693
rect 223803 169628 223804 169692
rect 223868 169628 223869 169692
rect 223803 169627 223869 169628
rect 223619 167924 223685 167925
rect 223619 167860 223620 167924
rect 223684 167860 223685 167924
rect 223619 167859 223685 167860
rect 222699 164660 222765 164661
rect 222699 164596 222700 164660
rect 222764 164596 222765 164660
rect 222699 164595 222765 164596
rect 224910 163165 224970 282235
rect 225234 262894 225854 298338
rect 226198 296730 226258 346155
rect 226014 296670 226258 296730
rect 226014 288829 226074 296670
rect 226195 289780 226261 289781
rect 226195 289716 226196 289780
rect 226260 289716 226261 289780
rect 226195 289715 226261 289716
rect 226011 288828 226077 288829
rect 226011 288764 226012 288828
rect 226076 288764 226077 288828
rect 226011 288763 226077 288764
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 226894 225854 262338
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 224907 163164 224973 163165
rect 224907 163100 224908 163164
rect 224972 163100 224973 163164
rect 224907 163099 224973 163100
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 115174 222134 150618
rect 221514 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 222134 115174
rect 221514 114854 222134 114938
rect 221514 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 222134 114854
rect 221514 79174 222134 114618
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -1306 222134 6618
rect 221514 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 222134 -1306
rect 221514 -1626 222134 -1542
rect 221514 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 222134 -1626
rect 221514 -7654 222134 -1862
rect 225234 154894 225854 190338
rect 226198 174453 226258 289715
rect 226934 272509 226994 347787
rect 227115 346764 227181 346765
rect 227115 346700 227116 346764
rect 227180 346700 227181 346764
rect 227115 346699 227181 346700
rect 226931 272508 226997 272509
rect 226931 272444 226932 272508
rect 226996 272444 226997 272508
rect 226931 272443 226997 272444
rect 227118 270877 227178 346699
rect 227299 345404 227365 345405
rect 227299 345340 227300 345404
rect 227364 345340 227365 345404
rect 227299 345339 227365 345340
rect 227115 270876 227181 270877
rect 227115 270812 227116 270876
rect 227180 270812 227181 270876
rect 227115 270811 227181 270812
rect 227302 269245 227362 345339
rect 227486 274141 227546 347923
rect 228219 345540 228285 345541
rect 228219 345476 228220 345540
rect 228284 345476 228285 345540
rect 228219 345475 228285 345476
rect 228222 287197 228282 345475
rect 228954 338614 229574 374058
rect 232674 378334 233294 388711
rect 232674 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 233294 378334
rect 232674 378014 233294 378098
rect 232674 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 233294 378014
rect 231163 353564 231229 353565
rect 231163 353500 231164 353564
rect 231228 353500 231229 353564
rect 231163 353499 231229 353500
rect 229875 351116 229941 351117
rect 229875 351052 229876 351116
rect 229940 351052 229941 351116
rect 229875 351051 229941 351052
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228219 287196 228285 287197
rect 228219 287132 228220 287196
rect 228284 287132 228285 287196
rect 228219 287131 228285 287132
rect 227483 274140 227549 274141
rect 227483 274076 227484 274140
rect 227548 274076 227549 274140
rect 227483 274075 227549 274076
rect 227299 269244 227365 269245
rect 227299 269180 227300 269244
rect 227364 269180 227365 269244
rect 227299 269179 227365 269180
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 226195 174452 226261 174453
rect 226195 174388 226196 174452
rect 226260 174388 226261 174452
rect 226195 174387 226261 174388
rect 228219 170644 228285 170645
rect 228219 170580 228220 170644
rect 228284 170580 228285 170644
rect 228219 170579 228285 170580
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 118894 225854 154338
rect 225234 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 225854 118894
rect 225234 118574 225854 118658
rect 225234 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 225854 118574
rect 225234 82894 225854 118338
rect 228222 86325 228282 170579
rect 228954 158614 229574 194058
rect 229878 166293 229938 351051
rect 230243 339556 230309 339557
rect 230243 339492 230244 339556
rect 230308 339492 230309 339556
rect 230243 339491 230309 339492
rect 230059 252516 230125 252517
rect 230059 252452 230060 252516
rect 230124 252452 230125 252516
rect 230059 252451 230125 252452
rect 229875 166292 229941 166293
rect 229875 166228 229876 166292
rect 229940 166228 229941 166292
rect 229875 166227 229941 166228
rect 230062 161397 230122 252451
rect 230246 251293 230306 339491
rect 230979 338740 231045 338741
rect 230979 338676 230980 338740
rect 231044 338676 231045 338740
rect 230979 338675 231045 338676
rect 230243 251292 230309 251293
rect 230243 251228 230244 251292
rect 230308 251228 230309 251292
rect 230243 251227 230309 251228
rect 230982 165205 231042 338675
rect 231166 244765 231226 353499
rect 231347 342820 231413 342821
rect 231347 342756 231348 342820
rect 231412 342756 231413 342820
rect 231347 342755 231413 342756
rect 231350 267613 231410 342755
rect 232674 342334 233294 377778
rect 236394 382054 237014 388711
rect 236394 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 237014 382054
rect 236394 381734 237014 381818
rect 236394 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 237014 381734
rect 234475 377500 234541 377501
rect 234475 377436 234476 377500
rect 234540 377436 234541 377500
rect 234475 377435 234541 377436
rect 234291 366484 234357 366485
rect 234291 366420 234292 366484
rect 234356 366420 234357 366484
rect 234291 366419 234357 366420
rect 234107 364988 234173 364989
rect 234107 364924 234108 364988
rect 234172 364924 234173 364988
rect 234107 364923 234173 364924
rect 232674 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 233294 342334
rect 232674 342014 233294 342098
rect 232674 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 233294 342014
rect 231531 341052 231597 341053
rect 231531 340988 231532 341052
rect 231596 340988 231597 341052
rect 231531 340987 231597 340988
rect 231534 285565 231594 340987
rect 232674 306334 233294 341778
rect 234110 309909 234170 364923
rect 234107 309908 234173 309909
rect 234107 309844 234108 309908
rect 234172 309844 234173 309908
rect 234107 309843 234173 309844
rect 232674 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 233294 306334
rect 232674 306014 233294 306098
rect 232674 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 233294 306014
rect 231531 285564 231597 285565
rect 231531 285500 231532 285564
rect 231596 285500 231597 285564
rect 231531 285499 231597 285500
rect 232674 270334 233294 305778
rect 234294 284885 234354 366419
rect 234478 287061 234538 377435
rect 235763 353836 235829 353837
rect 235763 353772 235764 353836
rect 235828 353772 235829 353836
rect 235763 353771 235829 353772
rect 235211 349212 235277 349213
rect 235211 349148 235212 349212
rect 235276 349148 235277 349212
rect 235211 349147 235277 349148
rect 234475 287060 234541 287061
rect 234475 286996 234476 287060
rect 234540 286996 234541 287060
rect 234475 286995 234541 286996
rect 234291 284884 234357 284885
rect 234291 284820 234292 284884
rect 234356 284820 234357 284884
rect 234291 284819 234357 284820
rect 232674 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 233294 270334
rect 232674 270014 233294 270098
rect 232674 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 233294 270014
rect 231347 267612 231413 267613
rect 231347 267548 231348 267612
rect 231412 267548 231413 267612
rect 231347 267547 231413 267548
rect 231163 244764 231229 244765
rect 231163 244700 231164 244764
rect 231228 244700 231229 244764
rect 231163 244699 231229 244700
rect 232674 234334 233294 269778
rect 232674 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 233294 234334
rect 232674 234014 233294 234098
rect 232674 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 233294 234014
rect 232674 198334 233294 233778
rect 234659 201924 234725 201925
rect 234659 201860 234660 201924
rect 234724 201860 234725 201924
rect 234659 201859 234725 201860
rect 232674 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 233294 198334
rect 232674 198014 233294 198098
rect 232674 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 233294 198014
rect 231163 171732 231229 171733
rect 231163 171668 231164 171732
rect 231228 171668 231229 171732
rect 231163 171667 231229 171668
rect 230979 165204 231045 165205
rect 230979 165140 230980 165204
rect 231044 165140 231045 165204
rect 230979 165139 231045 165140
rect 230059 161396 230125 161397
rect 230059 161332 230060 161396
rect 230124 161332 230125 161396
rect 230059 161331 230125 161332
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228219 86324 228285 86325
rect 228219 86260 228220 86324
rect 228284 86260 228285 86324
rect 228219 86259 228285 86260
rect 228954 86294 229574 86378
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -2266 225854 10338
rect 225234 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 225854 -2266
rect 225234 -2586 225854 -2502
rect 225234 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 225854 -2586
rect 225234 -7654 225854 -2822
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 231166 45525 231226 171667
rect 232674 162334 233294 197778
rect 232674 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 233294 162334
rect 232674 162014 233294 162098
rect 232674 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 233294 162014
rect 232674 126334 233294 161778
rect 234662 155957 234722 201859
rect 235214 156637 235274 349147
rect 235766 283797 235826 353771
rect 236394 346054 237014 381498
rect 240114 385774 240734 388711
rect 240114 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 240734 385774
rect 240114 385454 240734 385538
rect 240114 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 240734 385454
rect 239811 380220 239877 380221
rect 239811 380156 239812 380220
rect 239876 380156 239877 380220
rect 239811 380155 239877 380156
rect 239627 362268 239693 362269
rect 239627 362204 239628 362268
rect 239692 362204 239693 362268
rect 239627 362203 239693 362204
rect 239443 361044 239509 361045
rect 239443 360980 239444 361044
rect 239508 360980 239509 361044
rect 239443 360979 239509 360980
rect 239259 353428 239325 353429
rect 239259 353364 239260 353428
rect 239324 353364 239325 353428
rect 239259 353363 239325 353364
rect 236394 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 237014 346054
rect 236394 345734 237014 345818
rect 236394 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 237014 345734
rect 236394 310054 237014 345498
rect 237971 340236 238037 340237
rect 237971 340172 237972 340236
rect 238036 340172 238037 340236
rect 237971 340171 238037 340172
rect 238155 340236 238221 340237
rect 238155 340172 238156 340236
rect 238220 340172 238221 340236
rect 238155 340171 238221 340172
rect 236394 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 237014 310054
rect 236394 309734 237014 309818
rect 236394 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 237014 309734
rect 235763 283796 235829 283797
rect 235763 283732 235764 283796
rect 235828 283732 235829 283796
rect 235763 283731 235829 283732
rect 236394 274054 237014 309498
rect 236394 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 237014 274054
rect 236394 273734 237014 273818
rect 236394 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 237014 273734
rect 236394 238054 237014 273498
rect 237787 239188 237853 239189
rect 237787 239124 237788 239188
rect 237852 239124 237853 239188
rect 237787 239123 237853 239124
rect 236394 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 237014 238054
rect 237603 238100 237669 238101
rect 237603 238036 237604 238100
rect 237668 238036 237669 238100
rect 237603 238035 237669 238036
rect 236394 237734 237014 237818
rect 236394 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 237014 237734
rect 236394 202054 237014 237498
rect 237419 231572 237485 231573
rect 237419 231508 237420 231572
rect 237484 231508 237485 231572
rect 237419 231507 237485 231508
rect 237422 226949 237482 231507
rect 237606 231165 237666 238035
rect 237603 231164 237669 231165
rect 237603 231100 237604 231164
rect 237668 231100 237669 231164
rect 237603 231099 237669 231100
rect 237419 226948 237485 226949
rect 237419 226884 237420 226948
rect 237484 226884 237485 226948
rect 237419 226883 237485 226884
rect 237790 225589 237850 239123
rect 237974 236061 238034 340171
rect 238158 339557 238218 340171
rect 238155 339556 238221 339557
rect 238155 339492 238156 339556
rect 238220 339492 238221 339556
rect 238155 339491 238221 339492
rect 238339 246804 238405 246805
rect 238339 246740 238340 246804
rect 238404 246740 238405 246804
rect 238339 246739 238405 246740
rect 238155 237012 238221 237013
rect 238155 236948 238156 237012
rect 238220 236948 238221 237012
rect 238155 236947 238221 236948
rect 237971 236060 238037 236061
rect 237971 235996 237972 236060
rect 238036 235996 238037 236060
rect 237971 235995 238037 235996
rect 237971 234836 238037 234837
rect 237971 234772 237972 234836
rect 238036 234772 238037 234836
rect 237971 234771 238037 234772
rect 237787 225588 237853 225589
rect 237787 225524 237788 225588
rect 237852 225524 237853 225588
rect 237787 225523 237853 225524
rect 237974 207637 238034 234771
rect 237971 207636 238037 207637
rect 237971 207572 237972 207636
rect 238036 207572 238037 207636
rect 237971 207571 238037 207572
rect 236394 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 237014 202054
rect 236394 201734 237014 201818
rect 236394 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 237014 201734
rect 235395 185604 235461 185605
rect 235395 185540 235396 185604
rect 235460 185540 235461 185604
rect 235395 185539 235461 185540
rect 235398 168469 235458 185539
rect 235395 168468 235461 168469
rect 235395 168404 235396 168468
rect 235460 168404 235461 168468
rect 235395 168403 235461 168404
rect 236394 166054 237014 201498
rect 238158 195261 238218 236947
rect 238342 235245 238402 246739
rect 238339 235244 238405 235245
rect 238339 235180 238340 235244
rect 238404 235180 238405 235244
rect 238339 235179 238405 235180
rect 238523 226404 238589 226405
rect 238523 226340 238524 226404
rect 238588 226340 238589 226404
rect 238523 226339 238589 226340
rect 238155 195260 238221 195261
rect 238155 195196 238156 195260
rect 238220 195196 238221 195260
rect 238155 195195 238221 195196
rect 237971 193900 238037 193901
rect 237971 193836 237972 193900
rect 238036 193836 238037 193900
rect 237971 193835 238037 193836
rect 237419 192540 237485 192541
rect 237419 192476 237420 192540
rect 237484 192476 237485 192540
rect 237419 192475 237485 192476
rect 237422 187781 237482 192475
rect 237419 187780 237485 187781
rect 237419 187716 237420 187780
rect 237484 187716 237485 187780
rect 237419 187715 237485 187716
rect 236394 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 237014 166054
rect 236394 165734 237014 165818
rect 236394 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 237014 165734
rect 235579 159764 235645 159765
rect 235579 159700 235580 159764
rect 235644 159700 235645 159764
rect 235579 159699 235645 159700
rect 235211 156636 235277 156637
rect 235211 156572 235212 156636
rect 235276 156572 235277 156636
rect 235211 156571 235277 156572
rect 235395 156500 235461 156501
rect 235395 156436 235396 156500
rect 235460 156436 235461 156500
rect 235395 156435 235461 156436
rect 234659 155956 234725 155957
rect 234659 155892 234660 155956
rect 234724 155892 234725 155956
rect 234659 155891 234725 155892
rect 235211 154868 235277 154869
rect 235211 154804 235212 154868
rect 235276 154804 235277 154868
rect 235211 154803 235277 154804
rect 232674 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 233294 126334
rect 232674 126014 233294 126098
rect 232674 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 233294 126014
rect 232674 90334 233294 125778
rect 234659 120596 234725 120597
rect 234659 120532 234660 120596
rect 234724 120532 234725 120596
rect 234659 120531 234725 120532
rect 232674 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 233294 90334
rect 232674 90014 233294 90098
rect 232674 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 233294 90014
rect 232674 54334 233294 89778
rect 232674 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 233294 54334
rect 232674 54014 233294 54098
rect 232674 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 233294 54014
rect 231163 45524 231229 45525
rect 231163 45460 231164 45524
rect 231228 45460 231229 45524
rect 231163 45459 231229 45460
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 228954 -3226 229574 14058
rect 228954 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 229574 -3226
rect 228954 -3546 229574 -3462
rect 228954 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 229574 -3546
rect 228954 -7654 229574 -3782
rect 232674 18334 233294 53778
rect 232674 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 233294 18334
rect 232674 18014 233294 18098
rect 232674 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 233294 18014
rect 232674 -4186 233294 17778
rect 234662 7717 234722 120531
rect 235214 120189 235274 154803
rect 235211 120188 235277 120189
rect 235211 120124 235212 120188
rect 235276 120124 235277 120188
rect 235211 120123 235277 120124
rect 235398 115293 235458 156435
rect 235582 118557 235642 159699
rect 235763 158132 235829 158133
rect 235763 158068 235764 158132
rect 235828 158068 235829 158132
rect 235763 158067 235829 158068
rect 235766 119373 235826 158067
rect 236394 130054 237014 165498
rect 237974 160853 238034 193835
rect 238155 191044 238221 191045
rect 238155 190980 238156 191044
rect 238220 190980 238221 191044
rect 238155 190979 238221 190980
rect 237971 160852 238037 160853
rect 237971 160788 237972 160852
rect 238036 160788 238037 160852
rect 237971 160787 238037 160788
rect 238158 159765 238218 190979
rect 238339 188324 238405 188325
rect 238339 188260 238340 188324
rect 238404 188260 238405 188324
rect 238339 188259 238405 188260
rect 238342 161941 238402 188259
rect 238339 161940 238405 161941
rect 238339 161876 238340 161940
rect 238404 161876 238405 161940
rect 238339 161875 238405 161876
rect 238155 159764 238221 159765
rect 238155 159700 238156 159764
rect 238220 159700 238221 159764
rect 238155 159699 238221 159700
rect 238155 151604 238221 151605
rect 238155 151540 238156 151604
rect 238220 151540 238221 151604
rect 238155 151539 238221 151540
rect 237971 149972 238037 149973
rect 237971 149908 237972 149972
rect 238036 149908 238037 149972
rect 237971 149907 238037 149908
rect 236394 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 237014 130054
rect 236394 129734 237014 129818
rect 236394 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 237014 129734
rect 235763 119372 235829 119373
rect 235763 119308 235764 119372
rect 235828 119308 235829 119372
rect 235763 119307 235829 119308
rect 235579 118556 235645 118557
rect 235579 118492 235580 118556
rect 235644 118492 235645 118556
rect 235579 118491 235645 118492
rect 235395 115292 235461 115293
rect 235395 115228 235396 115292
rect 235460 115228 235461 115292
rect 235395 115227 235461 115228
rect 236394 94054 237014 129498
rect 237787 123860 237853 123861
rect 237787 123796 237788 123860
rect 237852 123796 237853 123860
rect 237787 123795 237853 123796
rect 237790 117469 237850 123795
rect 237974 118421 238034 149907
rect 238158 119373 238218 151539
rect 238526 141405 238586 226339
rect 239262 143170 239322 353363
rect 239446 143850 239506 360979
rect 239630 144601 239690 362203
rect 239814 145689 239874 380155
rect 240114 349774 240734 385218
rect 240114 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 240734 349774
rect 240114 349454 240734 349538
rect 240114 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 240734 349454
rect 240114 336713 240734 349218
rect 264954 374614 265574 388711
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 256003 339556 256069 339557
rect 256003 339492 256004 339556
rect 256068 339492 256069 339556
rect 256003 339491 256069 339492
rect 256006 339013 256066 339491
rect 256003 339012 256069 339013
rect 256003 338948 256004 339012
rect 256068 338948 256069 339012
rect 256003 338947 256069 338948
rect 264954 338614 265574 374058
rect 268674 378334 269294 388711
rect 268674 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 269294 378334
rect 268674 378014 269294 378098
rect 268674 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 269294 378014
rect 268674 342334 269294 377778
rect 268674 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 269294 342334
rect 268674 342014 269294 342098
rect 268674 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 269294 342014
rect 267595 340372 267661 340373
rect 267595 340308 267596 340372
rect 267660 340308 267661 340372
rect 267595 340307 267661 340308
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 267598 338605 267658 340307
rect 267595 338604 267661 338605
rect 267595 338540 267596 338604
rect 267660 338540 267661 338604
rect 267595 338539 267661 338540
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 336713 265574 338058
rect 268674 336713 269294 341778
rect 272394 382054 273014 388711
rect 272394 381818 272426 382054
rect 272662 381818 272746 382054
rect 272982 381818 273014 382054
rect 272394 381734 273014 381818
rect 272394 381498 272426 381734
rect 272662 381498 272746 381734
rect 272982 381498 273014 381734
rect 272394 346054 273014 381498
rect 272394 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 273014 346054
rect 272394 345734 273014 345818
rect 272394 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 273014 345734
rect 272394 336713 273014 345498
rect 276114 385774 276734 388711
rect 276114 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 276734 385774
rect 276114 385454 276734 385538
rect 276114 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 276734 385454
rect 276114 349774 276734 385218
rect 284891 375188 284957 375189
rect 284891 375124 284892 375188
rect 284956 375124 284957 375188
rect 284891 375123 284957 375124
rect 282131 374780 282197 374781
rect 282131 374716 282132 374780
rect 282196 374716 282197 374780
rect 282131 374715 282197 374716
rect 276114 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 276734 349774
rect 276114 349454 276734 349538
rect 276114 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 276734 349454
rect 274587 339556 274653 339557
rect 274587 339492 274588 339556
rect 274652 339492 274653 339556
rect 274587 339491 274653 339492
rect 274590 339013 274650 339491
rect 274587 339012 274653 339013
rect 274587 338948 274588 339012
rect 274652 338948 274653 339012
rect 274587 338947 274653 338948
rect 276114 336713 276734 349218
rect 279003 346900 279069 346901
rect 279003 346836 279004 346900
rect 279068 346836 279069 346900
rect 279003 346835 279069 346836
rect 279006 339421 279066 346835
rect 280659 345676 280725 345677
rect 280659 345612 280660 345676
rect 280724 345612 280725 345676
rect 280659 345611 280725 345612
rect 279555 341596 279621 341597
rect 279555 341532 279556 341596
rect 279620 341532 279621 341596
rect 279555 341531 279621 341532
rect 279003 339420 279069 339421
rect 279003 339356 279004 339420
rect 279068 339356 279069 339420
rect 279003 339355 279069 339356
rect 279558 338061 279618 341531
rect 280291 341188 280357 341189
rect 280291 341124 280292 341188
rect 280356 341124 280357 341188
rect 280291 341123 280357 341124
rect 279923 340644 279989 340645
rect 279923 340580 279924 340644
rect 279988 340580 279989 340644
rect 279923 340579 279989 340580
rect 279739 340372 279805 340373
rect 279739 340308 279740 340372
rect 279804 340308 279805 340372
rect 279739 340307 279805 340308
rect 279555 338060 279621 338061
rect 279555 337996 279556 338060
rect 279620 337996 279621 338060
rect 279555 337995 279621 337996
rect 279742 337925 279802 340307
rect 279926 338877 279986 340579
rect 280107 340236 280173 340237
rect 280107 340172 280108 340236
rect 280172 340172 280173 340236
rect 280107 340171 280173 340172
rect 279923 338876 279989 338877
rect 279923 338812 279924 338876
rect 279988 338812 279989 338876
rect 279923 338811 279989 338812
rect 279739 337924 279805 337925
rect 279739 337860 279740 337924
rect 279804 337860 279805 337924
rect 279739 337859 279805 337860
rect 259568 331174 259888 331206
rect 259568 330938 259610 331174
rect 259846 330938 259888 331174
rect 259568 330854 259888 330938
rect 259568 330618 259610 330854
rect 259846 330618 259888 330854
rect 259568 330586 259888 330618
rect 244208 327454 244528 327486
rect 244208 327218 244250 327454
rect 244486 327218 244528 327454
rect 244208 327134 244528 327218
rect 244208 326898 244250 327134
rect 244486 326898 244528 327134
rect 244208 326866 244528 326898
rect 274928 327454 275248 327486
rect 274928 327218 274970 327454
rect 275206 327218 275248 327454
rect 274928 327134 275248 327218
rect 274928 326898 274970 327134
rect 275206 326898 275248 327134
rect 274928 326866 275248 326898
rect 259568 295174 259888 295206
rect 259568 294938 259610 295174
rect 259846 294938 259888 295174
rect 259568 294854 259888 294938
rect 259568 294618 259610 294854
rect 259846 294618 259888 294854
rect 259568 294586 259888 294618
rect 244208 291454 244528 291486
rect 244208 291218 244250 291454
rect 244486 291218 244528 291454
rect 244208 291134 244528 291218
rect 244208 290898 244250 291134
rect 244486 290898 244528 291134
rect 244208 290866 244528 290898
rect 274928 291454 275248 291486
rect 274928 291218 274970 291454
rect 275206 291218 275248 291454
rect 274928 291134 275248 291218
rect 274928 290898 274970 291134
rect 275206 290898 275248 291134
rect 274928 290866 275248 290898
rect 259568 259174 259888 259206
rect 259568 258938 259610 259174
rect 259846 258938 259888 259174
rect 259568 258854 259888 258938
rect 259568 258618 259610 258854
rect 259846 258618 259888 258854
rect 259568 258586 259888 258618
rect 244208 255454 244528 255486
rect 244208 255218 244250 255454
rect 244486 255218 244528 255454
rect 244208 255134 244528 255218
rect 244208 254898 244250 255134
rect 244486 254898 244528 255134
rect 244208 254866 244528 254898
rect 274928 255454 275248 255486
rect 274928 255218 274970 255454
rect 275206 255218 275248 255454
rect 274928 255134 275248 255218
rect 274928 254898 274970 255134
rect 275206 254898 275248 255134
rect 274928 254866 275248 254898
rect 280110 238770 280170 340171
rect 280294 243541 280354 341123
rect 280662 335370 280722 345611
rect 280478 335310 280722 335370
rect 280478 309365 280538 335310
rect 280475 309364 280541 309365
rect 280475 309300 280476 309364
rect 280540 309300 280541 309364
rect 280475 309299 280541 309300
rect 282134 272373 282194 374715
rect 282315 373420 282381 373421
rect 282315 373356 282316 373420
rect 282380 373356 282381 373420
rect 282315 373355 282381 373356
rect 282318 274549 282378 373355
rect 282683 370564 282749 370565
rect 282683 370500 282684 370564
rect 282748 370500 282749 370564
rect 282683 370499 282749 370500
rect 282499 369068 282565 369069
rect 282499 369004 282500 369068
rect 282564 369004 282565 369068
rect 282499 369003 282565 369004
rect 282315 274548 282381 274549
rect 282315 274484 282316 274548
rect 282380 274484 282381 274548
rect 282315 274483 282381 274484
rect 282131 272372 282197 272373
rect 282131 272308 282132 272372
rect 282196 272308 282197 272372
rect 282131 272307 282197 272308
rect 282502 270741 282562 369003
rect 282686 273461 282746 370499
rect 282867 357508 282933 357509
rect 282867 357444 282868 357508
rect 282932 357444 282933 357508
rect 282867 357443 282933 357444
rect 282683 273460 282749 273461
rect 282683 273396 282684 273460
rect 282748 273396 282749 273460
rect 282683 273395 282749 273396
rect 282499 270740 282565 270741
rect 282499 270676 282500 270740
rect 282564 270676 282565 270740
rect 282499 270675 282565 270676
rect 280291 243540 280357 243541
rect 280291 243476 280292 243540
rect 280356 243476 280357 243540
rect 280291 243475 280357 243476
rect 280110 238710 280354 238770
rect 280294 233749 280354 238710
rect 280291 233748 280357 233749
rect 280291 233684 280292 233748
rect 280356 233684 280357 233748
rect 280291 233683 280357 233684
rect 259568 223174 259888 223206
rect 259568 222938 259610 223174
rect 259846 222938 259888 223174
rect 259568 222854 259888 222938
rect 259568 222618 259610 222854
rect 259846 222618 259888 222854
rect 259568 222586 259888 222618
rect 244208 219454 244528 219486
rect 244208 219218 244250 219454
rect 244486 219218 244528 219454
rect 244208 219134 244528 219218
rect 244208 218898 244250 219134
rect 244486 218898 244528 219134
rect 244208 218866 244528 218898
rect 274928 219454 275248 219486
rect 274928 219218 274970 219454
rect 275206 219218 275248 219454
rect 274928 219134 275248 219218
rect 274928 218898 274970 219134
rect 275206 218898 275248 219134
rect 274928 218866 275248 218898
rect 281763 214708 281829 214709
rect 281763 214644 281764 214708
rect 281828 214644 281829 214708
rect 281763 214643 281829 214644
rect 280843 208724 280909 208725
rect 280843 208660 280844 208724
rect 280908 208660 280909 208724
rect 280843 208659 280909 208660
rect 280659 197300 280725 197301
rect 280659 197236 280660 197300
rect 280724 197236 280725 197300
rect 280659 197235 280725 197236
rect 259568 187174 259888 187206
rect 259568 186938 259610 187174
rect 259846 186938 259888 187174
rect 259568 186854 259888 186938
rect 259568 186618 259610 186854
rect 259846 186618 259888 186854
rect 259568 186586 259888 186618
rect 244208 183454 244528 183486
rect 244208 183218 244250 183454
rect 244486 183218 244528 183454
rect 244208 183134 244528 183218
rect 244208 182898 244250 183134
rect 244486 182898 244528 183134
rect 244208 182866 244528 182898
rect 274928 183454 275248 183486
rect 274928 183218 274970 183454
rect 275206 183218 275248 183454
rect 274928 183134 275248 183218
rect 274928 182898 274970 183134
rect 275206 182898 275248 183134
rect 274928 182866 275248 182898
rect 259568 151174 259888 151206
rect 259568 150938 259610 151174
rect 259846 150938 259888 151174
rect 259568 150854 259888 150938
rect 259568 150618 259610 150854
rect 259846 150618 259888 150854
rect 259568 150586 259888 150618
rect 244208 147454 244528 147486
rect 244208 147218 244250 147454
rect 244486 147218 244528 147454
rect 244208 147134 244528 147218
rect 244208 146898 244250 147134
rect 244486 146898 244528 147134
rect 244208 146866 244528 146898
rect 274928 147454 275248 147486
rect 274928 147218 274970 147454
rect 275206 147218 275248 147454
rect 274928 147134 275248 147218
rect 274928 146898 274970 147134
rect 275206 146898 275248 147134
rect 274928 146866 275248 146898
rect 239811 145688 239877 145689
rect 239811 145624 239812 145688
rect 239876 145624 239877 145688
rect 239811 145623 239877 145624
rect 239627 144600 239693 144601
rect 239627 144536 239628 144600
rect 239692 144536 239693 144600
rect 239627 144535 239693 144536
rect 239446 143790 239874 143850
rect 239814 143513 239874 143790
rect 239811 143512 239877 143513
rect 239811 143448 239812 143512
rect 239876 143448 239877 143512
rect 239811 143447 239877 143448
rect 239262 143110 239690 143170
rect 239630 142425 239690 143110
rect 239627 142424 239693 142425
rect 239627 142360 239628 142424
rect 239692 142360 239693 142424
rect 239627 142359 239693 142360
rect 238523 141404 238589 141405
rect 238523 141340 238524 141404
rect 238588 141340 238589 141404
rect 238523 141339 238589 141340
rect 238339 136916 238405 136917
rect 238339 136852 238340 136916
rect 238404 136852 238405 136916
rect 238339 136851 238405 136852
rect 238342 123589 238402 136851
rect 238523 135828 238589 135829
rect 238523 135764 238524 135828
rect 238588 135764 238589 135828
rect 238523 135763 238589 135764
rect 238339 123588 238405 123589
rect 238339 123524 238340 123588
rect 238404 123524 238405 123588
rect 238339 123523 238405 123524
rect 238526 120053 238586 135763
rect 280107 135148 280173 135149
rect 280107 135084 280108 135148
rect 280172 135084 280173 135148
rect 280107 135083 280173 135084
rect 239627 134808 239693 134809
rect 239627 134744 239628 134808
rect 239692 134744 239693 134808
rect 239627 134743 239693 134744
rect 239443 133652 239509 133653
rect 239443 133588 239444 133652
rect 239508 133588 239509 133652
rect 239443 133587 239509 133588
rect 238523 120052 238589 120053
rect 238523 119988 238524 120052
rect 238588 119988 238589 120052
rect 238523 119987 238589 119988
rect 238155 119372 238221 119373
rect 238155 119308 238156 119372
rect 238220 119308 238221 119372
rect 238155 119307 238221 119308
rect 237971 118420 238037 118421
rect 237971 118356 237972 118420
rect 238036 118356 238037 118420
rect 237971 118355 238037 118356
rect 237787 117468 237853 117469
rect 237787 117404 237788 117468
rect 237852 117404 237853 117468
rect 237787 117403 237853 117404
rect 239446 98701 239506 133587
rect 239630 100741 239690 134743
rect 280110 134330 280170 135083
rect 278822 134270 280170 134330
rect 239811 132632 239877 132633
rect 239811 132568 239812 132632
rect 239876 132568 239877 132632
rect 239811 132567 239877 132568
rect 239627 100740 239693 100741
rect 239627 100676 239628 100740
rect 239692 100676 239693 100740
rect 239627 100675 239693 100676
rect 239443 98700 239509 98701
rect 239443 98636 239444 98700
rect 239508 98636 239509 98700
rect 239443 98635 239509 98636
rect 236394 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 237014 94054
rect 236394 93734 237014 93818
rect 236394 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 237014 93734
rect 236394 58054 237014 93498
rect 236394 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 237014 58054
rect 236394 57734 237014 57818
rect 236394 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 237014 57734
rect 236394 22054 237014 57498
rect 239814 33149 239874 132567
rect 240114 97774 240734 132447
rect 240114 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 240734 97774
rect 240114 97454 240734 97538
rect 240114 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 240734 97454
rect 240114 61774 240734 97218
rect 240114 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 240734 61774
rect 240114 61454 240734 61538
rect 240114 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 240734 61454
rect 239811 33148 239877 33149
rect 239811 33084 239812 33148
rect 239876 33084 239877 33148
rect 239811 33083 239877 33084
rect 236394 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 237014 22054
rect 236394 21734 237014 21818
rect 236394 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 237014 21734
rect 234659 7716 234725 7717
rect 234659 7652 234660 7716
rect 234724 7652 234725 7716
rect 234659 7651 234725 7652
rect 232674 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 233294 -4186
rect 232674 -4506 233294 -4422
rect 232674 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 233294 -4506
rect 232674 -7654 233294 -4742
rect 236394 -5146 237014 21498
rect 236394 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 237014 -5146
rect 236394 -5466 237014 -5382
rect 236394 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 237014 -5466
rect 236394 -7654 237014 -5702
rect 240114 25774 240734 61218
rect 240114 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 240734 25774
rect 240114 25454 240734 25538
rect 240114 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 240734 25454
rect 240114 -6106 240734 25218
rect 240114 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 240734 -6106
rect 240114 -6426 240734 -6342
rect 240114 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 240734 -6426
rect 240114 -7654 240734 -6662
rect 243834 101494 244454 119988
rect 243834 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 244454 101494
rect 243834 101174 244454 101258
rect 243834 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 244454 101174
rect 243834 65494 244454 100938
rect 243834 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 244454 65494
rect 243834 65174 244454 65258
rect 243834 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 244454 65174
rect 243834 29494 244454 64938
rect 243834 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 244454 29494
rect 243834 29174 244454 29258
rect 243834 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 244454 29174
rect 243834 -7066 244454 28938
rect 243834 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 244454 -7066
rect 243834 -7386 244454 -7302
rect 243834 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 244454 -7386
rect 243834 -7654 244454 -7622
rect 253794 111454 254414 132447
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -7654 254414 -902
rect 257514 115174 258134 132447
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -1306 258134 6618
rect 257514 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 258134 -1306
rect 257514 -1626 258134 -1542
rect 257514 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 258134 -1626
rect 257514 -7654 258134 -1862
rect 261234 118894 261854 132447
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -2266 261854 10338
rect 261234 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 261854 -2266
rect 261234 -2586 261854 -2502
rect 261234 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 261854 -2586
rect 261234 -7654 261854 -2822
rect 264954 122614 265574 132447
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 264954 -3226 265574 14058
rect 264954 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 265574 -3226
rect 264954 -3546 265574 -3462
rect 264954 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 265574 -3546
rect 264954 -7654 265574 -3782
rect 268674 126334 269294 132447
rect 268674 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 269294 126334
rect 268674 126014 269294 126098
rect 268674 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 269294 126014
rect 268674 90334 269294 125778
rect 268674 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 269294 90334
rect 268674 90014 269294 90098
rect 268674 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 269294 90014
rect 268674 54334 269294 89778
rect 268674 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 269294 54334
rect 268674 54014 269294 54098
rect 268674 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 269294 54014
rect 268674 18334 269294 53778
rect 268674 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 269294 18334
rect 268674 18014 269294 18098
rect 268674 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 269294 18014
rect 268674 -4186 269294 17778
rect 268674 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 269294 -4186
rect 268674 -4506 269294 -4422
rect 268674 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 269294 -4506
rect 268674 -7654 269294 -4742
rect 272394 130054 273014 132447
rect 272394 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 273014 130054
rect 272394 129734 273014 129818
rect 272394 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 273014 129734
rect 272394 94054 273014 129498
rect 272394 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 273014 94054
rect 272394 93734 273014 93818
rect 272394 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 273014 93734
rect 272394 58054 273014 93498
rect 272394 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 273014 58054
rect 272394 57734 273014 57818
rect 272394 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 273014 57734
rect 272394 22054 273014 57498
rect 272394 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 273014 22054
rect 272394 21734 273014 21818
rect 272394 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 273014 21734
rect 272394 -5146 273014 21498
rect 272394 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 273014 -5146
rect 272394 -5466 273014 -5382
rect 272394 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 273014 -5466
rect 272394 -7654 273014 -5702
rect 276114 97774 276734 132447
rect 276114 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 276734 97774
rect 276114 97454 276734 97538
rect 276114 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 276734 97454
rect 276114 61774 276734 97218
rect 278822 94485 278882 134270
rect 279834 101494 280454 132447
rect 279834 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 280454 101494
rect 279834 101174 280454 101258
rect 279834 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 280454 101174
rect 278819 94484 278885 94485
rect 278819 94420 278820 94484
rect 278884 94420 278885 94484
rect 278819 94419 278885 94420
rect 276114 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 276734 61774
rect 276114 61454 276734 61538
rect 276114 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 276734 61454
rect 276114 25774 276734 61218
rect 276114 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 276734 25774
rect 276114 25454 276734 25538
rect 276114 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 276734 25454
rect 276114 -6106 276734 25218
rect 276114 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 276734 -6106
rect 276114 -6426 276734 -6342
rect 276114 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 276734 -6426
rect 276114 -7654 276734 -6662
rect 279834 65494 280454 100938
rect 279834 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 280454 65494
rect 279834 65174 280454 65258
rect 279834 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 280454 65174
rect 279834 29494 280454 64938
rect 280662 44981 280722 197235
rect 280846 116653 280906 208659
rect 281579 198932 281645 198933
rect 281579 198868 281580 198932
rect 281644 198868 281645 198932
rect 281579 198867 281645 198868
rect 281027 191316 281093 191317
rect 281027 191252 281028 191316
rect 281092 191252 281093 191316
rect 281027 191251 281093 191252
rect 280843 116652 280909 116653
rect 280843 116588 280844 116652
rect 280908 116588 280909 116652
rect 280843 116587 280909 116588
rect 281030 104141 281090 191251
rect 281027 104140 281093 104141
rect 281027 104076 281028 104140
rect 281092 104076 281093 104140
rect 281027 104075 281093 104076
rect 281582 62797 281642 198867
rect 281766 114341 281826 214643
rect 282131 204916 282197 204917
rect 282131 204852 282132 204916
rect 282196 204852 282197 204916
rect 282131 204851 282197 204852
rect 281947 197844 282013 197845
rect 281947 197780 281948 197844
rect 282012 197780 282013 197844
rect 281947 197779 282013 197780
rect 281950 134741 282010 197779
rect 282134 169829 282194 204851
rect 282131 169828 282197 169829
rect 282131 169764 282132 169828
rect 282196 169764 282197 169828
rect 282131 169763 282197 169764
rect 282870 164661 282930 357443
rect 284339 355060 284405 355061
rect 284339 354996 284340 355060
rect 284404 354996 284405 355060
rect 284339 354995 284405 354996
rect 283051 353972 283117 353973
rect 283051 353908 283052 353972
rect 283116 353908 283117 353972
rect 283051 353907 283117 353908
rect 283054 166293 283114 353907
rect 283235 191860 283301 191861
rect 283235 191796 283236 191860
rect 283300 191796 283301 191860
rect 283235 191795 283301 191796
rect 283051 166292 283117 166293
rect 283051 166228 283052 166292
rect 283116 166228 283117 166292
rect 283051 166227 283117 166228
rect 282867 164660 282933 164661
rect 282867 164596 282868 164660
rect 282932 164596 282933 164660
rect 282867 164595 282933 164596
rect 281947 134740 282013 134741
rect 281947 134676 281948 134740
rect 282012 134676 282013 134740
rect 281947 134675 282013 134676
rect 281763 114340 281829 114341
rect 281763 114276 281764 114340
rect 281828 114276 281829 114340
rect 281763 114275 281829 114276
rect 283238 98837 283298 191795
rect 284342 165749 284402 354995
rect 284523 345676 284589 345677
rect 284523 345612 284524 345676
rect 284588 345612 284589 345676
rect 284523 345611 284589 345612
rect 284526 303381 284586 345611
rect 284523 303380 284589 303381
rect 284523 303316 284524 303380
rect 284588 303316 284589 303380
rect 284523 303315 284589 303316
rect 284523 291412 284589 291413
rect 284523 291348 284524 291412
rect 284588 291348 284589 291412
rect 284523 291347 284589 291348
rect 284339 165748 284405 165749
rect 284339 165684 284340 165748
rect 284404 165684 284405 165748
rect 284339 165683 284405 165684
rect 284526 120053 284586 291347
rect 284894 260133 284954 375123
rect 287835 371244 287901 371245
rect 287835 371180 287836 371244
rect 287900 371180 287901 371244
rect 287835 371179 287901 371180
rect 285811 353564 285877 353565
rect 285811 353500 285812 353564
rect 285876 353500 285877 353564
rect 285811 353499 285877 353500
rect 285627 296852 285693 296853
rect 285627 296788 285628 296852
rect 285692 296788 285693 296852
rect 285627 296787 285693 296788
rect 284891 260132 284957 260133
rect 284891 260068 284892 260132
rect 284956 260068 284957 260132
rect 284891 260067 284957 260068
rect 284707 196756 284773 196757
rect 284707 196692 284708 196756
rect 284772 196692 284773 196756
rect 284707 196691 284773 196692
rect 284523 120052 284589 120053
rect 284523 119988 284524 120052
rect 284588 119988 284589 120052
rect 284523 119987 284589 119988
rect 283235 98836 283301 98837
rect 283235 98772 283236 98836
rect 283300 98772 283301 98836
rect 283235 98771 283301 98772
rect 281579 62796 281645 62797
rect 281579 62732 281580 62796
rect 281644 62732 281645 62796
rect 281579 62731 281645 62732
rect 280659 44980 280725 44981
rect 280659 44916 280660 44980
rect 280724 44916 280725 44980
rect 280659 44915 280725 44916
rect 284710 29749 284770 196691
rect 284891 194036 284957 194037
rect 284891 193972 284892 194036
rect 284956 193972 284957 194036
rect 284891 193971 284957 193972
rect 284894 109717 284954 193971
rect 285630 119781 285690 296787
rect 285814 231573 285874 353499
rect 287651 345540 287717 345541
rect 287651 345476 287652 345540
rect 287716 345476 287717 345540
rect 287651 345475 287717 345476
rect 286915 341188 286981 341189
rect 286915 341124 286916 341188
rect 286980 341124 286981 341188
rect 286915 341123 286981 341124
rect 285995 336700 286061 336701
rect 285995 336636 285996 336700
rect 286060 336636 286061 336700
rect 285995 336635 286061 336636
rect 285998 244085 286058 336635
rect 285995 244084 286061 244085
rect 285995 244020 285996 244084
rect 286060 244020 286061 244084
rect 285995 244019 286061 244020
rect 285811 231572 285877 231573
rect 285811 231508 285812 231572
rect 285876 231508 285877 231572
rect 285811 231507 285877 231508
rect 286918 210085 286978 341123
rect 287283 297940 287349 297941
rect 287283 297876 287284 297940
rect 287348 297876 287349 297940
rect 287283 297875 287349 297876
rect 287099 297396 287165 297397
rect 287099 297332 287100 297396
rect 287164 297332 287165 297396
rect 287099 297331 287165 297332
rect 286915 210084 286981 210085
rect 286915 210020 286916 210084
rect 286980 210020 286981 210084
rect 286915 210019 286981 210020
rect 285811 200020 285877 200021
rect 285811 199956 285812 200020
rect 285876 199956 285877 200020
rect 285811 199955 285877 199956
rect 285627 119780 285693 119781
rect 285627 119716 285628 119780
rect 285692 119716 285693 119780
rect 285627 119715 285693 119716
rect 284891 109716 284957 109717
rect 284891 109652 284892 109716
rect 284956 109652 284957 109716
rect 284891 109651 284957 109652
rect 284707 29748 284773 29749
rect 284707 29684 284708 29748
rect 284772 29684 284773 29748
rect 284707 29683 284773 29684
rect 279834 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 280454 29494
rect 279834 29174 280454 29258
rect 279834 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 280454 29174
rect 279834 -7066 280454 28938
rect 285814 22813 285874 199955
rect 287102 119917 287162 297331
rect 287286 121413 287346 297875
rect 287467 296308 287533 296309
rect 287467 296244 287468 296308
rect 287532 296244 287533 296308
rect 287467 296243 287533 296244
rect 287283 121412 287349 121413
rect 287283 121348 287284 121412
rect 287348 121348 287349 121412
rect 287283 121347 287349 121348
rect 287470 121277 287530 296243
rect 287654 245717 287714 345475
rect 287838 299437 287898 371179
rect 289794 363454 290414 388711
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 288571 347580 288637 347581
rect 288571 347516 288572 347580
rect 288636 347516 288637 347580
rect 288571 347515 288637 347516
rect 288387 345404 288453 345405
rect 288387 345340 288388 345404
rect 288452 345340 288453 345404
rect 288387 345339 288453 345340
rect 287835 299436 287901 299437
rect 287835 299372 287836 299436
rect 287900 299372 287901 299436
rect 287835 299371 287901 299372
rect 287651 245716 287717 245717
rect 287651 245652 287652 245716
rect 287716 245652 287717 245716
rect 287651 245651 287717 245652
rect 288390 239733 288450 345339
rect 288574 249525 288634 347515
rect 289794 327454 290414 362898
rect 293514 367174 294134 388711
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 291331 346764 291397 346765
rect 291331 346700 291332 346764
rect 291396 346700 291397 346764
rect 291331 346699 291397 346700
rect 290779 346220 290845 346221
rect 290779 346156 290780 346220
rect 290844 346156 290845 346220
rect 290779 346155 290845 346156
rect 290595 341052 290661 341053
rect 290595 340988 290596 341052
rect 290660 340988 290661 341052
rect 290595 340987 290661 340988
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 288571 249524 288637 249525
rect 288571 249460 288572 249524
rect 288636 249460 288637 249524
rect 288571 249459 288637 249460
rect 288387 239732 288453 239733
rect 288387 239668 288388 239732
rect 288452 239668 288453 239732
rect 288387 239667 288453 239668
rect 289794 219454 290414 254898
rect 290598 245173 290658 340987
rect 290782 338061 290842 346155
rect 290779 338060 290845 338061
rect 290779 337996 290780 338060
rect 290844 337996 290845 338060
rect 290779 337995 290845 337996
rect 290963 337788 291029 337789
rect 290963 337724 290964 337788
rect 291028 337724 291029 337788
rect 290963 337723 291029 337724
rect 290966 316050 291026 337723
rect 290782 315990 291026 316050
rect 290595 245172 290661 245173
rect 290595 245108 290596 245172
rect 290660 245108 290661 245172
rect 290595 245107 290661 245108
rect 290782 241909 290842 315990
rect 291147 300660 291213 300661
rect 291147 300596 291148 300660
rect 291212 300596 291213 300660
rect 291147 300595 291213 300596
rect 290779 241908 290845 241909
rect 290779 241844 290780 241908
rect 290844 241844 290845 241908
rect 290779 241843 290845 241844
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 290779 188052 290845 188053
rect 290779 187988 290780 188052
rect 290844 187988 290845 188052
rect 290779 187987 290845 187988
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289491 176084 289557 176085
rect 289491 176020 289492 176084
rect 289556 176020 289557 176084
rect 289491 176019 289557 176020
rect 288939 174996 289005 174997
rect 288939 174932 288940 174996
rect 289004 174932 289005 174996
rect 288939 174931 289005 174932
rect 287467 121276 287533 121277
rect 287467 121212 287468 121276
rect 287532 121212 287533 121276
rect 287467 121211 287533 121212
rect 287099 119916 287165 119917
rect 287099 119852 287100 119916
rect 287164 119852 287165 119916
rect 287099 119851 287165 119852
rect 288942 112573 289002 174931
rect 289494 174589 289554 176019
rect 289491 174588 289557 174589
rect 289491 174524 289492 174588
rect 289556 174524 289557 174588
rect 289491 174523 289557 174524
rect 289794 147454 290414 182898
rect 290595 169556 290661 169557
rect 290595 169492 290596 169556
rect 290660 169492 290661 169556
rect 290595 169491 290661 169492
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 288939 112572 289005 112573
rect 288939 112508 288940 112572
rect 289004 112508 289005 112572
rect 288939 112507 289005 112508
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 290598 97613 290658 169491
rect 290782 140045 290842 187987
rect 290779 140044 290845 140045
rect 290779 139980 290780 140044
rect 290844 139980 290845 140044
rect 290779 139979 290845 139980
rect 291150 115293 291210 300595
rect 291334 240277 291394 346699
rect 291515 338604 291581 338605
rect 291515 338540 291516 338604
rect 291580 338540 291581 338604
rect 291515 338539 291581 338540
rect 291331 240276 291397 240277
rect 291331 240212 291332 240276
rect 291396 240212 291397 240276
rect 291331 240211 291397 240212
rect 291518 235381 291578 338539
rect 293514 331174 294134 366618
rect 297234 370894 297854 388711
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 295563 342820 295629 342821
rect 295563 342756 295564 342820
rect 295628 342756 295629 342820
rect 295563 342755 295629 342756
rect 295379 342548 295445 342549
rect 295379 342484 295380 342548
rect 295444 342484 295445 342548
rect 295379 342483 295445 342484
rect 294643 338468 294709 338469
rect 294643 338404 294644 338468
rect 294708 338404 294709 338468
rect 294643 338403 294709 338404
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 292619 300116 292685 300117
rect 292619 300052 292620 300116
rect 292684 300052 292685 300116
rect 292619 300051 292685 300052
rect 291515 235380 291581 235381
rect 291515 235316 291516 235380
rect 291580 235316 291581 235380
rect 291515 235315 291581 235316
rect 291883 185332 291949 185333
rect 291883 185268 291884 185332
rect 291948 185268 291949 185332
rect 291883 185267 291949 185268
rect 291699 171188 291765 171189
rect 291699 171124 291700 171188
rect 291764 171124 291765 171188
rect 291699 171123 291765 171124
rect 291331 169012 291397 169013
rect 291331 168948 291332 169012
rect 291396 168948 291397 169012
rect 291331 168947 291397 168948
rect 291334 116109 291394 168947
rect 291515 131204 291581 131205
rect 291515 131140 291516 131204
rect 291580 131140 291581 131204
rect 291515 131139 291581 131140
rect 291518 119237 291578 131139
rect 291515 119236 291581 119237
rect 291515 119172 291516 119236
rect 291580 119172 291581 119236
rect 291515 119171 291581 119172
rect 291331 116108 291397 116109
rect 291331 116044 291332 116108
rect 291396 116044 291397 116108
rect 291331 116043 291397 116044
rect 291147 115292 291213 115293
rect 291147 115228 291148 115292
rect 291212 115228 291213 115292
rect 291147 115227 291213 115228
rect 291702 103325 291762 171123
rect 291886 131613 291946 185267
rect 291883 131612 291949 131613
rect 291883 131548 291884 131612
rect 291948 131548 291949 131612
rect 291883 131547 291949 131548
rect 292622 120461 292682 300051
rect 293514 295174 294134 330618
rect 294459 301748 294525 301749
rect 294459 301684 294460 301748
rect 294524 301684 294525 301748
rect 294459 301683 294525 301684
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293355 162076 293421 162077
rect 293355 162012 293356 162076
rect 293420 162012 293421 162076
rect 293355 162011 293421 162012
rect 293358 154869 293418 162011
rect 293355 154868 293421 154869
rect 293355 154804 293356 154868
rect 293420 154804 293421 154868
rect 293355 154803 293421 154804
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 292619 120460 292685 120461
rect 292619 120396 292620 120460
rect 292684 120396 292685 120460
rect 292619 120395 292685 120396
rect 291883 118828 291949 118829
rect 291883 118764 291884 118828
rect 291948 118764 291949 118828
rect 291883 118763 291949 118764
rect 291886 112437 291946 118763
rect 293514 115174 294134 150618
rect 294275 125492 294341 125493
rect 294275 125428 294276 125492
rect 294340 125428 294341 125492
rect 294275 125427 294341 125428
rect 294278 119509 294338 125427
rect 294275 119508 294341 119509
rect 294275 119444 294276 119508
rect 294340 119444 294341 119508
rect 294275 119443 294341 119444
rect 294462 118557 294522 301683
rect 294646 231029 294706 338403
rect 295382 234293 295442 342483
rect 295566 239189 295626 342755
rect 296483 340916 296549 340917
rect 296483 340852 296484 340916
rect 296548 340852 296549 340916
rect 296483 340851 296549 340852
rect 295563 239188 295629 239189
rect 295563 239124 295564 239188
rect 295628 239124 295629 239188
rect 295563 239123 295629 239124
rect 296486 238770 296546 340851
rect 296851 339692 296917 339693
rect 296851 339628 296852 339692
rect 296916 339628 296917 339692
rect 296851 339627 296917 339628
rect 296486 238710 296730 238770
rect 296670 238645 296730 238710
rect 296667 238644 296733 238645
rect 296667 238580 296668 238644
rect 296732 238580 296733 238644
rect 296667 238579 296733 238580
rect 296854 238101 296914 339627
rect 297234 334894 297854 370338
rect 300954 374614 301574 388711
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 298139 349212 298205 349213
rect 298139 349148 298140 349212
rect 298204 349148 298205 349212
rect 298139 349147 298205 349148
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 296851 238100 296917 238101
rect 296851 238036 296852 238100
rect 296916 238036 296917 238100
rect 296851 238035 296917 238036
rect 295379 234292 295445 234293
rect 295379 234228 295380 234292
rect 295444 234228 295445 234292
rect 295379 234227 295445 234228
rect 294643 231028 294709 231029
rect 294643 230964 294644 231028
rect 294708 230964 294709 231028
rect 294643 230963 294709 230964
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 294827 182068 294893 182069
rect 294827 182004 294828 182068
rect 294892 182004 294893 182068
rect 294827 182003 294893 182004
rect 294643 177172 294709 177173
rect 294643 177108 294644 177172
rect 294708 177108 294709 177172
rect 294643 177107 294709 177108
rect 294459 118556 294525 118557
rect 294459 118492 294460 118556
rect 294524 118492 294525 118556
rect 294459 118491 294525 118492
rect 294646 115293 294706 177107
rect 294830 125085 294890 182003
rect 296115 178804 296181 178805
rect 296115 178740 296116 178804
rect 296180 178740 296181 178804
rect 296115 178739 296181 178740
rect 295931 173908 295997 173909
rect 295931 173844 295932 173908
rect 295996 173844 295997 173908
rect 295931 173843 295997 173844
rect 294827 125084 294893 125085
rect 294827 125020 294828 125084
rect 294892 125020 294893 125084
rect 294827 125019 294893 125020
rect 294643 115292 294709 115293
rect 294643 115228 294644 115292
rect 294708 115228 294709 115292
rect 294643 115227 294709 115228
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 291883 112436 291949 112437
rect 291883 112372 291884 112436
rect 291948 112372 291949 112436
rect 291883 112371 291949 112372
rect 291699 103324 291765 103325
rect 291699 103260 291700 103324
rect 291764 103260 291765 103324
rect 291699 103259 291765 103260
rect 290595 97612 290661 97613
rect 290595 97548 290596 97612
rect 290660 97548 290661 97612
rect 290595 97547 290661 97548
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 285811 22812 285877 22813
rect 285811 22748 285812 22812
rect 285876 22748 285877 22812
rect 285811 22747 285877 22748
rect 279834 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 280454 -7066
rect 279834 -7386 280454 -7302
rect 279834 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 280454 -7386
rect 279834 -7654 280454 -7622
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -7654 290414 -902
rect 293514 79174 294134 114618
rect 295934 109717 295994 173843
rect 296118 120869 296178 178739
rect 297234 154894 297854 190338
rect 298142 164117 298202 349147
rect 299427 347988 299493 347989
rect 299427 347924 299428 347988
rect 299492 347924 299493 347988
rect 299427 347923 299493 347924
rect 299430 241365 299490 347923
rect 299611 347852 299677 347853
rect 299611 347788 299612 347852
rect 299676 347788 299677 347852
rect 299611 347787 299677 347788
rect 299427 241364 299493 241365
rect 299427 241300 299428 241364
rect 299492 241300 299493 241364
rect 299427 241299 299493 241300
rect 299614 240821 299674 347787
rect 300954 338614 301574 374058
rect 304674 378334 305294 388711
rect 304674 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 305294 378334
rect 304674 378014 305294 378098
rect 304674 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 305294 378014
rect 303659 343908 303725 343909
rect 303659 343844 303660 343908
rect 303724 343844 303725 343908
rect 303659 343843 303725 343844
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 301819 338196 301885 338197
rect 301819 338132 301820 338196
rect 301884 338132 301885 338196
rect 301819 338131 301885 338132
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 299611 240820 299677 240821
rect 299611 240756 299612 240820
rect 299676 240756 299677 240820
rect 299611 240755 299677 240756
rect 300954 230614 301574 266058
rect 301822 233205 301882 338131
rect 303662 234837 303722 343843
rect 304674 342334 305294 377778
rect 308394 382054 309014 388711
rect 308394 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 309014 382054
rect 308394 381734 309014 381818
rect 308394 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 309014 381734
rect 308394 346054 309014 381498
rect 308394 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 309014 346054
rect 308394 345734 309014 345818
rect 308394 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 309014 345734
rect 306419 344860 306485 344861
rect 306419 344796 306420 344860
rect 306484 344796 306485 344860
rect 306419 344795 306485 344796
rect 304674 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 305294 342334
rect 304674 342014 305294 342098
rect 304674 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 305294 342014
rect 303843 339012 303909 339013
rect 303843 338948 303844 339012
rect 303908 338948 303909 339012
rect 303843 338947 303909 338948
rect 303659 234836 303725 234837
rect 303659 234772 303660 234836
rect 303724 234772 303725 234836
rect 303659 234771 303725 234772
rect 301819 233204 301885 233205
rect 301819 233140 301820 233204
rect 301884 233140 301885 233204
rect 301819 233139 301885 233140
rect 303846 232117 303906 338947
rect 304674 306334 305294 341778
rect 304674 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 305294 306334
rect 304674 306014 305294 306098
rect 304674 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 305294 306014
rect 304674 270334 305294 305778
rect 304674 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 305294 270334
rect 304674 270014 305294 270098
rect 304674 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 305294 270014
rect 304674 234334 305294 269778
rect 304674 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 305294 234334
rect 304674 234014 305294 234098
rect 304674 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 305294 234014
rect 303843 232116 303909 232117
rect 303843 232052 303844 232116
rect 303908 232052 303909 232116
rect 303843 232051 303909 232052
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300163 186420 300229 186421
rect 300163 186356 300164 186420
rect 300228 186356 300229 186420
rect 300163 186355 300229 186356
rect 298875 184244 298941 184245
rect 298875 184180 298876 184244
rect 298940 184180 298941 184244
rect 298875 184179 298941 184180
rect 298139 164116 298205 164117
rect 298139 164052 298140 164116
rect 298204 164052 298205 164116
rect 298139 164051 298205 164052
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 296115 120868 296181 120869
rect 296115 120804 296116 120868
rect 296180 120804 296181 120868
rect 296115 120803 296181 120804
rect 297234 118894 297854 154338
rect 298691 150516 298757 150517
rect 298691 150452 298692 150516
rect 298756 150452 298757 150516
rect 298691 150451 298757 150452
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 295931 109716 295997 109717
rect 295931 109652 295932 109716
rect 295996 109652 295997 109716
rect 295931 109651 295997 109652
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -1306 294134 6618
rect 293514 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 294134 -1306
rect 293514 -1626 294134 -1542
rect 293514 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 294134 -1626
rect 293514 -7654 294134 -1862
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 298694 19821 298754 150451
rect 298878 129437 298938 184179
rect 299979 176628 300045 176629
rect 299979 176564 299980 176628
rect 300044 176564 300045 176628
rect 299979 176563 300045 176564
rect 298875 129436 298941 129437
rect 298875 129372 298876 129436
rect 298940 129372 298941 129436
rect 298875 129371 298941 129372
rect 299982 114205 300042 176563
rect 300166 133789 300226 186355
rect 300954 158614 301574 194058
rect 304674 198334 305294 233778
rect 306422 230485 306482 344795
rect 308394 310054 309014 345498
rect 308394 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 309014 310054
rect 308394 309734 309014 309818
rect 308394 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 309014 309734
rect 308394 274054 309014 309498
rect 308394 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 309014 274054
rect 308394 273734 309014 273818
rect 308394 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 309014 273734
rect 308394 238054 309014 273498
rect 308394 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 309014 238054
rect 308394 237734 309014 237818
rect 308394 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 309014 237734
rect 306419 230484 306485 230485
rect 306419 230420 306420 230484
rect 306484 230420 306485 230484
rect 306419 230419 306485 230420
rect 304674 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 305294 198334
rect 304674 198014 305294 198098
rect 304674 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 305294 198014
rect 302923 190228 302989 190229
rect 302923 190164 302924 190228
rect 302988 190164 302989 190228
rect 302923 190163 302989 190164
rect 302739 177716 302805 177717
rect 302739 177652 302740 177716
rect 302804 177652 302805 177716
rect 302739 177651 302805 177652
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300163 133788 300229 133789
rect 300163 133724 300164 133788
rect 300228 133724 300229 133788
rect 300163 133723 300229 133724
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 299979 114204 300045 114205
rect 299979 114140 299980 114204
rect 300044 114140 300045 114204
rect 299979 114139 300045 114140
rect 300954 86614 301574 122058
rect 302742 116381 302802 177651
rect 302926 142765 302986 190163
rect 304211 173364 304277 173365
rect 304211 173300 304212 173364
rect 304276 173300 304277 173364
rect 304211 173299 304277 173300
rect 302923 142764 302989 142765
rect 302923 142700 302924 142764
rect 302988 142700 302989 142764
rect 302923 142699 302989 142700
rect 302739 116380 302805 116381
rect 302739 116316 302740 116380
rect 302804 116316 302805 116380
rect 302739 116315 302805 116316
rect 304214 107677 304274 173299
rect 304674 162334 305294 197778
rect 308394 202054 309014 237498
rect 308394 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 309014 202054
rect 308394 201734 309014 201818
rect 308394 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 309014 201734
rect 307155 181524 307221 181525
rect 307155 181460 307156 181524
rect 307220 181460 307221 181524
rect 307155 181459 307221 181460
rect 305499 174452 305565 174453
rect 305499 174388 305500 174452
rect 305564 174388 305565 174452
rect 305499 174387 305565 174388
rect 304674 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 305294 162334
rect 304674 162014 305294 162098
rect 304674 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 305294 162014
rect 304674 126334 305294 161778
rect 304674 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 305294 126334
rect 304674 126014 305294 126098
rect 304674 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 305294 126014
rect 304211 107676 304277 107677
rect 304211 107612 304212 107676
rect 304276 107612 304277 107676
rect 304211 107611 304277 107612
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 298691 19820 298757 19821
rect 298691 19756 298692 19820
rect 298756 19756 298757 19820
rect 298691 19755 298757 19756
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -2266 297854 10338
rect 297234 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 297854 -2266
rect 297234 -2586 297854 -2502
rect 297234 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 297854 -2586
rect 297234 -7654 297854 -2822
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 300954 -3226 301574 14058
rect 300954 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 301574 -3226
rect 300954 -3546 301574 -3462
rect 300954 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 301574 -3546
rect 300954 -7654 301574 -3782
rect 304674 90334 305294 125778
rect 305502 111077 305562 174387
rect 306419 152148 306485 152149
rect 306419 152084 306420 152148
rect 306484 152084 306485 152148
rect 306419 152083 306485 152084
rect 306422 151061 306482 152083
rect 306419 151060 306485 151061
rect 306419 150996 306420 151060
rect 306484 150996 306485 151060
rect 306419 150995 306485 150996
rect 306971 150924 307037 150925
rect 306971 150860 306972 150924
rect 307036 150860 307037 150924
rect 306971 150859 307037 150860
rect 305499 111076 305565 111077
rect 305499 111012 305500 111076
rect 305564 111012 305565 111076
rect 305499 111011 305565 111012
rect 304674 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 305294 90334
rect 304674 90014 305294 90098
rect 304674 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 305294 90014
rect 304674 54334 305294 89778
rect 306974 59669 307034 150859
rect 307158 123997 307218 181459
rect 308394 166054 309014 201498
rect 312114 385774 312734 388711
rect 312114 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 312734 385774
rect 312114 385454 312734 385538
rect 312114 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 312734 385454
rect 312114 349774 312734 385218
rect 312114 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 312734 349774
rect 312114 349454 312734 349538
rect 312114 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 312734 349454
rect 312114 313774 312734 349218
rect 312114 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 312734 313774
rect 312114 313454 312734 313538
rect 312114 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 312734 313454
rect 312114 277774 312734 313218
rect 312114 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 312734 277774
rect 312114 277454 312734 277538
rect 312114 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 312734 277454
rect 312114 241774 312734 277218
rect 312114 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 312734 241774
rect 312114 241454 312734 241538
rect 312114 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 312734 241454
rect 312114 205774 312734 241218
rect 312114 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 312734 205774
rect 312114 205454 312734 205538
rect 312114 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 312734 205454
rect 309731 180436 309797 180437
rect 309731 180372 309732 180436
rect 309796 180372 309797 180436
rect 309731 180371 309797 180372
rect 308394 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 309014 166054
rect 308394 165734 309014 165818
rect 308394 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 309014 165734
rect 308394 130054 309014 165498
rect 308394 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 309014 130054
rect 308394 129734 309014 129818
rect 308394 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 309014 129734
rect 307155 123996 307221 123997
rect 307155 123932 307156 123996
rect 307220 123932 307221 123996
rect 307155 123931 307221 123932
rect 308394 94054 309014 129498
rect 309734 121821 309794 180371
rect 311019 171732 311085 171733
rect 311019 171668 311020 171732
rect 311084 171668 311085 171732
rect 311019 171667 311085 171668
rect 309731 121820 309797 121821
rect 309731 121756 309732 121820
rect 309796 121756 309797 121820
rect 309731 121755 309797 121756
rect 311022 104413 311082 171667
rect 312114 169774 312734 205218
rect 315834 353494 316454 388711
rect 315834 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 316454 353494
rect 315834 353174 316454 353258
rect 315834 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 316454 353174
rect 315834 317494 316454 352938
rect 315834 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 316454 317494
rect 315834 317174 316454 317258
rect 315834 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 316454 317174
rect 315834 281494 316454 316938
rect 315834 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 316454 281494
rect 315834 281174 316454 281258
rect 315834 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 316454 281174
rect 315834 245494 316454 280938
rect 315834 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 316454 245494
rect 315834 245174 316454 245258
rect 315834 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 316454 245174
rect 315834 209494 316454 244938
rect 315834 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 316454 209494
rect 315834 209174 316454 209258
rect 315834 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 316454 209174
rect 313963 187508 314029 187509
rect 313963 187444 313964 187508
rect 314028 187444 314029 187508
rect 313963 187443 314029 187444
rect 312114 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 312734 169774
rect 312114 169454 312734 169538
rect 312114 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 312734 169454
rect 312114 133774 312734 169218
rect 313779 151604 313845 151605
rect 313779 151540 313780 151604
rect 313844 151540 313845 151604
rect 313779 151539 313845 151540
rect 312114 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 312734 133774
rect 312114 133454 312734 133538
rect 312114 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 312734 133454
rect 311019 104412 311085 104413
rect 311019 104348 311020 104412
rect 311084 104348 311085 104412
rect 311019 104347 311085 104348
rect 308394 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 309014 94054
rect 308394 93734 309014 93818
rect 308394 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 309014 93734
rect 306971 59668 307037 59669
rect 306971 59604 306972 59668
rect 307036 59604 307037 59668
rect 306971 59603 307037 59604
rect 304674 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 305294 54334
rect 304674 54014 305294 54098
rect 304674 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 305294 54014
rect 304674 18334 305294 53778
rect 304674 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 305294 18334
rect 304674 18014 305294 18098
rect 304674 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 305294 18014
rect 304674 -4186 305294 17778
rect 304674 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 305294 -4186
rect 304674 -4506 305294 -4422
rect 304674 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 305294 -4506
rect 304674 -7654 305294 -4742
rect 308394 58054 309014 93498
rect 308394 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 309014 58054
rect 308394 57734 309014 57818
rect 308394 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 309014 57734
rect 308394 22054 309014 57498
rect 308394 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 309014 22054
rect 308394 21734 309014 21818
rect 308394 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 309014 21734
rect 308394 -5146 309014 21498
rect 308394 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 309014 -5146
rect 308394 -5466 309014 -5382
rect 308394 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 309014 -5466
rect 308394 -7654 309014 -5702
rect 312114 97774 312734 133218
rect 313782 99517 313842 151539
rect 313966 135965 314026 187443
rect 315834 173494 316454 208938
rect 325794 363454 326414 388711
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 319299 184788 319365 184789
rect 319299 184724 319300 184788
rect 319364 184724 319365 184788
rect 319299 184723 319365 184724
rect 315834 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 316454 173494
rect 315834 173174 316454 173258
rect 315834 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 316454 173174
rect 315834 137494 316454 172938
rect 315834 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 316454 137494
rect 315834 137174 316454 137258
rect 315834 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 316454 137174
rect 313963 135964 314029 135965
rect 313963 135900 313964 135964
rect 314028 135900 314029 135964
rect 313963 135899 314029 135900
rect 315834 101494 316454 136938
rect 319302 130525 319362 184723
rect 325794 183454 326414 218898
rect 329514 367174 330134 388711
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 327763 188596 327829 188597
rect 327763 188532 327764 188596
rect 327828 188532 327829 188596
rect 327763 188531 327829 188532
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 322059 172820 322125 172821
rect 322059 172756 322060 172820
rect 322124 172756 322125 172820
rect 322059 172755 322125 172756
rect 319299 130524 319365 130525
rect 319299 130460 319300 130524
rect 319364 130460 319365 130524
rect 319299 130459 319365 130460
rect 322062 106589 322122 172755
rect 323531 172276 323597 172277
rect 323531 172212 323532 172276
rect 323596 172212 323597 172276
rect 323531 172211 323597 172212
rect 322059 106588 322125 106589
rect 322059 106524 322060 106588
rect 322124 106524 322125 106588
rect 322059 106523 322125 106524
rect 323534 105501 323594 172211
rect 325794 147454 326414 182898
rect 327579 178260 327645 178261
rect 327579 178196 327580 178260
rect 327644 178196 327645 178260
rect 327579 178195 327645 178196
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 327582 119373 327642 178195
rect 327766 141405 327826 188531
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 327763 141404 327829 141405
rect 327763 141340 327764 141404
rect 327828 141340 327829 141404
rect 327763 141339 327829 141340
rect 327579 119372 327645 119373
rect 327579 119308 327580 119372
rect 327644 119308 327645 119372
rect 327579 119307 327645 119308
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 323531 105500 323597 105501
rect 323531 105436 323532 105500
rect 323596 105436 323597 105500
rect 323531 105435 323597 105436
rect 315834 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 316454 101494
rect 315834 101174 316454 101258
rect 315834 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 316454 101174
rect 313779 99516 313845 99517
rect 313779 99452 313780 99516
rect 313844 99452 313845 99516
rect 313779 99451 313845 99452
rect 312114 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 312734 97774
rect 312114 97454 312734 97538
rect 312114 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 312734 97454
rect 312114 61774 312734 97218
rect 312114 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 312734 61774
rect 312114 61454 312734 61538
rect 312114 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 312734 61454
rect 312114 25774 312734 61218
rect 312114 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 312734 25774
rect 312114 25454 312734 25538
rect 312114 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 312734 25454
rect 312114 -6106 312734 25218
rect 312114 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 312734 -6106
rect 312114 -6426 312734 -6342
rect 312114 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 312734 -6426
rect 312114 -7654 312734 -6662
rect 315834 65494 316454 100938
rect 315834 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 316454 65494
rect 315834 65174 316454 65258
rect 315834 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 316454 65174
rect 315834 29494 316454 64938
rect 315834 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 316454 29494
rect 315834 29174 316454 29258
rect 315834 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 316454 29174
rect 315834 -7066 316454 28938
rect 315834 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 316454 -7066
rect 315834 -7386 316454 -7302
rect 315834 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 316454 -7386
rect 315834 -7654 316454 -7622
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -7654 326414 -902
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -1306 330134 6618
rect 329514 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 330134 -1306
rect 329514 -1626 330134 -1542
rect 329514 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 330134 -1626
rect 329514 -7654 330134 -1862
rect 333234 370894 333854 388711
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 336954 374614 337574 388711
rect 338619 381852 338685 381853
rect 338619 381788 338620 381852
rect 338684 381788 338685 381852
rect 338619 381787 338685 381788
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 338622 278357 338682 381787
rect 340674 378334 341294 388711
rect 340674 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 341294 378334
rect 340674 378014 341294 378098
rect 340674 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 341294 378014
rect 340674 342334 341294 377778
rect 340674 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 341294 342334
rect 340674 342014 341294 342098
rect 340674 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 341294 342014
rect 340674 306334 341294 341778
rect 340674 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 341294 306334
rect 340674 306014 341294 306098
rect 340674 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 341294 306014
rect 338619 278356 338685 278357
rect 338619 278292 338620 278356
rect 338684 278292 338685 278356
rect 338619 278291 338685 278292
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 334571 185876 334637 185877
rect 334571 185812 334572 185876
rect 334636 185812 334637 185876
rect 334571 185811 334637 185812
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 334574 134469 334634 185811
rect 335859 182612 335925 182613
rect 335859 182548 335860 182612
rect 335924 182548 335925 182612
rect 335859 182547 335925 182548
rect 334755 179212 334821 179213
rect 334755 179148 334756 179212
rect 334820 179148 334821 179212
rect 334755 179147 334821 179148
rect 334758 152693 334818 179147
rect 334755 152692 334821 152693
rect 334755 152628 334756 152692
rect 334820 152628 334821 152692
rect 334755 152627 334821 152628
rect 334571 134468 334637 134469
rect 334571 134404 334572 134468
rect 334636 134404 334637 134468
rect 334571 134403 334637 134404
rect 335862 126173 335922 182547
rect 336954 158614 337574 194058
rect 340674 270334 341294 305778
rect 340674 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 341294 270334
rect 340674 270014 341294 270098
rect 340674 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 341294 270014
rect 340674 234334 341294 269778
rect 340674 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 341294 234334
rect 340674 234014 341294 234098
rect 340674 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 341294 234014
rect 340674 198334 341294 233778
rect 340674 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 341294 198334
rect 340674 198014 341294 198098
rect 340674 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 341294 198014
rect 338619 186964 338685 186965
rect 338619 186900 338620 186964
rect 338684 186900 338685 186964
rect 338619 186899 338685 186900
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 335859 126172 335925 126173
rect 335859 126108 335860 126172
rect 335924 126108 335925 126172
rect 335859 126107 335925 126108
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -2266 333854 10338
rect 333234 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 333854 -2266
rect 333234 -2586 333854 -2502
rect 333234 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 333854 -2586
rect 333234 -7654 333854 -2822
rect 336954 122614 337574 158058
rect 338622 137325 338682 186899
rect 340674 162334 341294 197778
rect 344394 382054 345014 388711
rect 345611 388652 345677 388653
rect 345611 388588 345612 388652
rect 345676 388588 345677 388652
rect 345611 388587 345677 388588
rect 344394 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 345014 382054
rect 344394 381734 345014 381818
rect 344394 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 345014 381734
rect 344394 346054 345014 381498
rect 344394 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 345014 346054
rect 344394 345734 345014 345818
rect 344394 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 345014 345734
rect 344394 310054 345014 345498
rect 344394 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 345014 310054
rect 344394 309734 345014 309818
rect 344394 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 345014 309734
rect 344394 274054 345014 309498
rect 344394 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 345014 274054
rect 344394 273734 345014 273818
rect 344394 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 345014 273734
rect 344394 238054 345014 273498
rect 345614 270197 345674 388587
rect 348114 385774 348734 388711
rect 349659 387972 349725 387973
rect 349659 387908 349660 387972
rect 349724 387908 349725 387972
rect 349659 387907 349725 387908
rect 348114 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 348734 385774
rect 348114 385454 348734 385538
rect 348114 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 348734 385454
rect 346899 384572 346965 384573
rect 346899 384508 346900 384572
rect 346964 384508 346965 384572
rect 346899 384507 346965 384508
rect 346902 276181 346962 384507
rect 348114 349774 348734 385218
rect 348114 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 348734 349774
rect 348114 349454 348734 349538
rect 348114 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 348734 349454
rect 348114 313774 348734 349218
rect 348114 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 348734 313774
rect 348114 313454 348734 313538
rect 348114 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 348734 313454
rect 348114 277774 348734 313218
rect 348114 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 348734 277774
rect 348114 277454 348734 277538
rect 348114 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 348734 277454
rect 346899 276180 346965 276181
rect 346899 276116 346900 276180
rect 346964 276116 346965 276180
rect 346899 276115 346965 276116
rect 345611 270196 345677 270197
rect 345611 270132 345612 270196
rect 345676 270132 345677 270196
rect 345611 270131 345677 270132
rect 344394 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 345014 238054
rect 344394 237734 345014 237818
rect 344394 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 345014 237734
rect 344394 202054 345014 237498
rect 344394 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 345014 202054
rect 344394 201734 345014 201818
rect 344394 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 345014 201734
rect 342851 183700 342917 183701
rect 342851 183636 342852 183700
rect 342916 183636 342917 183700
rect 342851 183635 342917 183636
rect 340674 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 341294 162334
rect 340674 162014 341294 162098
rect 340674 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 341294 162014
rect 338619 137324 338685 137325
rect 338619 137260 338620 137324
rect 338684 137260 338685 137324
rect 338619 137259 338685 137260
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 336954 -3226 337574 14058
rect 336954 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 337574 -3226
rect 336954 -3546 337574 -3462
rect 336954 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 337574 -3546
rect 336954 -7654 337574 -3782
rect 340674 126334 341294 161778
rect 342854 128349 342914 183635
rect 344394 166054 345014 201498
rect 348114 241774 348734 277218
rect 349662 275637 349722 387907
rect 349843 385796 349909 385797
rect 349843 385732 349844 385796
rect 349908 385732 349909 385796
rect 349843 385731 349909 385732
rect 349846 281077 349906 385731
rect 351131 384708 351197 384709
rect 351131 384644 351132 384708
rect 351196 384644 351197 384708
rect 351131 384643 351197 384644
rect 349843 281076 349909 281077
rect 349843 281012 349844 281076
rect 349908 281012 349909 281076
rect 349843 281011 349909 281012
rect 351134 276725 351194 384643
rect 351315 372060 351381 372061
rect 351315 371996 351316 372060
rect 351380 371996 351381 372060
rect 351315 371995 351381 371996
rect 351131 276724 351197 276725
rect 351131 276660 351132 276724
rect 351196 276660 351197 276724
rect 351131 276659 351197 276660
rect 349659 275636 349725 275637
rect 349659 275572 349660 275636
rect 349724 275572 349725 275636
rect 349659 275571 349725 275572
rect 351318 275093 351378 371995
rect 351834 353494 352454 388711
rect 356651 384844 356717 384845
rect 356651 384780 356652 384844
rect 356716 384780 356717 384844
rect 356651 384779 356717 384780
rect 354627 384028 354693 384029
rect 354627 383964 354628 384028
rect 354692 383964 354693 384028
rect 354627 383963 354693 383964
rect 353891 383892 353957 383893
rect 353891 383828 353892 383892
rect 353956 383828 353957 383892
rect 353891 383827 353957 383828
rect 352971 379268 353037 379269
rect 352971 379204 352972 379268
rect 353036 379204 353037 379268
rect 352971 379203 353037 379204
rect 352787 367708 352853 367709
rect 352787 367644 352788 367708
rect 352852 367644 352853 367708
rect 352787 367643 352853 367644
rect 351834 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 352454 353494
rect 351834 353174 352454 353258
rect 351834 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 352454 353174
rect 351834 317494 352454 352938
rect 351834 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 352454 317494
rect 351834 317174 352454 317258
rect 351834 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 352454 317174
rect 351834 281494 352454 316938
rect 351834 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 352454 281494
rect 351834 281174 352454 281258
rect 351834 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 352454 281174
rect 351315 275092 351381 275093
rect 351315 275028 351316 275092
rect 351380 275028 351381 275092
rect 351315 275027 351381 275028
rect 348114 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 348734 241774
rect 348114 241454 348734 241538
rect 348114 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 348734 241454
rect 348114 205774 348734 241218
rect 348114 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 348734 205774
rect 348114 205454 348734 205538
rect 348114 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 348734 205454
rect 346899 189684 346965 189685
rect 346899 189620 346900 189684
rect 346964 189620 346965 189684
rect 346899 189619 346965 189620
rect 345611 189140 345677 189141
rect 345611 189076 345612 189140
rect 345676 189076 345677 189140
rect 345611 189075 345677 189076
rect 344394 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 345014 166054
rect 344394 165734 345014 165818
rect 344394 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 345014 165734
rect 344394 130054 345014 165498
rect 345614 139229 345674 189075
rect 346902 140317 346962 189619
rect 348114 169774 348734 205218
rect 351834 245494 352454 280938
rect 352790 274005 352850 367643
rect 352974 288149 353034 379203
rect 352971 288148 353037 288149
rect 352971 288084 352972 288148
rect 353036 288084 353037 288148
rect 352971 288083 353037 288084
rect 353894 279445 353954 383827
rect 354630 383670 354690 383963
rect 354446 383610 354690 383670
rect 354075 376548 354141 376549
rect 354075 376484 354076 376548
rect 354140 376484 354141 376548
rect 354075 376483 354141 376484
rect 354078 288693 354138 376483
rect 354259 365260 354325 365261
rect 354259 365196 354260 365260
rect 354324 365196 354325 365260
rect 354259 365195 354325 365196
rect 354075 288692 354141 288693
rect 354075 288628 354076 288692
rect 354140 288628 354141 288692
rect 354075 288627 354141 288628
rect 354262 284341 354322 365195
rect 354259 284340 354325 284341
rect 354259 284276 354260 284340
rect 354324 284276 354325 284340
rect 354259 284275 354325 284276
rect 354446 280669 354506 383610
rect 355179 381988 355245 381989
rect 355179 381924 355180 381988
rect 355244 381924 355245 381988
rect 355179 381923 355245 381924
rect 355182 285973 355242 381923
rect 355547 379404 355613 379405
rect 355547 379340 355548 379404
rect 355612 379340 355613 379404
rect 355547 379339 355613 379340
rect 355363 363628 355429 363629
rect 355363 363564 355364 363628
rect 355428 363564 355429 363628
rect 355363 363563 355429 363564
rect 355179 285972 355245 285973
rect 355179 285908 355180 285972
rect 355244 285908 355245 285972
rect 355179 285907 355245 285908
rect 354443 280668 354509 280669
rect 354443 280604 354444 280668
rect 354508 280604 354509 280668
rect 354443 280603 354509 280604
rect 353891 279444 353957 279445
rect 353891 279380 353892 279444
rect 353956 279380 353957 279444
rect 353891 279379 353957 279380
rect 352787 274004 352853 274005
rect 352787 273940 352788 274004
rect 352852 273940 352853 274004
rect 352787 273939 352853 273940
rect 355366 271829 355426 363563
rect 355550 287605 355610 379339
rect 355547 287604 355613 287605
rect 355547 287540 355548 287604
rect 355612 287540 355613 287604
rect 355547 287539 355613 287540
rect 356654 277269 356714 384779
rect 356835 382260 356901 382261
rect 356835 382196 356836 382260
rect 356900 382196 356901 382260
rect 356835 382195 356901 382196
rect 356838 283253 356898 382195
rect 357203 375460 357269 375461
rect 357203 375396 357204 375460
rect 357268 375396 357269 375460
rect 357203 375395 357269 375396
rect 357019 365396 357085 365397
rect 357019 365332 357020 365396
rect 357084 365332 357085 365396
rect 357019 365331 357085 365332
rect 356835 283252 356901 283253
rect 356835 283188 356836 283252
rect 356900 283188 356901 283252
rect 356835 283187 356901 283188
rect 356651 277268 356717 277269
rect 356651 277204 356652 277268
rect 356716 277204 356717 277268
rect 356651 277203 356717 277204
rect 357022 272917 357082 365331
rect 357206 289237 357266 375395
rect 357203 289236 357269 289237
rect 357203 289172 357204 289236
rect 357268 289172 357269 289236
rect 357203 289171 357269 289172
rect 357019 272916 357085 272917
rect 357019 272852 357020 272916
rect 357084 272852 357085 272916
rect 357019 272851 357085 272852
rect 355363 271828 355429 271829
rect 355363 271764 355364 271828
rect 355428 271764 355429 271828
rect 355363 271763 355429 271764
rect 357942 271285 358002 390219
rect 361619 386884 361685 386885
rect 361619 386820 361620 386884
rect 361684 386820 361685 386884
rect 361619 386819 361685 386820
rect 362907 386884 362973 386885
rect 362907 386820 362908 386884
rect 362972 386820 362973 386884
rect 362907 386819 362973 386820
rect 360147 386748 360213 386749
rect 360147 386684 360148 386748
rect 360212 386684 360213 386748
rect 360147 386683 360213 386684
rect 358123 383076 358189 383077
rect 358123 383012 358124 383076
rect 358188 383012 358189 383076
rect 358123 383011 358189 383012
rect 358126 282165 358186 383011
rect 360150 345813 360210 386683
rect 360331 386476 360397 386477
rect 360331 386412 360332 386476
rect 360396 386412 360397 386476
rect 360331 386411 360397 386412
rect 360147 345812 360213 345813
rect 360147 345748 360148 345812
rect 360212 345748 360213 345812
rect 360147 345747 360213 345748
rect 358123 282164 358189 282165
rect 358123 282100 358124 282164
rect 358188 282100 358189 282164
rect 358123 282099 358189 282100
rect 357939 271284 358005 271285
rect 357939 271220 357940 271284
rect 358004 271220 358005 271284
rect 357939 271219 358005 271220
rect 351834 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 352454 245494
rect 351834 245174 352454 245258
rect 351834 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 352454 245174
rect 351834 209494 352454 244938
rect 351834 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 352454 209494
rect 351834 209174 352454 209258
rect 351834 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 352454 209174
rect 349659 183156 349725 183157
rect 349659 183092 349660 183156
rect 349724 183092 349725 183156
rect 349659 183091 349725 183092
rect 348114 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 348734 169774
rect 348114 169454 348734 169538
rect 348114 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 348734 169454
rect 346899 140316 346965 140317
rect 346899 140252 346900 140316
rect 346964 140252 346965 140316
rect 346899 140251 346965 140252
rect 345611 139228 345677 139229
rect 345611 139164 345612 139228
rect 345676 139164 345677 139228
rect 345611 139163 345677 139164
rect 344394 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 345014 130054
rect 344394 129734 345014 129818
rect 344394 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 345014 129734
rect 342851 128348 342917 128349
rect 342851 128284 342852 128348
rect 342916 128284 342917 128348
rect 342851 128283 342917 128284
rect 340674 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 341294 126334
rect 340674 126014 341294 126098
rect 340674 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 341294 126014
rect 340674 90334 341294 125778
rect 340674 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 341294 90334
rect 340674 90014 341294 90098
rect 340674 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 341294 90014
rect 340674 54334 341294 89778
rect 340674 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 341294 54334
rect 340674 54014 341294 54098
rect 340674 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 341294 54014
rect 340674 18334 341294 53778
rect 340674 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 341294 18334
rect 340674 18014 341294 18098
rect 340674 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 341294 18014
rect 340674 -4186 341294 17778
rect 340674 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 341294 -4186
rect 340674 -4506 341294 -4422
rect 340674 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 341294 -4506
rect 340674 -7654 341294 -4742
rect 344394 94054 345014 129498
rect 344394 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 345014 94054
rect 344394 93734 345014 93818
rect 344394 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 345014 93734
rect 344394 58054 345014 93498
rect 344394 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 345014 58054
rect 344394 57734 345014 57818
rect 344394 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 345014 57734
rect 344394 22054 345014 57498
rect 344394 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 345014 22054
rect 344394 21734 345014 21818
rect 344394 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 345014 21734
rect 344394 -5146 345014 21498
rect 344394 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 345014 -5146
rect 344394 -5466 345014 -5382
rect 344394 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 345014 -5466
rect 344394 -7654 345014 -5702
rect 348114 133774 348734 169218
rect 348114 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 348734 133774
rect 348114 133454 348734 133538
rect 348114 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 348734 133454
rect 348114 97774 348734 133218
rect 349662 127261 349722 183091
rect 351131 179892 351197 179893
rect 351131 179828 351132 179892
rect 351196 179828 351197 179892
rect 351131 179827 351197 179828
rect 349659 127260 349725 127261
rect 349659 127196 349660 127260
rect 349724 127196 349725 127260
rect 349659 127195 349725 127196
rect 351134 120733 351194 179827
rect 351834 173494 352454 208938
rect 353891 180980 353957 180981
rect 353891 180916 353892 180980
rect 353956 180916 353957 180980
rect 353891 180915 353957 180916
rect 351834 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 352454 173494
rect 351834 173174 352454 173258
rect 351834 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 352454 173174
rect 351834 137494 352454 172938
rect 351834 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 352454 137494
rect 351834 137174 352454 137258
rect 351834 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 352454 137174
rect 351131 120732 351197 120733
rect 351131 120668 351132 120732
rect 351196 120668 351197 120732
rect 351131 120667 351197 120668
rect 348114 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 348734 97774
rect 348114 97454 348734 97538
rect 348114 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 348734 97454
rect 348114 61774 348734 97218
rect 348114 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 348734 61774
rect 348114 61454 348734 61538
rect 348114 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 348734 61454
rect 348114 25774 348734 61218
rect 348114 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 348734 25774
rect 348114 25454 348734 25538
rect 348114 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 348734 25454
rect 348114 -6106 348734 25218
rect 348114 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 348734 -6106
rect 348114 -6426 348734 -6342
rect 348114 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 348734 -6426
rect 348114 -7654 348734 -6662
rect 351834 101494 352454 136938
rect 353894 122909 353954 180915
rect 355179 178668 355245 178669
rect 355179 178604 355180 178668
rect 355244 178604 355245 178668
rect 355179 178603 355245 178604
rect 353891 122908 353957 122909
rect 353891 122844 353892 122908
rect 353956 122844 353957 122908
rect 353891 122843 353957 122844
rect 355182 119645 355242 178603
rect 356651 175540 356717 175541
rect 356651 175476 356652 175540
rect 356716 175476 356717 175540
rect 356651 175475 356717 175476
rect 355179 119644 355245 119645
rect 355179 119580 355180 119644
rect 355244 119580 355245 119644
rect 355179 119579 355245 119580
rect 356654 112709 356714 175475
rect 357939 174588 358005 174589
rect 357939 174524 357940 174588
rect 358004 174524 358005 174588
rect 357939 174523 358005 174524
rect 357387 141404 357453 141405
rect 357387 141340 357388 141404
rect 357452 141340 357453 141404
rect 357387 141339 357453 141340
rect 357390 138141 357450 141339
rect 357571 140044 357637 140045
rect 357571 139980 357572 140044
rect 357636 139980 357637 140044
rect 357571 139979 357637 139980
rect 357387 138140 357453 138141
rect 357387 138076 357388 138140
rect 357452 138076 357453 138140
rect 357387 138075 357453 138076
rect 357387 137324 357453 137325
rect 357387 137260 357388 137324
rect 357452 137260 357453 137324
rect 357387 137259 357453 137260
rect 357390 134877 357450 137259
rect 357574 137053 357634 139979
rect 357571 137052 357637 137053
rect 357571 136988 357572 137052
rect 357636 136988 357637 137052
rect 357571 136987 357637 136988
rect 357387 134876 357453 134877
rect 357387 134812 357388 134876
rect 357452 134812 357453 134876
rect 357387 134811 357453 134812
rect 357387 134468 357453 134469
rect 357387 134404 357388 134468
rect 357452 134404 357453 134468
rect 357387 134403 357453 134404
rect 357390 132701 357450 134403
rect 357387 132700 357453 132701
rect 357387 132636 357388 132700
rect 357452 132636 357453 132700
rect 357387 132635 357453 132636
rect 357571 120868 357637 120869
rect 357571 120804 357572 120868
rect 357636 120804 357637 120868
rect 357571 120803 357637 120804
rect 357387 119372 357453 119373
rect 357387 119308 357388 119372
rect 357452 119308 357453 119372
rect 357387 119307 357453 119308
rect 357390 117469 357450 119307
rect 357574 118557 357634 120803
rect 357571 118556 357637 118557
rect 357571 118492 357572 118556
rect 357636 118492 357637 118556
rect 357571 118491 357637 118492
rect 357387 117468 357453 117469
rect 357387 117404 357388 117468
rect 357452 117404 357453 117468
rect 357387 117403 357453 117404
rect 357942 113117 358002 174523
rect 360334 169149 360394 386411
rect 361622 349077 361682 386819
rect 361619 349076 361685 349077
rect 361619 349012 361620 349076
rect 361684 349012 361685 349076
rect 361619 349011 361685 349012
rect 362910 348941 362970 386819
rect 384114 385774 384734 388711
rect 384114 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 384734 385774
rect 384114 385454 384734 385538
rect 384114 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 384734 385454
rect 384114 349774 384734 385218
rect 384114 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 384734 349774
rect 384114 349454 384734 349538
rect 384114 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 384734 349454
rect 362907 348940 362973 348941
rect 362907 348876 362908 348940
rect 362972 348876 362973 348940
rect 362907 348875 362973 348876
rect 384114 348433 384734 349218
rect 420114 385774 420734 388711
rect 420114 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 420734 385774
rect 420114 385454 420734 385538
rect 420114 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 420734 385454
rect 420114 349774 420734 385218
rect 420114 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 420734 349774
rect 456114 385774 456734 388711
rect 456114 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 456734 385774
rect 456114 385454 456734 385538
rect 456114 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 456734 385454
rect 456114 349740 456734 385218
rect 492114 385774 492734 388711
rect 492114 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 492734 385774
rect 492114 385454 492734 385538
rect 492114 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 492734 385454
rect 492114 349774 492734 385218
rect 420114 349454 420734 349538
rect 420114 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 420734 349454
rect 420114 348433 420734 349218
rect 492114 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 492734 349774
rect 492114 349454 492734 349538
rect 492114 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 492734 349454
rect 492114 348433 492734 349218
rect 379568 331174 379888 331206
rect 379568 330938 379610 331174
rect 379846 330938 379888 331174
rect 379568 330854 379888 330938
rect 379568 330618 379610 330854
rect 379846 330618 379888 330854
rect 379568 330586 379888 330618
rect 410288 331174 410608 331206
rect 410288 330938 410330 331174
rect 410566 330938 410608 331174
rect 410288 330854 410608 330938
rect 410288 330618 410330 330854
rect 410566 330618 410608 330854
rect 410288 330586 410608 330618
rect 441008 331174 441328 331206
rect 441008 330938 441050 331174
rect 441286 330938 441328 331174
rect 441008 330854 441328 330938
rect 441008 330618 441050 330854
rect 441286 330618 441328 330854
rect 441008 330586 441328 330618
rect 471728 331174 472048 331206
rect 471728 330938 471770 331174
rect 472006 330938 472048 331174
rect 471728 330854 472048 330938
rect 471728 330618 471770 330854
rect 472006 330618 472048 330854
rect 471728 330586 472048 330618
rect 364208 327454 364528 327486
rect 364208 327218 364250 327454
rect 364486 327218 364528 327454
rect 364208 327134 364528 327218
rect 364208 326898 364250 327134
rect 364486 326898 364528 327134
rect 364208 326866 364528 326898
rect 394928 327454 395248 327486
rect 394928 327218 394970 327454
rect 395206 327218 395248 327454
rect 394928 327134 395248 327218
rect 394928 326898 394970 327134
rect 395206 326898 395248 327134
rect 394928 326866 395248 326898
rect 425648 327454 425968 327486
rect 425648 327218 425690 327454
rect 425926 327218 425968 327454
rect 425648 327134 425968 327218
rect 425648 326898 425690 327134
rect 425926 326898 425968 327134
rect 425648 326866 425968 326898
rect 456368 327454 456688 327486
rect 456368 327218 456410 327454
rect 456646 327218 456688 327454
rect 456368 327134 456688 327218
rect 456368 326898 456410 327134
rect 456646 326898 456688 327134
rect 456368 326866 456688 326898
rect 487088 327454 487408 327486
rect 487088 327218 487130 327454
rect 487366 327218 487408 327454
rect 487088 327134 487408 327218
rect 487088 326898 487130 327134
rect 487366 326898 487408 327134
rect 487088 326866 487408 326898
rect 379568 295174 379888 295206
rect 379568 294938 379610 295174
rect 379846 294938 379888 295174
rect 379568 294854 379888 294938
rect 379568 294618 379610 294854
rect 379846 294618 379888 294854
rect 379568 294586 379888 294618
rect 410288 295174 410608 295206
rect 410288 294938 410330 295174
rect 410566 294938 410608 295174
rect 410288 294854 410608 294938
rect 410288 294618 410330 294854
rect 410566 294618 410608 294854
rect 410288 294586 410608 294618
rect 441008 295174 441328 295206
rect 441008 294938 441050 295174
rect 441286 294938 441328 295174
rect 441008 294854 441328 294938
rect 441008 294618 441050 294854
rect 441286 294618 441328 294854
rect 441008 294586 441328 294618
rect 471728 295174 472048 295206
rect 471728 294938 471770 295174
rect 472006 294938 472048 295174
rect 471728 294854 472048 294938
rect 471728 294618 471770 294854
rect 472006 294618 472048 294854
rect 471728 294586 472048 294618
rect 364208 291454 364528 291486
rect 364208 291218 364250 291454
rect 364486 291218 364528 291454
rect 364208 291134 364528 291218
rect 364208 290898 364250 291134
rect 364486 290898 364528 291134
rect 364208 290866 364528 290898
rect 394928 291454 395248 291486
rect 394928 291218 394970 291454
rect 395206 291218 395248 291454
rect 394928 291134 395248 291218
rect 394928 290898 394970 291134
rect 395206 290898 395248 291134
rect 394928 290866 395248 290898
rect 425648 291454 425968 291486
rect 425648 291218 425690 291454
rect 425926 291218 425968 291454
rect 425648 291134 425968 291218
rect 425648 290898 425690 291134
rect 425926 290898 425968 291134
rect 425648 290866 425968 290898
rect 456368 291454 456688 291486
rect 456368 291218 456410 291454
rect 456646 291218 456688 291454
rect 456368 291134 456688 291218
rect 456368 290898 456410 291134
rect 456646 290898 456688 291134
rect 456368 290866 456688 290898
rect 487088 291454 487408 291486
rect 487088 291218 487130 291454
rect 487366 291218 487408 291454
rect 487088 291134 487408 291218
rect 487088 290898 487130 291134
rect 487366 290898 487408 291134
rect 487088 290866 487408 290898
rect 379568 259174 379888 259206
rect 379568 258938 379610 259174
rect 379846 258938 379888 259174
rect 379568 258854 379888 258938
rect 379568 258618 379610 258854
rect 379846 258618 379888 258854
rect 379568 258586 379888 258618
rect 410288 259174 410608 259206
rect 410288 258938 410330 259174
rect 410566 258938 410608 259174
rect 410288 258854 410608 258938
rect 410288 258618 410330 258854
rect 410566 258618 410608 258854
rect 410288 258586 410608 258618
rect 441008 259174 441328 259206
rect 441008 258938 441050 259174
rect 441286 258938 441328 259174
rect 441008 258854 441328 258938
rect 441008 258618 441050 258854
rect 441286 258618 441328 258854
rect 441008 258586 441328 258618
rect 471728 259174 472048 259206
rect 471728 258938 471770 259174
rect 472006 258938 472048 259174
rect 471728 258854 472048 258938
rect 471728 258618 471770 258854
rect 472006 258618 472048 258854
rect 471728 258586 472048 258618
rect 364208 255454 364528 255486
rect 364208 255218 364250 255454
rect 364486 255218 364528 255454
rect 364208 255134 364528 255218
rect 364208 254898 364250 255134
rect 364486 254898 364528 255134
rect 364208 254866 364528 254898
rect 394928 255454 395248 255486
rect 394928 255218 394970 255454
rect 395206 255218 395248 255454
rect 394928 255134 395248 255218
rect 394928 254898 394970 255134
rect 395206 254898 395248 255134
rect 394928 254866 395248 254898
rect 425648 255454 425968 255486
rect 425648 255218 425690 255454
rect 425926 255218 425968 255454
rect 425648 255134 425968 255218
rect 425648 254898 425690 255134
rect 425926 254898 425968 255134
rect 425648 254866 425968 254898
rect 456368 255454 456688 255486
rect 456368 255218 456410 255454
rect 456646 255218 456688 255454
rect 456368 255134 456688 255218
rect 456368 254898 456410 255134
rect 456646 254898 456688 255134
rect 456368 254866 456688 254898
rect 487088 255454 487408 255486
rect 487088 255218 487130 255454
rect 487366 255218 487408 255454
rect 487088 255134 487408 255218
rect 487088 254898 487130 255134
rect 487366 254898 487408 255134
rect 487088 254866 487408 254898
rect 379568 223174 379888 223206
rect 379568 222938 379610 223174
rect 379846 222938 379888 223174
rect 379568 222854 379888 222938
rect 379568 222618 379610 222854
rect 379846 222618 379888 222854
rect 379568 222586 379888 222618
rect 410288 223174 410608 223206
rect 410288 222938 410330 223174
rect 410566 222938 410608 223174
rect 410288 222854 410608 222938
rect 410288 222618 410330 222854
rect 410566 222618 410608 222854
rect 410288 222586 410608 222618
rect 441008 223174 441328 223206
rect 441008 222938 441050 223174
rect 441286 222938 441328 223174
rect 441008 222854 441328 222938
rect 441008 222618 441050 222854
rect 441286 222618 441328 222854
rect 441008 222586 441328 222618
rect 471728 223174 472048 223206
rect 471728 222938 471770 223174
rect 472006 222938 472048 223174
rect 471728 222854 472048 222938
rect 471728 222618 471770 222854
rect 472006 222618 472048 222854
rect 471728 222586 472048 222618
rect 364208 219454 364528 219486
rect 364208 219218 364250 219454
rect 364486 219218 364528 219454
rect 364208 219134 364528 219218
rect 364208 218898 364250 219134
rect 364486 218898 364528 219134
rect 364208 218866 364528 218898
rect 394928 219454 395248 219486
rect 394928 219218 394970 219454
rect 395206 219218 395248 219454
rect 394928 219134 395248 219218
rect 394928 218898 394970 219134
rect 395206 218898 395248 219134
rect 394928 218866 395248 218898
rect 425648 219454 425968 219486
rect 425648 219218 425690 219454
rect 425926 219218 425968 219454
rect 425648 219134 425968 219218
rect 425648 218898 425690 219134
rect 425926 218898 425968 219134
rect 425648 218866 425968 218898
rect 456368 219454 456688 219486
rect 456368 219218 456410 219454
rect 456646 219218 456688 219454
rect 456368 219134 456688 219218
rect 456368 218898 456410 219134
rect 456646 218898 456688 219134
rect 456368 218866 456688 218898
rect 487088 219454 487408 219486
rect 487088 219218 487130 219454
rect 487366 219218 487408 219454
rect 487088 219134 487408 219218
rect 487088 218898 487130 219134
rect 487366 218898 487408 219134
rect 487088 218866 487408 218898
rect 379568 187174 379888 187206
rect 379568 186938 379610 187174
rect 379846 186938 379888 187174
rect 379568 186854 379888 186938
rect 379568 186618 379610 186854
rect 379846 186618 379888 186854
rect 379568 186586 379888 186618
rect 410288 187174 410608 187206
rect 410288 186938 410330 187174
rect 410566 186938 410608 187174
rect 410288 186854 410608 186938
rect 410288 186618 410330 186854
rect 410566 186618 410608 186854
rect 410288 186586 410608 186618
rect 441008 187174 441328 187206
rect 441008 186938 441050 187174
rect 441286 186938 441328 187174
rect 441008 186854 441328 186938
rect 441008 186618 441050 186854
rect 441286 186618 441328 186854
rect 441008 186586 441328 186618
rect 471728 187174 472048 187206
rect 471728 186938 471770 187174
rect 472006 186938 472048 187174
rect 471728 186854 472048 186938
rect 471728 186618 471770 186854
rect 472006 186618 472048 186854
rect 471728 186586 472048 186618
rect 364208 183454 364528 183486
rect 364208 183218 364250 183454
rect 364486 183218 364528 183454
rect 364208 183134 364528 183218
rect 364208 182898 364250 183134
rect 364486 182898 364528 183134
rect 364208 182866 364528 182898
rect 394928 183454 395248 183486
rect 394928 183218 394970 183454
rect 395206 183218 395248 183454
rect 394928 183134 395248 183218
rect 394928 182898 394970 183134
rect 395206 182898 395248 183134
rect 394928 182866 395248 182898
rect 425648 183454 425968 183486
rect 425648 183218 425690 183454
rect 425926 183218 425968 183454
rect 425648 183134 425968 183218
rect 425648 182898 425690 183134
rect 425926 182898 425968 183134
rect 425648 182866 425968 182898
rect 456368 183454 456688 183486
rect 456368 183218 456410 183454
rect 456646 183218 456688 183454
rect 456368 183134 456688 183218
rect 456368 182898 456410 183134
rect 456646 182898 456688 183134
rect 456368 182866 456688 182898
rect 487088 183454 487408 183486
rect 487088 183218 487130 183454
rect 487366 183218 487408 183454
rect 487088 183134 487408 183218
rect 487088 182898 487130 183134
rect 487366 182898 487408 183134
rect 487088 182866 487408 182898
rect 407619 181388 407685 181389
rect 407619 181324 407620 181388
rect 407684 181324 407685 181388
rect 407619 181323 407685 181324
rect 360331 169148 360397 169149
rect 360331 169084 360332 169148
rect 360396 169084 360397 169148
rect 360331 169083 360397 169084
rect 397794 147454 398414 179799
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 379568 115174 379888 115206
rect 379568 114938 379610 115174
rect 379846 114938 379888 115174
rect 379568 114854 379888 114938
rect 379568 114618 379610 114854
rect 379846 114618 379888 114854
rect 379568 114586 379888 114618
rect 357939 113116 358005 113117
rect 357939 113052 357940 113116
rect 358004 113052 358005 113116
rect 357939 113051 358005 113052
rect 356651 112708 356717 112709
rect 356651 112644 356652 112708
rect 356716 112644 356717 112708
rect 356651 112643 356717 112644
rect 364208 111454 364528 111486
rect 364208 111218 364250 111454
rect 364486 111218 364528 111454
rect 364208 111134 364528 111218
rect 364208 110898 364250 111134
rect 364486 110898 364528 111134
rect 364208 110866 364528 110898
rect 394928 111454 395248 111486
rect 394928 111218 394970 111454
rect 395206 111218 395248 111454
rect 394928 111134 395248 111218
rect 394928 110898 394970 111134
rect 395206 110898 395248 111134
rect 394928 110866 395248 110898
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 351834 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 352454 101494
rect 351834 101174 352454 101258
rect 351834 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 352454 101174
rect 351834 65494 352454 100938
rect 351834 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 352454 65494
rect 351834 65174 352454 65258
rect 351834 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 352454 65174
rect 351834 29494 352454 64938
rect 351834 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 352454 29494
rect 351834 29174 352454 29258
rect 351834 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 352454 29174
rect 351834 -7066 352454 28938
rect 351834 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 352454 -7066
rect 351834 -7386 352454 -7302
rect 351834 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 352454 -7386
rect 351834 -7654 352454 -7622
rect 361794 75454 362414 100479
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -7654 362414 -902
rect 365514 79174 366134 100479
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -1306 366134 6618
rect 365514 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 366134 -1306
rect 365514 -1626 366134 -1542
rect 365514 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 366134 -1626
rect 365514 -7654 366134 -1862
rect 369234 82894 369854 100479
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -2266 369854 10338
rect 369234 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 369854 -2266
rect 369234 -2586 369854 -2502
rect 369234 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 369854 -2586
rect 369234 -7654 369854 -2822
rect 372954 86614 373574 100479
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 372954 -3226 373574 14058
rect 372954 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 373574 -3226
rect 372954 -3546 373574 -3462
rect 372954 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 373574 -3546
rect 372954 -7654 373574 -3782
rect 376674 90334 377294 100479
rect 376674 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 377294 90334
rect 376674 90014 377294 90098
rect 376674 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 377294 90014
rect 376674 54334 377294 89778
rect 376674 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 377294 54334
rect 376674 54014 377294 54098
rect 376674 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 377294 54014
rect 376674 18334 377294 53778
rect 376674 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 377294 18334
rect 376674 18014 377294 18098
rect 376674 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 377294 18014
rect 376674 -4186 377294 17778
rect 376674 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 377294 -4186
rect 376674 -4506 377294 -4422
rect 376674 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 377294 -4506
rect 376674 -7654 377294 -4742
rect 380394 94054 381014 100479
rect 380394 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 381014 94054
rect 380394 93734 381014 93818
rect 380394 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 381014 93734
rect 380394 58054 381014 93498
rect 380394 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 381014 58054
rect 380394 57734 381014 57818
rect 380394 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 381014 57734
rect 380394 22054 381014 57498
rect 380394 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 381014 22054
rect 380394 21734 381014 21818
rect 380394 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 381014 21734
rect 380394 -5146 381014 21498
rect 380394 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 381014 -5146
rect 380394 -5466 381014 -5382
rect 380394 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 381014 -5466
rect 380394 -7654 381014 -5702
rect 384114 97774 384734 100479
rect 384114 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 384734 97774
rect 384114 97454 384734 97538
rect 384114 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 384734 97454
rect 384114 61774 384734 97218
rect 384114 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 384734 61774
rect 384114 61454 384734 61538
rect 384114 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 384734 61454
rect 384114 25774 384734 61218
rect 384114 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 384734 25774
rect 384114 25454 384734 25538
rect 384114 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 384734 25454
rect 384114 -6106 384734 25218
rect 384114 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 384734 -6106
rect 384114 -6426 384734 -6342
rect 384114 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 384734 -6426
rect 384114 -7654 384734 -6662
rect 387834 65494 388454 100479
rect 387834 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 388454 65494
rect 387834 65174 388454 65258
rect 387834 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 388454 65174
rect 387834 29494 388454 64938
rect 387834 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 388454 29494
rect 387834 29174 388454 29258
rect 387834 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 388454 29174
rect 387834 -7066 388454 28938
rect 387834 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 388454 -7066
rect 387834 -7386 388454 -7302
rect 387834 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 388454 -7386
rect 387834 -7654 388454 -7622
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -7654 398414 -902
rect 401514 151174 402134 179799
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -1306 402134 6618
rect 401514 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 402134 -1306
rect 401514 -1626 402134 -1542
rect 401514 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 402134 -1626
rect 401514 -7654 402134 -1862
rect 405234 154894 405854 179799
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 407622 144805 407682 181323
rect 408954 158614 409574 179799
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 407619 144804 407685 144805
rect 407619 144740 407620 144804
rect 407684 144740 407685 144804
rect 407619 144739 407685 144740
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -2266 405854 10338
rect 405234 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 405854 -2266
rect 405234 -2586 405854 -2502
rect 405234 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 405854 -2586
rect 405234 -7654 405854 -2822
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 408954 -3226 409574 14058
rect 408954 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 409574 -3226
rect 408954 -3546 409574 -3462
rect 408954 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 409574 -3546
rect 408954 -7654 409574 -3782
rect 412674 162334 413294 179799
rect 412674 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 413294 162334
rect 412674 162014 413294 162098
rect 412674 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 413294 162014
rect 412674 126334 413294 161778
rect 412674 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 413294 126334
rect 412674 126014 413294 126098
rect 412674 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 413294 126014
rect 412674 90334 413294 125778
rect 412674 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 413294 90334
rect 412674 90014 413294 90098
rect 412674 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 413294 90014
rect 412674 54334 413294 89778
rect 412674 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 413294 54334
rect 412674 54014 413294 54098
rect 412674 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 413294 54014
rect 412674 18334 413294 53778
rect 412674 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 413294 18334
rect 412674 18014 413294 18098
rect 412674 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 413294 18014
rect 412674 -4186 413294 17778
rect 412674 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 413294 -4186
rect 412674 -4506 413294 -4422
rect 412674 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 413294 -4506
rect 412674 -7654 413294 -4742
rect 416394 166054 417014 179799
rect 416394 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 417014 166054
rect 416394 165734 417014 165818
rect 416394 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 417014 165734
rect 416394 130054 417014 165498
rect 416394 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 417014 130054
rect 416394 129734 417014 129818
rect 416394 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 417014 129734
rect 416394 94054 417014 129498
rect 416394 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 417014 94054
rect 416394 93734 417014 93818
rect 416394 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 417014 93734
rect 416394 58054 417014 93498
rect 416394 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 417014 58054
rect 416394 57734 417014 57818
rect 416394 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 417014 57734
rect 416394 22054 417014 57498
rect 416394 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 417014 22054
rect 416394 21734 417014 21818
rect 416394 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 417014 21734
rect 416394 -5146 417014 21498
rect 416394 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 417014 -5146
rect 416394 -5466 417014 -5382
rect 416394 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 417014 -5466
rect 416394 -7654 417014 -5702
rect 420114 169774 420734 179799
rect 420114 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 420734 169774
rect 420114 169454 420734 169538
rect 420114 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 420734 169454
rect 420114 133774 420734 169218
rect 420114 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 420734 133774
rect 420114 133454 420734 133538
rect 420114 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 420734 133454
rect 420114 97774 420734 133218
rect 420114 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 420734 97774
rect 420114 97454 420734 97538
rect 420114 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 420734 97454
rect 420114 61774 420734 97218
rect 420114 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 420734 61774
rect 420114 61454 420734 61538
rect 420114 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 420734 61454
rect 420114 25774 420734 61218
rect 420114 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 420734 25774
rect 420114 25454 420734 25538
rect 420114 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 420734 25454
rect 420114 -6106 420734 25218
rect 420114 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 420734 -6106
rect 420114 -6426 420734 -6342
rect 420114 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 420734 -6426
rect 420114 -7654 420734 -6662
rect 423834 173494 424454 179799
rect 423834 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 424454 173494
rect 423834 173174 424454 173258
rect 423834 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 424454 173174
rect 423834 137494 424454 172938
rect 423834 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 424454 137494
rect 423834 137174 424454 137258
rect 423834 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 424454 137174
rect 423834 101494 424454 136938
rect 423834 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 424454 101494
rect 423834 101174 424454 101258
rect 423834 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 424454 101174
rect 423834 65494 424454 100938
rect 423834 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 424454 65494
rect 423834 65174 424454 65258
rect 423834 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 424454 65174
rect 423834 29494 424454 64938
rect 423834 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 424454 29494
rect 423834 29174 424454 29258
rect 423834 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 424454 29174
rect 423834 -7066 424454 28938
rect 423834 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 424454 -7066
rect 423834 -7386 424454 -7302
rect 423834 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 424454 -7386
rect 423834 -7654 424454 -7622
rect 433794 147454 434414 179799
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -7654 434414 -902
rect 437514 151174 438134 179799
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -1306 438134 6618
rect 437514 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 438134 -1306
rect 437514 -1626 438134 -1542
rect 437514 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 438134 -1626
rect 437514 -7654 438134 -1862
rect 441234 154894 441854 179799
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -2266 441854 10338
rect 441234 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 441854 -2266
rect 441234 -2586 441854 -2502
rect 441234 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 441854 -2586
rect 441234 -7654 441854 -2822
rect 444954 158614 445574 179799
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 444954 -3226 445574 14058
rect 444954 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 445574 -3226
rect 444954 -3546 445574 -3462
rect 444954 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 445574 -3546
rect 444954 -7654 445574 -3782
rect 448674 162334 449294 179799
rect 448674 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 449294 162334
rect 448674 162014 449294 162098
rect 448674 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 449294 162014
rect 448674 126334 449294 161778
rect 448674 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 449294 126334
rect 448674 126014 449294 126098
rect 448674 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 449294 126014
rect 448674 90334 449294 125778
rect 448674 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 449294 90334
rect 448674 90014 449294 90098
rect 448674 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 449294 90014
rect 448674 54334 449294 89778
rect 448674 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 449294 54334
rect 448674 54014 449294 54098
rect 448674 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 449294 54014
rect 448674 18334 449294 53778
rect 448674 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 449294 18334
rect 448674 18014 449294 18098
rect 448674 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 449294 18014
rect 448674 -4186 449294 17778
rect 448674 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 449294 -4186
rect 448674 -4506 449294 -4422
rect 448674 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 449294 -4506
rect 448674 -7654 449294 -4742
rect 452394 166054 453014 179799
rect 452394 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 453014 166054
rect 452394 165734 453014 165818
rect 452394 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 453014 165734
rect 452394 130054 453014 165498
rect 452394 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 453014 130054
rect 452394 129734 453014 129818
rect 452394 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 453014 129734
rect 452394 94054 453014 129498
rect 452394 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 453014 94054
rect 452394 93734 453014 93818
rect 452394 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 453014 93734
rect 452394 58054 453014 93498
rect 452394 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 453014 58054
rect 452394 57734 453014 57818
rect 452394 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 453014 57734
rect 452394 22054 453014 57498
rect 452394 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 453014 22054
rect 452394 21734 453014 21818
rect 452394 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 453014 21734
rect 452394 -5146 453014 21498
rect 452394 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 453014 -5146
rect 452394 -5466 453014 -5382
rect 452394 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 453014 -5466
rect 452394 -7654 453014 -5702
rect 456114 169774 456734 179799
rect 456114 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 456734 169774
rect 456114 169454 456734 169538
rect 456114 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 456734 169454
rect 456114 133774 456734 169218
rect 456114 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 456734 133774
rect 456114 133454 456734 133538
rect 456114 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 456734 133454
rect 456114 97774 456734 133218
rect 456114 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 456734 97774
rect 456114 97454 456734 97538
rect 456114 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 456734 97454
rect 456114 61774 456734 97218
rect 456114 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 456734 61774
rect 456114 61454 456734 61538
rect 456114 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 456734 61454
rect 456114 25774 456734 61218
rect 456114 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 456734 25774
rect 456114 25454 456734 25538
rect 456114 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 456734 25454
rect 456114 -6106 456734 25218
rect 456114 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 456734 -6106
rect 456114 -6426 456734 -6342
rect 456114 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 456734 -6426
rect 456114 -7654 456734 -6662
rect 459834 173494 460454 179799
rect 459834 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 460454 173494
rect 459834 173174 460454 173258
rect 459834 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 460454 173174
rect 459834 137494 460454 172938
rect 459834 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 460454 137494
rect 459834 137174 460454 137258
rect 459834 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 460454 137174
rect 459834 101494 460454 136938
rect 459834 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 460454 101494
rect 459834 101174 460454 101258
rect 459834 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 460454 101174
rect 459834 65494 460454 100938
rect 459834 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 460454 65494
rect 459834 65174 460454 65258
rect 459834 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 460454 65174
rect 459834 29494 460454 64938
rect 459834 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 460454 29494
rect 459834 29174 460454 29258
rect 459834 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 460454 29174
rect 459834 -7066 460454 28938
rect 459834 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 460454 -7066
rect 459834 -7386 460454 -7302
rect 459834 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 460454 -7386
rect 459834 -7654 460454 -7622
rect 469794 147454 470414 179799
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -7654 470414 -902
rect 473514 151174 474134 179799
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -1306 474134 6618
rect 473514 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 474134 -1306
rect 473514 -1626 474134 -1542
rect 473514 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 474134 -1626
rect 473514 -7654 474134 -1862
rect 477234 154894 477854 179799
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -2266 477854 10338
rect 477234 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 477854 -2266
rect 477234 -2586 477854 -2502
rect 477234 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 477854 -2586
rect 477234 -7654 477854 -2822
rect 480954 158614 481574 179799
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 480954 -3226 481574 14058
rect 480954 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 481574 -3226
rect 480954 -3546 481574 -3462
rect 480954 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 481574 -3546
rect 480954 -7654 481574 -3782
rect 484674 162334 485294 179799
rect 484674 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 485294 162334
rect 484674 162014 485294 162098
rect 484674 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 485294 162014
rect 484674 126334 485294 161778
rect 484674 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 485294 126334
rect 484674 126014 485294 126098
rect 484674 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 485294 126014
rect 484674 90334 485294 125778
rect 484674 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 485294 90334
rect 484674 90014 485294 90098
rect 484674 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 485294 90014
rect 484674 54334 485294 89778
rect 484674 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 485294 54334
rect 484674 54014 485294 54098
rect 484674 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 485294 54014
rect 484674 18334 485294 53778
rect 484674 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 485294 18334
rect 484674 18014 485294 18098
rect 484674 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 485294 18014
rect 484674 -4186 485294 17778
rect 484674 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 485294 -4186
rect 484674 -4506 485294 -4422
rect 484674 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 485294 -4506
rect 484674 -7654 485294 -4742
rect 488394 166054 489014 179799
rect 488394 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 489014 166054
rect 488394 165734 489014 165818
rect 488394 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 489014 165734
rect 488394 130054 489014 165498
rect 488394 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 489014 130054
rect 488394 129734 489014 129818
rect 488394 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 489014 129734
rect 488394 94054 489014 129498
rect 488394 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 489014 94054
rect 488394 93734 489014 93818
rect 488394 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 489014 93734
rect 488394 58054 489014 93498
rect 488394 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 489014 58054
rect 488394 57734 489014 57818
rect 488394 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 489014 57734
rect 488394 22054 489014 57498
rect 488394 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 489014 22054
rect 488394 21734 489014 21818
rect 488394 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 489014 21734
rect 488394 -5146 489014 21498
rect 488394 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 489014 -5146
rect 488394 -5466 489014 -5382
rect 488394 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 489014 -5466
rect 488394 -7654 489014 -5702
rect 492114 169774 492734 179799
rect 492114 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 492734 169774
rect 492114 169454 492734 169538
rect 492114 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 492734 169454
rect 492114 133774 492734 169218
rect 492114 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 492734 133774
rect 492114 133454 492734 133538
rect 492114 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 492734 133454
rect 492114 97774 492734 133218
rect 492114 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 492734 97774
rect 492114 97454 492734 97538
rect 492114 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 492734 97454
rect 492114 61774 492734 97218
rect 492114 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 492734 61774
rect 492114 61454 492734 61538
rect 492114 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 492734 61454
rect 492114 25774 492734 61218
rect 492114 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 492734 25774
rect 492114 25454 492734 25538
rect 492114 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 492734 25454
rect 492114 -6106 492734 25218
rect 492114 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 492734 -6106
rect 492114 -6426 492734 -6342
rect 492114 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 492734 -6426
rect 492114 -7654 492734 -6662
rect 495834 173494 496454 179799
rect 499622 176085 499682 534107
rect 499803 531452 499869 531453
rect 499803 531388 499804 531452
rect 499868 531388 499869 531452
rect 499803 531387 499869 531388
rect 499806 177309 499866 531387
rect 499987 520300 500053 520301
rect 499987 520236 499988 520300
rect 500052 520236 500053 520300
rect 499987 520235 500053 520236
rect 499990 478410 500050 520235
rect 500174 482901 500234 599659
rect 504219 598092 504285 598093
rect 504219 598028 504220 598092
rect 504284 598028 504285 598092
rect 504219 598027 504285 598028
rect 502379 550628 502445 550629
rect 502379 550564 502380 550628
rect 502444 550564 502445 550628
rect 502379 550563 502445 550564
rect 501275 529276 501341 529277
rect 501275 529212 501276 529276
rect 501340 529212 501341 529276
rect 501275 529211 501341 529212
rect 500723 521932 500789 521933
rect 500723 521868 500724 521932
rect 500788 521868 500789 521932
rect 500723 521867 500789 521868
rect 500539 521660 500605 521661
rect 500539 521596 500540 521660
rect 500604 521596 500605 521660
rect 500539 521595 500605 521596
rect 500355 520708 500421 520709
rect 500355 520644 500356 520708
rect 500420 520644 500421 520708
rect 500355 520643 500421 520644
rect 500358 519485 500418 520643
rect 500542 519757 500602 521595
rect 500539 519756 500605 519757
rect 500539 519692 500540 519756
rect 500604 519692 500605 519756
rect 500539 519691 500605 519692
rect 500726 519621 500786 521867
rect 501091 520028 501157 520029
rect 501091 519964 501092 520028
rect 501156 519964 501157 520028
rect 501091 519963 501157 519964
rect 500723 519620 500789 519621
rect 500723 519556 500724 519620
rect 500788 519556 500789 519620
rect 500723 519555 500789 519556
rect 500355 519484 500421 519485
rect 500355 519420 500356 519484
rect 500420 519420 500421 519484
rect 500355 519419 500421 519420
rect 500171 482900 500237 482901
rect 500171 482836 500172 482900
rect 500236 482836 500237 482900
rect 500171 482835 500237 482836
rect 500539 482220 500605 482221
rect 500539 482156 500540 482220
rect 500604 482156 500605 482220
rect 500539 482155 500605 482156
rect 499990 478350 500418 478410
rect 500358 475285 500418 478350
rect 500355 475284 500421 475285
rect 500355 475220 500356 475284
rect 500420 475220 500421 475284
rect 500355 475219 500421 475220
rect 500542 475010 500602 482155
rect 500174 474950 500602 475010
rect 499803 177308 499869 177309
rect 499803 177244 499804 177308
rect 499868 177244 499869 177308
rect 499803 177243 499869 177244
rect 499619 176084 499685 176085
rect 499619 176020 499620 176084
rect 499684 176020 499685 176084
rect 499619 176019 499685 176020
rect 500174 175133 500234 474950
rect 500355 474604 500421 474605
rect 500355 474540 500356 474604
rect 500420 474540 500421 474604
rect 500355 474539 500421 474540
rect 500358 388109 500418 474539
rect 501094 390013 501154 519963
rect 501278 454613 501338 529211
rect 501643 528596 501709 528597
rect 501643 528532 501644 528596
rect 501708 528532 501709 528596
rect 501643 528531 501709 528532
rect 501459 526556 501525 526557
rect 501459 526492 501460 526556
rect 501524 526492 501525 526556
rect 501459 526491 501525 526492
rect 501462 481405 501522 526491
rect 501459 481404 501525 481405
rect 501459 481340 501460 481404
rect 501524 481340 501525 481404
rect 501459 481339 501525 481340
rect 501275 454612 501341 454613
rect 501275 454548 501276 454612
rect 501340 454548 501341 454612
rect 501275 454547 501341 454548
rect 501091 390012 501157 390013
rect 501091 389948 501092 390012
rect 501156 389948 501157 390012
rect 501091 389947 501157 389948
rect 500355 388108 500421 388109
rect 500355 388044 500356 388108
rect 500420 388044 500421 388108
rect 500355 388043 500421 388044
rect 500171 175132 500237 175133
rect 500171 175068 500172 175132
rect 500236 175068 500237 175132
rect 500171 175067 500237 175068
rect 501646 174997 501706 528531
rect 502382 480181 502442 550563
rect 503667 546548 503733 546549
rect 503667 546484 503668 546548
rect 503732 546484 503733 546548
rect 503667 546483 503733 546484
rect 502563 545052 502629 545053
rect 502563 544988 502564 545052
rect 502628 544988 502629 545052
rect 502563 544987 502629 544988
rect 502566 480453 502626 544987
rect 502931 540972 502997 540973
rect 502931 540908 502932 540972
rect 502996 540908 502997 540972
rect 502931 540907 502997 540908
rect 502747 526828 502813 526829
rect 502747 526764 502748 526828
rect 502812 526764 502813 526828
rect 502747 526763 502813 526764
rect 502563 480452 502629 480453
rect 502563 480388 502564 480452
rect 502628 480388 502629 480452
rect 502563 480387 502629 480388
rect 502379 480180 502445 480181
rect 502379 480116 502380 480180
rect 502444 480116 502445 480180
rect 502379 480115 502445 480116
rect 502750 479365 502810 526763
rect 502934 520301 502994 540907
rect 503115 521388 503181 521389
rect 503115 521324 503116 521388
rect 503180 521324 503181 521388
rect 503115 521323 503181 521324
rect 502931 520300 502997 520301
rect 502931 520236 502932 520300
rect 502996 520236 502997 520300
rect 502931 520235 502997 520236
rect 503118 509250 503178 521323
rect 502934 509190 503178 509250
rect 502747 479364 502813 479365
rect 502747 479300 502748 479364
rect 502812 479300 502813 479364
rect 502747 479299 502813 479300
rect 502934 479093 502994 509190
rect 503115 481404 503181 481405
rect 503115 481340 503116 481404
rect 503180 481340 503181 481404
rect 503115 481339 503181 481340
rect 502931 479092 502997 479093
rect 502931 479028 502932 479092
rect 502996 479028 502997 479092
rect 502931 479027 502997 479028
rect 503118 178805 503178 481339
rect 503670 178941 503730 546483
rect 503851 523156 503917 523157
rect 503851 523092 503852 523156
rect 503916 523092 503917 523156
rect 503851 523091 503917 523092
rect 503667 178940 503733 178941
rect 503667 178876 503668 178940
rect 503732 178876 503733 178940
rect 503667 178875 503733 178876
rect 503115 178804 503181 178805
rect 503115 178740 503116 178804
rect 503180 178740 503181 178804
rect 503115 178739 503181 178740
rect 501643 174996 501709 174997
rect 501643 174932 501644 174996
rect 501708 174932 501709 174996
rect 501643 174931 501709 174932
rect 503854 174861 503914 523091
rect 504035 519620 504101 519621
rect 504035 519556 504036 519620
rect 504100 519556 504101 519620
rect 504035 519555 504101 519556
rect 504038 512005 504098 519555
rect 504035 512004 504101 512005
rect 504035 511940 504036 512004
rect 504100 511940 504101 512004
rect 504035 511939 504101 511940
rect 504035 511868 504101 511869
rect 504035 511804 504036 511868
rect 504100 511804 504101 511868
rect 504035 511803 504101 511804
rect 504038 179349 504098 511803
rect 504222 354381 504282 598027
rect 505794 579454 506414 600207
rect 506979 598092 507045 598093
rect 506979 598028 506980 598092
rect 507044 598028 507045 598092
rect 506979 598027 507045 598028
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505139 557292 505205 557293
rect 505139 557228 505140 557292
rect 505204 557228 505205 557292
rect 505139 557227 505205 557228
rect 505142 478821 505202 557227
rect 505794 543454 506414 578898
rect 506611 547908 506677 547909
rect 506611 547844 506612 547908
rect 506676 547844 506677 547908
rect 506611 547843 506677 547844
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505323 521252 505389 521253
rect 505323 521188 505324 521252
rect 505388 521188 505389 521252
rect 505323 521187 505389 521188
rect 505139 478820 505205 478821
rect 505139 478756 505140 478820
rect 505204 478756 505205 478820
rect 505139 478755 505205 478756
rect 505326 475829 505386 521187
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505323 475828 505389 475829
rect 505323 475764 505324 475828
rect 505388 475764 505389 475828
rect 505323 475763 505389 475764
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 504219 354380 504285 354381
rect 504219 354316 504220 354380
rect 504284 354316 504285 354380
rect 504219 354315 504285 354316
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 504035 179348 504101 179349
rect 504035 179284 504036 179348
rect 504100 179284 504101 179348
rect 504035 179283 504101 179284
rect 503851 174860 503917 174861
rect 503851 174796 503852 174860
rect 503916 174796 503917 174860
rect 503851 174795 503917 174796
rect 495834 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 496454 173494
rect 495834 173174 496454 173258
rect 495834 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 496454 173174
rect 495834 137494 496454 172938
rect 495834 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 496454 137494
rect 495834 137174 496454 137258
rect 495834 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 496454 137174
rect 495834 101494 496454 136938
rect 495834 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 496454 101494
rect 495834 101174 496454 101258
rect 495834 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 496454 101174
rect 495834 65494 496454 100938
rect 495834 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 496454 65494
rect 495834 65174 496454 65258
rect 495834 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 496454 65174
rect 495834 29494 496454 64938
rect 495834 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 496454 29494
rect 495834 29174 496454 29258
rect 495834 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 496454 29174
rect 495834 -7066 496454 28938
rect 495834 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 496454 -7066
rect 495834 -7386 496454 -7302
rect 495834 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 496454 -7386
rect 495834 -7654 496454 -7622
rect 505794 147454 506414 182898
rect 506614 174589 506674 547843
rect 506795 541108 506861 541109
rect 506795 541044 506796 541108
rect 506860 541044 506861 541108
rect 506795 541043 506861 541044
rect 506798 175269 506858 541043
rect 506982 354245 507042 598027
rect 509514 583174 510134 599988
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 507899 554844 507965 554845
rect 507899 554780 507900 554844
rect 507964 554780 507965 554844
rect 507899 554779 507965 554780
rect 507163 519756 507229 519757
rect 507163 519692 507164 519756
rect 507228 519692 507229 519756
rect 507163 519691 507229 519692
rect 507166 483989 507226 519691
rect 507163 483988 507229 483989
rect 507163 483924 507164 483988
rect 507228 483924 507229 483988
rect 507163 483923 507229 483924
rect 506979 354244 507045 354245
rect 506979 354180 506980 354244
rect 507044 354180 507045 354244
rect 506979 354179 507045 354180
rect 506795 175268 506861 175269
rect 506795 175204 506796 175268
rect 506860 175204 506861 175268
rect 506795 175203 506861 175204
rect 507902 174725 507962 554779
rect 509187 550764 509253 550765
rect 509187 550700 509188 550764
rect 509252 550700 509253 550764
rect 509187 550699 509253 550700
rect 509190 550490 509250 550699
rect 509006 550430 509250 550490
rect 508267 546276 508333 546277
rect 508267 546212 508268 546276
rect 508332 546212 508333 546276
rect 508267 546211 508333 546212
rect 508083 521116 508149 521117
rect 508083 521052 508084 521116
rect 508148 521052 508149 521116
rect 508083 521051 508149 521052
rect 507899 174724 507965 174725
rect 507899 174660 507900 174724
rect 507964 174660 507965 174724
rect 507899 174659 507965 174660
rect 506611 174588 506677 174589
rect 506611 174524 506612 174588
rect 506676 174524 506677 174588
rect 506611 174523 506677 174524
rect 508086 159221 508146 521051
rect 508270 484261 508330 546211
rect 508451 520844 508517 520845
rect 508451 520780 508452 520844
rect 508516 520780 508517 520844
rect 508451 520779 508517 520780
rect 508267 484260 508333 484261
rect 508267 484196 508268 484260
rect 508332 484196 508333 484260
rect 508267 484195 508333 484196
rect 508454 475013 508514 520779
rect 509006 514770 509066 550430
rect 509514 547174 510134 582618
rect 513234 586894 513854 600207
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 512131 559060 512197 559061
rect 512131 558996 512132 559060
rect 512196 558996 512197 559060
rect 512131 558995 512197 558996
rect 511027 550084 511093 550085
rect 511027 550020 511028 550084
rect 511092 550020 511093 550084
rect 511027 550019 511093 550020
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509006 514710 509250 514770
rect 509190 505110 509250 514710
rect 509006 505050 509250 505110
rect 509514 511174 510134 546618
rect 510659 540700 510725 540701
rect 510659 540636 510660 540700
rect 510724 540636 510725 540700
rect 510659 540635 510725 540636
rect 510475 532812 510541 532813
rect 510475 532748 510476 532812
rect 510540 532748 510541 532812
rect 510475 532747 510541 532748
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 508451 475012 508517 475013
rect 508451 474948 508452 475012
rect 508516 474948 508517 475012
rect 508451 474947 508517 474948
rect 508451 258908 508517 258909
rect 508451 258844 508452 258908
rect 508516 258844 508517 258908
rect 508451 258843 508517 258844
rect 508083 159220 508149 159221
rect 508083 159156 508084 159220
rect 508148 159156 508149 159220
rect 508083 159155 508149 159156
rect 508454 153781 508514 258843
rect 509006 176357 509066 505050
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509003 176356 509069 176357
rect 509003 176292 509004 176356
rect 509068 176292 509069 176356
rect 509003 176291 509069 176292
rect 508451 153780 508517 153781
rect 508451 153716 508452 153780
rect 508516 153716 508517 153780
rect 508451 153715 508517 153716
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -7654 506414 -902
rect 509514 151174 510134 186618
rect 510478 176629 510538 532747
rect 510662 179077 510722 540635
rect 510843 513500 510909 513501
rect 510843 513436 510844 513500
rect 510908 513436 510909 513500
rect 510843 513435 510909 513436
rect 510659 179076 510725 179077
rect 510659 179012 510660 179076
rect 510724 179012 510725 179076
rect 510659 179011 510725 179012
rect 510475 176628 510541 176629
rect 510475 176564 510476 176628
rect 510540 176564 510541 176628
rect 510475 176563 510541 176564
rect 510846 176221 510906 513435
rect 511030 478005 511090 550019
rect 511947 527236 512013 527237
rect 511947 527172 511948 527236
rect 512012 527172 512013 527236
rect 511947 527171 512013 527172
rect 511211 519348 511277 519349
rect 511211 519284 511212 519348
rect 511276 519284 511277 519348
rect 511211 519283 511277 519284
rect 511214 480317 511274 519283
rect 511211 480316 511277 480317
rect 511211 480252 511212 480316
rect 511276 480252 511277 480316
rect 511211 480251 511277 480252
rect 511950 480270 512010 527171
rect 512134 481405 512194 558995
rect 513234 550894 513854 586338
rect 516954 590614 517574 600207
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 515259 558244 515325 558245
rect 515259 558180 515260 558244
rect 515324 558180 515325 558244
rect 515259 558179 515325 558180
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 512315 526964 512381 526965
rect 512315 526900 512316 526964
rect 512380 526900 512381 526964
rect 512315 526899 512381 526900
rect 512131 481404 512197 481405
rect 512131 481340 512132 481404
rect 512196 481340 512197 481404
rect 512131 481339 512197 481340
rect 511950 480210 512194 480270
rect 511027 478004 511093 478005
rect 511027 477940 511028 478004
rect 511092 477940 511093 478004
rect 511027 477939 511093 477940
rect 512134 177853 512194 480210
rect 512318 472837 512378 526899
rect 512499 524516 512565 524517
rect 512499 524452 512500 524516
rect 512564 524452 512565 524516
rect 512499 524451 512565 524452
rect 512502 482221 512562 524451
rect 513234 514894 513854 550338
rect 514155 549132 514221 549133
rect 514155 549068 514156 549132
rect 514220 549068 514221 549132
rect 514155 549067 514221 549068
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 512499 482220 512565 482221
rect 512499 482156 512500 482220
rect 512564 482156 512565 482220
rect 512499 482155 512565 482156
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 512315 472836 512381 472837
rect 512315 472772 512316 472836
rect 512380 472772 512381 472836
rect 512315 472771 512381 472772
rect 513234 442894 513854 478338
rect 514158 473925 514218 549067
rect 514339 539204 514405 539205
rect 514339 539140 514340 539204
rect 514404 539140 514405 539204
rect 514339 539139 514405 539140
rect 514342 525877 514402 539139
rect 514707 532812 514773 532813
rect 514707 532748 514708 532812
rect 514772 532748 514773 532812
rect 514707 532747 514773 532748
rect 514523 526148 514589 526149
rect 514523 526084 514524 526148
rect 514588 526084 514589 526148
rect 514523 526083 514589 526084
rect 514339 525876 514405 525877
rect 514339 525812 514340 525876
rect 514404 525812 514405 525876
rect 514339 525811 514405 525812
rect 514155 473924 514221 473925
rect 514155 473860 514156 473924
rect 514220 473860 514221 473924
rect 514155 473859 514221 473860
rect 514526 470933 514586 526083
rect 514710 514725 514770 532747
rect 514891 527236 514957 527237
rect 514891 527172 514892 527236
rect 514956 527172 514957 527236
rect 514891 527171 514957 527172
rect 514707 514724 514773 514725
rect 514707 514660 514708 514724
rect 514772 514660 514773 514724
rect 514707 514659 514773 514660
rect 514707 505340 514773 505341
rect 514707 505276 514708 505340
rect 514772 505276 514773 505340
rect 514707 505275 514773 505276
rect 514523 470932 514589 470933
rect 514523 470868 514524 470932
rect 514588 470868 514589 470932
rect 514523 470867 514589 470868
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 512131 177852 512197 177853
rect 512131 177788 512132 177852
rect 512196 177788 512197 177852
rect 512131 177787 512197 177788
rect 510843 176220 510909 176221
rect 510843 176156 510844 176220
rect 510908 176156 510909 176220
rect 510843 176155 510909 176156
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -1306 510134 6618
rect 509514 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 510134 -1306
rect 509514 -1626 510134 -1542
rect 509514 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 510134 -1626
rect 509514 -7654 510134 -1862
rect 513234 154894 513854 190338
rect 514710 174453 514770 505275
rect 514894 180029 514954 527171
rect 515075 520300 515141 520301
rect 515075 520236 515076 520300
rect 515140 520236 515141 520300
rect 515075 520235 515141 520236
rect 514891 180028 514957 180029
rect 514891 179964 514892 180028
rect 514956 179964 514957 180028
rect 514891 179963 514957 179964
rect 515078 177581 515138 520235
rect 515262 470661 515322 558179
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516179 543420 516245 543421
rect 516179 543356 516180 543420
rect 516244 543356 516245 543420
rect 516179 543355 516245 543356
rect 515259 470660 515325 470661
rect 515259 470596 515260 470660
rect 515324 470596 515325 470660
rect 515259 470595 515325 470596
rect 516182 469845 516242 543355
rect 516363 519620 516429 519621
rect 516363 519556 516364 519620
rect 516428 519556 516429 519620
rect 516363 519555 516429 519556
rect 516366 478277 516426 519555
rect 516954 518614 517574 554058
rect 520674 594334 521294 600207
rect 520674 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 521294 594334
rect 520674 594014 521294 594098
rect 520674 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 521294 594014
rect 520674 558334 521294 593778
rect 524394 598054 525014 599988
rect 524394 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 525014 598054
rect 524394 597734 525014 597818
rect 524394 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 525014 597734
rect 524394 562054 525014 597498
rect 524394 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 525014 562054
rect 524394 561734 525014 561818
rect 524394 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 525014 561734
rect 523171 558516 523237 558517
rect 523171 558452 523172 558516
rect 523236 558452 523237 558516
rect 523171 558451 523237 558452
rect 520674 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 521294 558334
rect 520674 558014 521294 558098
rect 520674 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 521294 558014
rect 519307 547500 519373 547501
rect 519307 547436 519308 547500
rect 519372 547436 519373 547500
rect 519307 547435 519373 547436
rect 518387 536620 518453 536621
rect 518387 536556 518388 536620
rect 518452 536556 518453 536620
rect 518387 536555 518453 536556
rect 518019 527236 518085 527237
rect 518019 527172 518020 527236
rect 518084 527172 518085 527236
rect 518019 527171 518085 527172
rect 517835 523156 517901 523157
rect 517835 523092 517836 523156
rect 517900 523092 517901 523156
rect 517835 523091 517901 523092
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516363 478276 516429 478277
rect 516363 478212 516364 478276
rect 516428 478212 516429 478276
rect 516363 478211 516429 478212
rect 516179 469844 516245 469845
rect 516179 469780 516180 469844
rect 516244 469780 516245 469844
rect 516179 469779 516245 469780
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 515075 177580 515141 177581
rect 515075 177516 515076 177580
rect 515140 177516 515141 177580
rect 515075 177515 515141 177516
rect 514707 174452 514773 174453
rect 514707 174388 514708 174452
rect 514772 174388 514773 174452
rect 514707 174387 514773 174388
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -2266 513854 10338
rect 513234 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 513854 -2266
rect 513234 -2586 513854 -2502
rect 513234 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 513854 -2586
rect 513234 -7654 513854 -2822
rect 516954 158614 517574 194058
rect 517838 180165 517898 523091
rect 518022 262037 518082 527171
rect 518203 521796 518269 521797
rect 518203 521732 518204 521796
rect 518268 521732 518269 521796
rect 518203 521731 518269 521732
rect 518206 268021 518266 521731
rect 518390 481269 518450 536555
rect 518939 532812 519005 532813
rect 518939 532748 518940 532812
rect 519004 532748 519005 532812
rect 518939 532747 519005 532748
rect 518387 481268 518453 481269
rect 518387 481204 518388 481268
rect 518452 481204 518453 481268
rect 518387 481203 518453 481204
rect 518942 279989 519002 532747
rect 519123 523020 519189 523021
rect 519123 522956 519124 523020
rect 519188 522956 519189 523020
rect 519123 522955 519189 522956
rect 519126 435301 519186 522955
rect 519310 473381 519370 547435
rect 520411 537708 520477 537709
rect 520411 537644 520412 537708
rect 520476 537644 520477 537708
rect 520411 537643 520477 537644
rect 519491 536348 519557 536349
rect 519491 536284 519492 536348
rect 519556 536284 519557 536348
rect 519491 536283 519557 536284
rect 519494 478549 519554 536283
rect 520227 522884 520293 522885
rect 520227 522820 520228 522884
rect 520292 522820 520293 522884
rect 520227 522819 520293 522820
rect 519491 478548 519557 478549
rect 519491 478484 519492 478548
rect 519556 478484 519557 478548
rect 519491 478483 519557 478484
rect 519307 473380 519373 473381
rect 519307 473316 519308 473380
rect 519372 473316 519373 473380
rect 519307 473315 519373 473316
rect 519123 435300 519189 435301
rect 519123 435236 519124 435300
rect 519188 435236 519189 435300
rect 519123 435235 519189 435236
rect 520230 435029 520290 522819
rect 520414 473109 520474 537643
rect 520674 522334 521294 557778
rect 522987 554844 523053 554845
rect 522987 554780 522988 554844
rect 523052 554780 523053 554844
rect 522987 554779 523053 554780
rect 521699 539748 521765 539749
rect 521699 539684 521700 539748
rect 521764 539684 521765 539748
rect 521699 539683 521765 539684
rect 520674 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 521294 522334
rect 520674 522014 521294 522098
rect 520674 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 521294 522014
rect 520674 486334 521294 521778
rect 520674 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 521294 486334
rect 520674 486014 521294 486098
rect 520674 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 521294 486014
rect 520411 473108 520477 473109
rect 520411 473044 520412 473108
rect 520476 473044 520477 473108
rect 520411 473043 520477 473044
rect 520674 450334 521294 485778
rect 520674 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 521294 450334
rect 520674 450014 521294 450098
rect 520674 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 521294 450014
rect 520227 435028 520293 435029
rect 520227 434964 520228 435028
rect 520292 434964 520293 435028
rect 520227 434963 520293 434964
rect 520674 414334 521294 449778
rect 520674 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 521294 414334
rect 520674 414014 521294 414098
rect 520674 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 521294 414014
rect 520674 378334 521294 413778
rect 520674 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 521294 378334
rect 520674 378014 521294 378098
rect 520674 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 521294 378014
rect 520674 342334 521294 377778
rect 520674 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 521294 342334
rect 520674 342014 521294 342098
rect 520674 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 521294 342014
rect 520674 306334 521294 341778
rect 520674 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 521294 306334
rect 520674 306014 521294 306098
rect 520674 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 521294 306014
rect 518939 279988 519005 279989
rect 518939 279924 518940 279988
rect 519004 279924 519005 279988
rect 518939 279923 519005 279924
rect 520674 270334 521294 305778
rect 520674 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 521294 270334
rect 520674 270014 521294 270098
rect 520674 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 521294 270014
rect 518203 268020 518269 268021
rect 518203 267956 518204 268020
rect 518268 267956 518269 268020
rect 518203 267955 518269 267956
rect 518019 262036 518085 262037
rect 518019 261972 518020 262036
rect 518084 261972 518085 262036
rect 518019 261971 518085 261972
rect 520674 234334 521294 269778
rect 520674 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 521294 234334
rect 520674 234014 521294 234098
rect 520674 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 521294 234014
rect 520674 198334 521294 233778
rect 520674 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 521294 198334
rect 520674 198014 521294 198098
rect 520674 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 521294 198014
rect 517835 180164 517901 180165
rect 517835 180100 517836 180164
rect 517900 180100 517901 180164
rect 517835 180099 517901 180100
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 516954 -3226 517574 14058
rect 516954 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 517574 -3226
rect 516954 -3546 517574 -3462
rect 516954 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 517574 -3546
rect 516954 -7654 517574 -3782
rect 520674 162334 521294 197778
rect 521702 177717 521762 539683
rect 521883 539612 521949 539613
rect 521883 539548 521884 539612
rect 521948 539548 521949 539612
rect 521883 539547 521949 539548
rect 521886 309909 521946 539547
rect 522067 531452 522133 531453
rect 522067 531388 522068 531452
rect 522132 531388 522133 531452
rect 522067 531387 522133 531388
rect 522070 315893 522130 531387
rect 522251 519484 522317 519485
rect 522251 519420 522252 519484
rect 522316 519420 522317 519484
rect 522251 519419 522317 519420
rect 522254 484805 522314 519419
rect 522251 484804 522317 484805
rect 522251 484740 522252 484804
rect 522316 484740 522317 484804
rect 522251 484739 522317 484740
rect 522067 315892 522133 315893
rect 522067 315828 522068 315892
rect 522132 315828 522133 315892
rect 522067 315827 522133 315828
rect 521883 309908 521949 309909
rect 521883 309844 521884 309908
rect 521948 309844 521949 309908
rect 521883 309843 521949 309844
rect 522990 177989 523050 554779
rect 523174 470117 523234 558451
rect 523539 527236 523605 527237
rect 523539 527172 523540 527236
rect 523604 527172 523605 527236
rect 523539 527171 523605 527172
rect 523171 470116 523237 470117
rect 523171 470052 523172 470116
rect 523236 470052 523237 470116
rect 523171 470051 523237 470052
rect 523542 467941 523602 527171
rect 524394 526054 525014 561498
rect 528114 565774 528734 600207
rect 528114 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 528734 565774
rect 528114 565454 528734 565538
rect 528114 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 528734 565454
rect 525379 557156 525445 557157
rect 525379 557092 525380 557156
rect 525444 557092 525445 557156
rect 525379 557091 525445 557092
rect 524394 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 525014 526054
rect 524394 525734 525014 525818
rect 524394 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 525014 525734
rect 524394 490054 525014 525498
rect 525195 522612 525261 522613
rect 525195 522548 525196 522612
rect 525260 522548 525261 522612
rect 525195 522547 525261 522548
rect 524394 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 525014 490054
rect 524394 489734 525014 489818
rect 524394 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 525014 489734
rect 523539 467940 523605 467941
rect 523539 467876 523540 467940
rect 523604 467876 523605 467940
rect 523539 467875 523605 467876
rect 524394 454054 525014 489498
rect 524394 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 525014 454054
rect 524394 453734 525014 453818
rect 524394 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 525014 453734
rect 524394 418054 525014 453498
rect 525198 436117 525258 522547
rect 525382 476373 525442 557091
rect 526115 536484 526181 536485
rect 526115 536420 526116 536484
rect 526180 536420 526181 536484
rect 526115 536419 526181 536420
rect 525747 531452 525813 531453
rect 525747 531388 525748 531452
rect 525812 531388 525813 531452
rect 525747 531387 525813 531388
rect 525379 476372 525445 476373
rect 525379 476308 525380 476372
rect 525444 476308 525445 476372
rect 525379 476307 525445 476308
rect 525195 436116 525261 436117
rect 525195 436052 525196 436116
rect 525260 436052 525261 436116
rect 525195 436051 525261 436052
rect 524394 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 525014 418054
rect 524394 417734 525014 417818
rect 524394 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 525014 417734
rect 524394 382054 525014 417498
rect 524394 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 525014 382054
rect 524394 381734 525014 381818
rect 524394 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 525014 381734
rect 524394 346054 525014 381498
rect 524394 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 525014 346054
rect 524394 345734 525014 345818
rect 524394 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 525014 345734
rect 524394 310054 525014 345498
rect 524394 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 525014 310054
rect 524394 309734 525014 309818
rect 524394 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 525014 309734
rect 524394 274054 525014 309498
rect 524394 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 525014 274054
rect 524394 273734 525014 273818
rect 524394 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 525014 273734
rect 524394 238054 525014 273498
rect 524394 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 525014 238054
rect 524394 237734 525014 237818
rect 524394 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 525014 237734
rect 524394 202054 525014 237498
rect 524394 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 525014 202054
rect 524394 201734 525014 201818
rect 524394 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 525014 201734
rect 522987 177988 523053 177989
rect 522987 177924 522988 177988
rect 523052 177924 523053 177988
rect 522987 177923 523053 177924
rect 521699 177716 521765 177717
rect 521699 177652 521700 177716
rect 521764 177652 521765 177716
rect 521699 177651 521765 177652
rect 520674 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 521294 162334
rect 520674 162014 521294 162098
rect 520674 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 521294 162014
rect 520674 126334 521294 161778
rect 520674 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 521294 126334
rect 520674 126014 521294 126098
rect 520674 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 521294 126014
rect 520674 90334 521294 125778
rect 520674 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 521294 90334
rect 520674 90014 521294 90098
rect 520674 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 521294 90014
rect 520674 54334 521294 89778
rect 520674 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 521294 54334
rect 520674 54014 521294 54098
rect 520674 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 521294 54014
rect 520674 18334 521294 53778
rect 520674 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 521294 18334
rect 520674 18014 521294 18098
rect 520674 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 521294 18014
rect 520674 -4186 521294 17778
rect 520674 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 521294 -4186
rect 520674 -4506 521294 -4422
rect 520674 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 521294 -4506
rect 520674 -7654 521294 -4742
rect 524394 166054 525014 201498
rect 525750 180573 525810 531387
rect 525931 523156 525997 523157
rect 525931 523092 525932 523156
rect 525996 523092 525997 523156
rect 525931 523091 525997 523092
rect 525747 180572 525813 180573
rect 525747 180508 525748 180572
rect 525812 180508 525813 180572
rect 525747 180507 525813 180508
rect 525934 177445 525994 523091
rect 526118 470389 526178 536419
rect 528114 529774 528734 565218
rect 531834 569494 532454 600207
rect 533291 598092 533357 598093
rect 533291 598028 533292 598092
rect 533356 598028 533357 598092
rect 533291 598027 533357 598028
rect 534579 598092 534645 598093
rect 534579 598028 534580 598092
rect 534644 598028 534645 598092
rect 534579 598027 534645 598028
rect 531834 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 532454 569494
rect 531834 569174 532454 569258
rect 531834 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 532454 569174
rect 529059 548996 529125 548997
rect 529059 548932 529060 548996
rect 529124 548932 529125 548996
rect 529059 548931 529125 548932
rect 528114 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 528734 529774
rect 528114 529454 528734 529538
rect 528114 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 528734 529454
rect 527403 524244 527469 524245
rect 527403 524180 527404 524244
rect 527468 524180 527469 524244
rect 527403 524179 527469 524180
rect 527219 521252 527285 521253
rect 527219 521188 527220 521252
rect 527284 521188 527285 521252
rect 527219 521187 527285 521188
rect 526299 519756 526365 519757
rect 526299 519692 526300 519756
rect 526364 519692 526365 519756
rect 526299 519691 526365 519692
rect 526302 480861 526362 519691
rect 526299 480860 526365 480861
rect 526299 480796 526300 480860
rect 526364 480796 526365 480860
rect 526299 480795 526365 480796
rect 526115 470388 526181 470389
rect 526115 470324 526116 470388
rect 526180 470324 526181 470388
rect 526115 470323 526181 470324
rect 525931 177444 525997 177445
rect 525931 177380 525932 177444
rect 525996 177380 525997 177444
rect 525931 177379 525997 177380
rect 527222 176493 527282 521187
rect 527406 477733 527466 524179
rect 528114 493774 528734 529218
rect 528114 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 528734 493774
rect 528114 493454 528734 493538
rect 528114 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 528734 493454
rect 527403 477732 527469 477733
rect 527403 477668 527404 477732
rect 527468 477668 527469 477732
rect 527403 477667 527469 477668
rect 528114 457774 528734 493218
rect 529062 473653 529122 548931
rect 531834 533494 532454 568938
rect 532739 542060 532805 542061
rect 532739 541996 532740 542060
rect 532804 541996 532805 542060
rect 532739 541995 532805 541996
rect 531834 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 532454 533494
rect 531834 533174 532454 533258
rect 531834 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 532454 533174
rect 529979 531452 530045 531453
rect 529979 531388 529980 531452
rect 530044 531388 530045 531452
rect 529979 531387 530045 531388
rect 529243 520028 529309 520029
rect 529243 519964 529244 520028
rect 529308 519964 529309 520028
rect 529243 519963 529309 519964
rect 529246 481541 529306 519963
rect 529243 481540 529309 481541
rect 529243 481476 529244 481540
rect 529308 481476 529309 481540
rect 529243 481475 529309 481476
rect 529059 473652 529125 473653
rect 529059 473588 529060 473652
rect 529124 473588 529125 473652
rect 529059 473587 529125 473588
rect 528114 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 528734 457774
rect 528114 457454 528734 457538
rect 528114 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 528734 457454
rect 528114 421774 528734 457218
rect 528114 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 528734 421774
rect 528114 421454 528734 421538
rect 528114 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 528734 421454
rect 528114 385774 528734 421218
rect 528114 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 528734 385774
rect 528114 385454 528734 385538
rect 528114 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 528734 385454
rect 528114 349774 528734 385218
rect 528114 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 528734 349774
rect 528114 349454 528734 349538
rect 528114 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 528734 349454
rect 528114 313774 528734 349218
rect 528114 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 528734 313774
rect 528114 313454 528734 313538
rect 528114 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 528734 313454
rect 528114 277774 528734 313218
rect 528114 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 528734 277774
rect 528114 277454 528734 277538
rect 528114 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 528734 277454
rect 528114 241774 528734 277218
rect 528114 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 528734 241774
rect 528114 241454 528734 241538
rect 528114 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 528734 241454
rect 528114 205774 528734 241218
rect 528114 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 528734 205774
rect 528114 205454 528734 205538
rect 528114 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 528734 205454
rect 527219 176492 527285 176493
rect 527219 176428 527220 176492
rect 527284 176428 527285 176492
rect 527219 176427 527285 176428
rect 524394 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 525014 166054
rect 524394 165734 525014 165818
rect 524394 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 525014 165734
rect 524394 130054 525014 165498
rect 524394 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 525014 130054
rect 524394 129734 525014 129818
rect 524394 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 525014 129734
rect 524394 94054 525014 129498
rect 524394 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 525014 94054
rect 524394 93734 525014 93818
rect 524394 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 525014 93734
rect 524394 58054 525014 93498
rect 524394 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 525014 58054
rect 524394 57734 525014 57818
rect 524394 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 525014 57734
rect 524394 22054 525014 57498
rect 524394 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 525014 22054
rect 524394 21734 525014 21818
rect 524394 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 525014 21734
rect 524394 -5146 525014 21498
rect 524394 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 525014 -5146
rect 524394 -5466 525014 -5382
rect 524394 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 525014 -5466
rect 524394 -7654 525014 -5702
rect 528114 169774 528734 205218
rect 529982 180301 530042 531387
rect 530163 525332 530229 525333
rect 530163 525268 530164 525332
rect 530228 525268 530229 525332
rect 530163 525267 530229 525268
rect 530166 474741 530226 525267
rect 530531 521660 530597 521661
rect 530531 521596 530532 521660
rect 530596 521596 530597 521660
rect 530531 521595 530597 521596
rect 530163 474740 530229 474741
rect 530163 474676 530164 474740
rect 530228 474676 530229 474740
rect 530163 474675 530229 474676
rect 530534 356013 530594 521595
rect 531451 520980 531517 520981
rect 531451 520916 531452 520980
rect 531516 520916 531517 520980
rect 531451 520915 531517 520916
rect 531454 474469 531514 520915
rect 531834 497494 532454 532938
rect 531834 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 532454 497494
rect 531834 497174 532454 497258
rect 531834 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 532454 497174
rect 531451 474468 531517 474469
rect 531451 474404 531452 474468
rect 531516 474404 531517 474468
rect 531451 474403 531517 474404
rect 531834 461494 532454 496938
rect 532742 477461 532802 541995
rect 532739 477460 532805 477461
rect 532739 477396 532740 477460
rect 532804 477396 532805 477460
rect 532739 477395 532805 477396
rect 531834 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 532454 461494
rect 531834 461174 532454 461258
rect 531834 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 532454 461174
rect 531834 425494 532454 460938
rect 531834 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 532454 425494
rect 531834 425174 532454 425258
rect 531834 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 532454 425174
rect 531834 389494 532454 424938
rect 531834 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 532454 389494
rect 531834 389174 532454 389258
rect 531834 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 532454 389174
rect 530531 356012 530597 356013
rect 530531 355948 530532 356012
rect 530596 355948 530597 356012
rect 530531 355947 530597 355948
rect 531834 353494 532454 388938
rect 533294 356013 533354 598027
rect 534027 537844 534093 537845
rect 534027 537780 534028 537844
rect 534092 537780 534093 537844
rect 534027 537779 534093 537780
rect 534030 476917 534090 537779
rect 534027 476916 534093 476917
rect 534027 476852 534028 476916
rect 534092 476852 534093 476916
rect 534027 476851 534093 476852
rect 534582 356013 534642 598027
rect 535499 535532 535565 535533
rect 535499 535468 535500 535532
rect 535564 535468 535565 535532
rect 535499 535467 535565 535468
rect 533291 356012 533357 356013
rect 533291 355948 533292 356012
rect 533356 355948 533357 356012
rect 533291 355947 533357 355948
rect 534579 356012 534645 356013
rect 534579 355948 534580 356012
rect 534644 355948 534645 356012
rect 534579 355947 534645 355948
rect 531834 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 532454 353494
rect 531834 353174 532454 353258
rect 531834 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 532454 353174
rect 531834 317494 532454 352938
rect 531834 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 532454 317494
rect 531834 317174 532454 317258
rect 531834 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 532454 317174
rect 531834 281494 532454 316938
rect 531834 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 532454 281494
rect 531834 281174 532454 281258
rect 531834 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 532454 281174
rect 531834 245494 532454 280938
rect 531834 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 532454 245494
rect 531834 245174 532454 245258
rect 531834 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 532454 245174
rect 531834 209494 532454 244938
rect 531834 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 532454 209494
rect 531834 209174 532454 209258
rect 531834 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 532454 209174
rect 529979 180300 530045 180301
rect 529979 180236 529980 180300
rect 530044 180236 530045 180300
rect 529979 180235 530045 180236
rect 528114 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 528734 169774
rect 528114 169454 528734 169538
rect 528114 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 528734 169454
rect 528114 133774 528734 169218
rect 528114 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 528734 133774
rect 528114 133454 528734 133538
rect 528114 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 528734 133454
rect 528114 97774 528734 133218
rect 528114 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 528734 97774
rect 528114 97454 528734 97538
rect 528114 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 528734 97454
rect 528114 61774 528734 97218
rect 528114 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 528734 61774
rect 528114 61454 528734 61538
rect 528114 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 528734 61454
rect 528114 25774 528734 61218
rect 528114 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 528734 25774
rect 528114 25454 528734 25538
rect 528114 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 528734 25454
rect 528114 -6106 528734 25218
rect 528114 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 528734 -6106
rect 528114 -6426 528734 -6342
rect 528114 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 528734 -6426
rect 528114 -7654 528734 -6662
rect 531834 173494 532454 208938
rect 535502 180437 535562 535467
rect 536787 528052 536853 528053
rect 536787 527988 536788 528052
rect 536852 527988 536853 528052
rect 536787 527987 536853 527988
rect 535683 525196 535749 525197
rect 535683 525132 535684 525196
rect 535748 525132 535749 525196
rect 535683 525131 535749 525132
rect 535686 471749 535746 525131
rect 535683 471748 535749 471749
rect 535683 471684 535684 471748
rect 535748 471684 535749 471748
rect 535683 471683 535749 471684
rect 536790 453525 536850 527987
rect 536971 523972 537037 523973
rect 536971 523908 536972 523972
rect 537036 523908 537037 523972
rect 536971 523907 537037 523908
rect 536974 474197 537034 523907
rect 536971 474196 537037 474197
rect 536971 474132 536972 474196
rect 537036 474132 537037 474196
rect 536971 474131 537037 474132
rect 536787 453524 536853 453525
rect 536787 453460 536788 453524
rect 536852 453460 536853 453524
rect 536787 453459 536853 453460
rect 538262 374781 538322 601699
rect 538811 600404 538877 600405
rect 538811 600340 538812 600404
rect 538876 600340 538877 600404
rect 538811 600339 538877 600340
rect 538443 520436 538509 520437
rect 538443 520372 538444 520436
rect 538508 520372 538509 520436
rect 538443 520371 538509 520372
rect 538446 472021 538506 520371
rect 538627 473244 538693 473245
rect 538627 473180 538628 473244
rect 538692 473180 538693 473244
rect 538627 473179 538693 473180
rect 538443 472020 538509 472021
rect 538443 471956 538444 472020
rect 538508 471956 538509 472020
rect 538443 471955 538509 471956
rect 538630 379405 538690 473179
rect 538814 388653 538874 600339
rect 538811 388652 538877 388653
rect 538811 388588 538812 388652
rect 538876 388588 538877 388652
rect 538811 388587 538877 388588
rect 538627 379404 538693 379405
rect 538627 379340 538628 379404
rect 538692 379340 538693 379404
rect 538627 379339 538693 379340
rect 538259 374780 538325 374781
rect 538259 374716 538260 374780
rect 538324 374716 538325 374780
rect 538259 374715 538325 374716
rect 539366 369069 539426 604963
rect 539547 603668 539613 603669
rect 539547 603604 539548 603668
rect 539612 603604 539613 603668
rect 539547 603603 539613 603604
rect 539550 600405 539610 603603
rect 539547 600404 539613 600405
rect 539547 600340 539548 600404
rect 539612 600340 539613 600404
rect 539547 600339 539613 600340
rect 539547 551716 539613 551717
rect 539547 551652 539548 551716
rect 539612 551652 539613 551716
rect 539547 551651 539613 551652
rect 539550 472565 539610 551651
rect 539731 541924 539797 541925
rect 539731 541860 539732 541924
rect 539796 541860 539797 541924
rect 539731 541859 539797 541860
rect 539734 476645 539794 541859
rect 539731 476644 539797 476645
rect 539731 476580 539732 476644
rect 539796 476580 539797 476644
rect 539731 476579 539797 476580
rect 539547 472564 539613 472565
rect 539547 472500 539548 472564
rect 539612 472500 539613 472564
rect 539547 472499 539613 472500
rect 541022 373421 541082 614483
rect 541203 611828 541269 611829
rect 541203 611764 541204 611828
rect 541268 611764 541269 611828
rect 541203 611763 541269 611764
rect 541019 373420 541085 373421
rect 541019 373356 541020 373420
rect 541084 373356 541085 373420
rect 541019 373355 541085 373356
rect 541206 370565 541266 611763
rect 541794 579454 542414 614898
rect 542859 613188 542925 613189
rect 542859 613124 542860 613188
rect 542924 613124 542925 613188
rect 542859 613123 542925 613124
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541203 370564 541269 370565
rect 541203 370500 541204 370564
rect 541268 370500 541269 370564
rect 541203 370499 541269 370500
rect 539363 369068 539429 369069
rect 539363 369004 539364 369068
rect 539428 369004 539429 369068
rect 539363 369003 539429 369004
rect 541794 363454 542414 398898
rect 542675 371380 542741 371381
rect 542675 371316 542676 371380
rect 542740 371316 542741 371380
rect 542675 371315 542741 371316
rect 542678 365261 542738 371315
rect 542862 367709 542922 613123
rect 543411 610468 543477 610469
rect 543411 610404 543412 610468
rect 543476 610404 543477 610468
rect 543411 610403 543477 610404
rect 543043 607748 543109 607749
rect 543043 607684 543044 607748
rect 543108 607684 543109 607748
rect 543043 607683 543109 607684
rect 542859 367708 542925 367709
rect 542859 367644 542860 367708
rect 542924 367644 542925 367708
rect 542859 367643 542925 367644
rect 542675 365260 542741 365261
rect 542675 365196 542676 365260
rect 542740 365196 542741 365260
rect 542675 365195 542741 365196
rect 543046 363629 543106 607683
rect 543227 606388 543293 606389
rect 543227 606324 543228 606388
rect 543292 606324 543293 606388
rect 543227 606323 543293 606324
rect 543230 390285 543290 606323
rect 543227 390284 543293 390285
rect 543227 390220 543228 390284
rect 543292 390220 543293 390284
rect 543227 390219 543293 390220
rect 543227 389196 543293 389197
rect 543227 389132 543228 389196
rect 543292 389132 543293 389196
rect 543227 389131 543293 389132
rect 543230 372061 543290 389131
rect 543227 372060 543293 372061
rect 543227 371996 543228 372060
rect 543292 371996 543293 372060
rect 543227 371995 543293 371996
rect 543414 365397 543474 610403
rect 543782 384845 543842 621283
rect 545514 619174 546134 654618
rect 549234 706758 549854 711590
rect 549234 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 549854 706758
rect 549234 706438 549854 706522
rect 549234 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 549854 706438
rect 549234 694894 549854 706202
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 547643 647324 547709 647325
rect 547643 647260 547644 647324
rect 547708 647260 547709 647324
rect 547643 647259 547709 647260
rect 546539 619988 546605 619989
rect 546539 619924 546540 619988
rect 546604 619924 546605 619988
rect 546539 619923 546605 619924
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 544331 418300 544397 418301
rect 544331 418236 544332 418300
rect 544396 418236 544397 418300
rect 544331 418235 544397 418236
rect 543779 384844 543845 384845
rect 543779 384780 543780 384844
rect 543844 384780 543845 384844
rect 543779 384779 543845 384780
rect 543411 365396 543477 365397
rect 543411 365332 543412 365396
rect 543476 365332 543477 365396
rect 543411 365331 543477 365332
rect 543043 363628 543109 363629
rect 543043 363564 543044 363628
rect 543108 363564 543109 363628
rect 543043 363563 543109 363564
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 542859 276724 542925 276725
rect 542859 276660 542860 276724
rect 542924 276660 542925 276724
rect 542859 276659 542925 276660
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 535499 180436 535565 180437
rect 535499 180372 535500 180436
rect 535564 180372 535565 180436
rect 535499 180371 535565 180372
rect 531834 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 532454 173494
rect 531834 173174 532454 173258
rect 531834 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 532454 173174
rect 531834 137494 532454 172938
rect 531834 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 532454 137494
rect 531834 137174 532454 137258
rect 531834 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 532454 137174
rect 531834 101494 532454 136938
rect 531834 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 532454 101494
rect 531834 101174 532454 101258
rect 531834 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 532454 101174
rect 531834 65494 532454 100938
rect 531834 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 532454 65494
rect 531834 65174 532454 65258
rect 531834 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 532454 65174
rect 531834 29494 532454 64938
rect 531834 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 532454 29494
rect 531834 29174 532454 29258
rect 531834 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 532454 29174
rect 531834 -7066 532454 28938
rect 531834 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 532454 -7066
rect 531834 -7386 532454 -7302
rect 531834 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 532454 -7386
rect 531834 -7654 532454 -7622
rect 541794 147454 542414 182898
rect 542862 154325 542922 276659
rect 544334 155413 544394 418235
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 546542 384709 546602 619923
rect 547091 471476 547157 471477
rect 547091 471412 547092 471476
rect 547156 471412 547157 471476
rect 547091 471411 547157 471412
rect 546539 384708 546605 384709
rect 546539 384644 546540 384708
rect 546604 384644 546605 384708
rect 546539 384643 546605 384644
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 544331 155412 544397 155413
rect 544331 155348 544332 155412
rect 544396 155348 544397 155412
rect 544331 155347 544397 155348
rect 542859 154324 542925 154325
rect 542859 154260 542860 154324
rect 542924 154260 542925 154324
rect 542859 154259 542925 154260
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -7654 542414 -902
rect 545514 151174 546134 186618
rect 547094 155957 547154 471411
rect 547646 379405 547706 647259
rect 549234 622894 549854 658338
rect 552954 707718 553574 711590
rect 552954 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 553574 707718
rect 552954 707398 553574 707482
rect 552954 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 553574 707398
rect 552954 698614 553574 707162
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 550771 649908 550837 649909
rect 550771 649844 550772 649908
rect 550836 649844 550837 649908
rect 550771 649843 550837 649844
rect 550035 643108 550101 643109
rect 550035 643044 550036 643108
rect 550100 643044 550101 643108
rect 550035 643043 550101 643044
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 548379 524516 548445 524517
rect 548379 524452 548380 524516
rect 548444 524452 548445 524516
rect 548379 524451 548445 524452
rect 547643 379404 547709 379405
rect 547643 379340 547644 379404
rect 547708 379340 547709 379404
rect 547643 379339 547709 379340
rect 548382 156501 548442 524451
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 550038 381989 550098 643043
rect 550774 625170 550834 649843
rect 550590 625110 550834 625170
rect 552954 626614 553574 662058
rect 556674 708678 557294 711590
rect 556674 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 557294 708678
rect 556674 708358 557294 708442
rect 556674 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 557294 708358
rect 556674 666334 557294 708122
rect 560394 709638 561014 711590
rect 560394 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 561014 709638
rect 560394 709318 561014 709402
rect 560394 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 561014 709318
rect 558131 683908 558197 683909
rect 558131 683844 558132 683908
rect 558196 683844 558197 683908
rect 558131 683843 558197 683844
rect 556674 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 557294 666334
rect 556674 666014 557294 666098
rect 556674 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 557294 666014
rect 555371 630868 555437 630869
rect 555371 630804 555372 630868
rect 555436 630804 555437 630868
rect 555371 630803 555437 630804
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 550035 381988 550101 381989
rect 550035 381924 550036 381988
rect 550100 381924 550101 381988
rect 550035 381923 550101 381924
rect 550590 376549 550650 625110
rect 550771 624068 550837 624069
rect 550771 624004 550772 624068
rect 550836 624004 550837 624068
rect 550771 624003 550837 624004
rect 550774 381853 550834 624003
rect 550955 618628 551021 618629
rect 550955 618564 550956 618628
rect 551020 618564 551021 618628
rect 550955 618563 551021 618564
rect 550958 384573 551018 618563
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 551139 577692 551205 577693
rect 551139 577628 551140 577692
rect 551204 577628 551205 577692
rect 551139 577627 551205 577628
rect 550955 384572 551021 384573
rect 550955 384508 550956 384572
rect 551020 384508 551021 384572
rect 550955 384507 551021 384508
rect 550771 381852 550837 381853
rect 550771 381788 550772 381852
rect 550836 381788 550837 381852
rect 550771 381787 550837 381788
rect 550587 376548 550653 376549
rect 550587 376484 550588 376548
rect 550652 376484 550653 376548
rect 550587 376483 550653 376484
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 548379 156500 548445 156501
rect 548379 156436 548380 156500
rect 548444 156436 548445 156500
rect 548379 156435 548445 156436
rect 547091 155956 547157 155957
rect 547091 155892 547092 155956
rect 547156 155892 547157 155956
rect 547091 155891 547157 155892
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -1306 546134 6618
rect 545514 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 546134 -1306
rect 545514 -1626 546134 -1542
rect 545514 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 546134 -1626
rect 545514 -7654 546134 -1862
rect 549234 154894 549854 190338
rect 551142 157045 551202 577627
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 551139 157044 551205 157045
rect 551139 156980 551140 157044
rect 551204 156980 551205 157044
rect 551139 156979 551205 156980
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -2266 549854 10338
rect 549234 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 549854 -2266
rect 549234 -2586 549854 -2502
rect 549234 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 549854 -2586
rect 549234 -7654 549854 -2822
rect 552954 122614 553574 158058
rect 555374 157589 555434 630803
rect 556674 630334 557294 665778
rect 556674 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 557294 630334
rect 556674 630014 557294 630098
rect 556674 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 557294 630014
rect 556674 594334 557294 629778
rect 556674 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 557294 594334
rect 556674 594014 557294 594098
rect 556674 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 557294 594014
rect 556674 558334 557294 593778
rect 556674 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 557294 558334
rect 556674 558014 557294 558098
rect 556674 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 557294 558014
rect 556674 522334 557294 557778
rect 556674 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 557294 522334
rect 556674 522014 557294 522098
rect 556674 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 557294 522014
rect 556674 486334 557294 521778
rect 556674 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 557294 486334
rect 556674 486014 557294 486098
rect 556674 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 557294 486014
rect 556674 450334 557294 485778
rect 556674 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 557294 450334
rect 556674 450014 557294 450098
rect 556674 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 557294 450014
rect 556674 414334 557294 449778
rect 556674 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 557294 414334
rect 556674 414014 557294 414098
rect 556674 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 557294 414014
rect 556674 378334 557294 413778
rect 556674 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 557294 378334
rect 556674 378014 557294 378098
rect 556674 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 557294 378014
rect 556674 342334 557294 377778
rect 556674 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 557294 342334
rect 556674 342014 557294 342098
rect 556674 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 557294 342014
rect 556674 306334 557294 341778
rect 556674 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 557294 306334
rect 556674 306014 557294 306098
rect 556674 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 557294 306014
rect 556674 270334 557294 305778
rect 556674 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 557294 270334
rect 556674 270014 557294 270098
rect 556674 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 557294 270014
rect 556674 234334 557294 269778
rect 556674 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 557294 234334
rect 556674 234014 557294 234098
rect 556674 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 557294 234014
rect 556674 198334 557294 233778
rect 556674 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 557294 198334
rect 556674 198014 557294 198098
rect 556674 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 557294 198014
rect 556674 162334 557294 197778
rect 556674 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 557294 162334
rect 556674 162014 557294 162098
rect 556674 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 557294 162014
rect 555371 157588 555437 157589
rect 555371 157524 555372 157588
rect 555436 157524 555437 157588
rect 555371 157523 555437 157524
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 552954 -3226 553574 14058
rect 552954 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 553574 -3226
rect 552954 -3546 553574 -3462
rect 552954 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 553574 -3546
rect 552954 -7654 553574 -3782
rect 556674 126334 557294 161778
rect 558134 158133 558194 683843
rect 560394 670054 561014 709082
rect 560394 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 561014 670054
rect 560394 669734 561014 669818
rect 560394 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 561014 669734
rect 560394 634054 561014 669498
rect 560394 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 561014 634054
rect 560394 633734 561014 633818
rect 560394 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 561014 633734
rect 560394 598054 561014 633498
rect 560394 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 561014 598054
rect 560394 597734 561014 597818
rect 560394 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 561014 597734
rect 560394 562054 561014 597498
rect 560394 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 561014 562054
rect 560394 561734 561014 561818
rect 560394 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 561014 561734
rect 560394 526054 561014 561498
rect 560394 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 561014 526054
rect 560394 525734 561014 525818
rect 560394 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 561014 525734
rect 560394 490054 561014 525498
rect 560394 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 561014 490054
rect 560394 489734 561014 489818
rect 560394 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 561014 489734
rect 560394 454054 561014 489498
rect 560394 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 561014 454054
rect 560394 453734 561014 453818
rect 560394 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 561014 453734
rect 560394 418054 561014 453498
rect 560394 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 561014 418054
rect 560394 417734 561014 417818
rect 560394 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 561014 417734
rect 560394 382054 561014 417498
rect 560394 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 561014 382054
rect 560394 381734 561014 381818
rect 560394 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 561014 381734
rect 560394 346054 561014 381498
rect 560394 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 561014 346054
rect 560394 345734 561014 345818
rect 560394 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 561014 345734
rect 560394 310054 561014 345498
rect 560394 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 561014 310054
rect 560394 309734 561014 309818
rect 560394 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 561014 309734
rect 560394 274054 561014 309498
rect 560394 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 561014 274054
rect 560394 273734 561014 273818
rect 560394 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 561014 273734
rect 560394 238054 561014 273498
rect 560394 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 561014 238054
rect 560394 237734 561014 237818
rect 560394 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 561014 237734
rect 560394 202054 561014 237498
rect 560394 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 561014 202054
rect 560394 201734 561014 201818
rect 560394 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 561014 201734
rect 560394 166054 561014 201498
rect 560394 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 561014 166054
rect 560394 165734 561014 165818
rect 560394 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 561014 165734
rect 558131 158132 558197 158133
rect 558131 158068 558132 158132
rect 558196 158068 558197 158132
rect 558131 158067 558197 158068
rect 556674 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 557294 126334
rect 556674 126014 557294 126098
rect 556674 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 557294 126014
rect 556674 90334 557294 125778
rect 556674 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 557294 90334
rect 556674 90014 557294 90098
rect 556674 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 557294 90014
rect 556674 54334 557294 89778
rect 556674 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 557294 54334
rect 556674 54014 557294 54098
rect 556674 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 557294 54014
rect 556674 18334 557294 53778
rect 556674 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 557294 18334
rect 556674 18014 557294 18098
rect 556674 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 557294 18014
rect 556674 -4186 557294 17778
rect 556674 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 557294 -4186
rect 556674 -4506 557294 -4422
rect 556674 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 557294 -4506
rect 556674 -7654 557294 -4742
rect 560394 130054 561014 165498
rect 560394 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 561014 130054
rect 560394 129734 561014 129818
rect 560394 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 561014 129734
rect 560394 94054 561014 129498
rect 560394 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 561014 94054
rect 560394 93734 561014 93818
rect 560394 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 561014 93734
rect 560394 58054 561014 93498
rect 560394 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 561014 58054
rect 560394 57734 561014 57818
rect 560394 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 561014 57734
rect 560394 22054 561014 57498
rect 560394 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 561014 22054
rect 560394 21734 561014 21818
rect 560394 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 561014 21734
rect 560394 -5146 561014 21498
rect 560394 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 561014 -5146
rect 560394 -5466 561014 -5382
rect 560394 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 561014 -5466
rect 560394 -7654 561014 -5702
rect 564114 710598 564734 711590
rect 564114 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 564734 710598
rect 564114 710278 564734 710362
rect 564114 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 564734 710278
rect 564114 673774 564734 710042
rect 564114 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 564734 673774
rect 564114 673454 564734 673538
rect 564114 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 564734 673454
rect 564114 637774 564734 673218
rect 564114 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 564734 637774
rect 564114 637454 564734 637538
rect 564114 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 564734 637454
rect 564114 601774 564734 637218
rect 564114 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 564734 601774
rect 564114 601454 564734 601538
rect 564114 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 564734 601454
rect 564114 565774 564734 601218
rect 564114 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 564734 565774
rect 564114 565454 564734 565538
rect 564114 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 564734 565454
rect 564114 529774 564734 565218
rect 564114 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 564734 529774
rect 564114 529454 564734 529538
rect 564114 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 564734 529454
rect 564114 493774 564734 529218
rect 564114 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 564734 493774
rect 564114 493454 564734 493538
rect 564114 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 564734 493454
rect 564114 457774 564734 493218
rect 564114 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 564734 457774
rect 564114 457454 564734 457538
rect 564114 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 564734 457454
rect 564114 421774 564734 457218
rect 564114 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 564734 421774
rect 564114 421454 564734 421538
rect 564114 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 564734 421454
rect 564114 385774 564734 421218
rect 564114 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 564734 385774
rect 564114 385454 564734 385538
rect 564114 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 564734 385454
rect 564114 349774 564734 385218
rect 564114 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 564734 349774
rect 564114 349454 564734 349538
rect 564114 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 564734 349454
rect 564114 313774 564734 349218
rect 564114 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 564734 313774
rect 564114 313454 564734 313538
rect 564114 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 564734 313454
rect 564114 277774 564734 313218
rect 564114 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 564734 277774
rect 564114 277454 564734 277538
rect 564114 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 564734 277454
rect 564114 241774 564734 277218
rect 564114 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 564734 241774
rect 564114 241454 564734 241538
rect 564114 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 564734 241454
rect 564114 205774 564734 241218
rect 564114 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 564734 205774
rect 564114 205454 564734 205538
rect 564114 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 564734 205454
rect 564114 169774 564734 205218
rect 564114 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 564734 169774
rect 564114 169454 564734 169538
rect 564114 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 564734 169454
rect 564114 133774 564734 169218
rect 564114 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 564734 133774
rect 564114 133454 564734 133538
rect 564114 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 564734 133454
rect 564114 97774 564734 133218
rect 564114 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 564734 97774
rect 564114 97454 564734 97538
rect 564114 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 564734 97454
rect 564114 61774 564734 97218
rect 564114 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 564734 61774
rect 564114 61454 564734 61538
rect 564114 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 564734 61454
rect 564114 25774 564734 61218
rect 564114 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 564734 25774
rect 564114 25454 564734 25538
rect 564114 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 564734 25454
rect 564114 -6106 564734 25218
rect 564114 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 564734 -6106
rect 564114 -6426 564734 -6342
rect 564114 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 564734 -6426
rect 564114 -7654 564734 -6662
rect 567834 711558 568454 711590
rect 567834 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 568454 711558
rect 567834 711238 568454 711322
rect 567834 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 568454 711238
rect 567834 677494 568454 711002
rect 567834 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 568454 677494
rect 567834 677174 568454 677258
rect 567834 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 568454 677174
rect 567834 641494 568454 676938
rect 567834 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 568454 641494
rect 567834 641174 568454 641258
rect 567834 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 568454 641174
rect 567834 605494 568454 640938
rect 567834 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 568454 605494
rect 567834 605174 568454 605258
rect 567834 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 568454 605174
rect 567834 569494 568454 604938
rect 567834 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 568454 569494
rect 567834 569174 568454 569258
rect 567834 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 568454 569174
rect 567834 533494 568454 568938
rect 567834 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 568454 533494
rect 567834 533174 568454 533258
rect 567834 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 568454 533174
rect 567834 497494 568454 532938
rect 567834 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 568454 497494
rect 567834 497174 568454 497258
rect 567834 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 568454 497174
rect 567834 461494 568454 496938
rect 567834 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 568454 461494
rect 567834 461174 568454 461258
rect 567834 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 568454 461174
rect 567834 425494 568454 460938
rect 567834 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 568454 425494
rect 567834 425174 568454 425258
rect 567834 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 568454 425174
rect 567834 389494 568454 424938
rect 567834 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 568454 389494
rect 567834 389174 568454 389258
rect 567834 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 568454 389174
rect 567834 353494 568454 388938
rect 567834 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 568454 353494
rect 567834 353174 568454 353258
rect 567834 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 568454 353174
rect 567834 317494 568454 352938
rect 567834 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 568454 317494
rect 567834 317174 568454 317258
rect 567834 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 568454 317174
rect 567834 281494 568454 316938
rect 567834 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 568454 281494
rect 567834 281174 568454 281258
rect 567834 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 568454 281174
rect 567834 245494 568454 280938
rect 567834 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 568454 245494
rect 567834 245174 568454 245258
rect 567834 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 568454 245174
rect 567834 209494 568454 244938
rect 567834 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 568454 209494
rect 567834 209174 568454 209258
rect 567834 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 568454 209174
rect 567834 173494 568454 208938
rect 567834 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 568454 173494
rect 567834 173174 568454 173258
rect 567834 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 568454 173174
rect 567834 137494 568454 172938
rect 567834 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 568454 137494
rect 567834 137174 568454 137258
rect 567834 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 568454 137174
rect 567834 101494 568454 136938
rect 567834 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 568454 101494
rect 567834 101174 568454 101258
rect 567834 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 568454 101174
rect 567834 65494 568454 100938
rect 567834 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 568454 65494
rect 567834 65174 568454 65258
rect 567834 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 568454 65174
rect 567834 29494 568454 64938
rect 567834 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 568454 29494
rect 567834 29174 568454 29258
rect 567834 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 568454 29174
rect 567834 -7066 568454 28938
rect 567834 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 568454 -7066
rect 567834 -7386 568454 -7302
rect 567834 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 568454 -7386
rect 567834 -7654 568454 -7622
rect 577794 704838 578414 711590
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 581514 705798 582134 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 581514 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 582134 705798
rect 581514 705478 582134 705562
rect 581514 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 582134 705478
rect 581514 691174 582134 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 580211 591020 580277 591021
rect 580211 590956 580212 591020
rect 580276 590956 580277 591020
rect 580211 590955 580277 590956
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 580214 380221 580274 590955
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 580395 537844 580461 537845
rect 580395 537780 580396 537844
rect 580460 537780 580461 537844
rect 580395 537779 580461 537780
rect 580211 380220 580277 380221
rect 580211 380156 580212 380220
rect 580276 380156 580277 380220
rect 580211 380155 580277 380156
rect 580211 365124 580277 365125
rect 580211 365060 580212 365124
rect 580276 365060 580277 365124
rect 580211 365059 580277 365060
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 580214 162077 580274 365059
rect 580398 362269 580458 537779
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 580579 484668 580645 484669
rect 580579 484604 580580 484668
rect 580644 484604 580645 484668
rect 580579 484603 580645 484604
rect 580395 362268 580461 362269
rect 580395 362204 580396 362268
rect 580460 362204 580461 362268
rect 580395 362203 580461 362204
rect 580582 361045 580642 484603
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 580579 361044 580645 361045
rect 580579 360980 580580 361044
rect 580644 360980 580645 361044
rect 580579 360979 580645 360980
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 580395 312084 580461 312085
rect 580395 312020 580396 312084
rect 580460 312020 580461 312084
rect 580395 312019 580461 312020
rect 580398 276725 580458 312019
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 580395 276724 580461 276725
rect 580395 276660 580396 276724
rect 580460 276660 580461 276724
rect 580395 276659 580461 276660
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 580211 162076 580277 162077
rect 580211 162012 580212 162076
rect 580276 162012 580277 162076
rect 580211 162011 580277 162012
rect 581514 151174 582134 186618
rect 580211 151060 580277 151061
rect 580211 150996 580212 151060
rect 580276 150996 580277 151060
rect 580211 150995 580277 150996
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 580214 139365 580274 150995
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 580211 139364 580277 139365
rect 580211 139300 580212 139364
rect 580276 139300 580277 139364
rect 580211 139299 580277 139300
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 580211 112844 580277 112845
rect 580211 112780 580212 112844
rect 580276 112780 580277 112844
rect 580211 112779 580277 112780
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 580214 100741 580274 112779
rect 580211 100740 580277 100741
rect 580211 100676 580212 100740
rect 580276 100676 580277 100740
rect 580211 100675 580277 100676
rect 580211 98700 580277 98701
rect 580211 98636 580212 98700
rect 580276 98636 580277 98700
rect 580211 98635 580277 98636
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 580214 72997 580274 98635
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 580211 72996 580277 72997
rect 580211 72932 580212 72996
rect 580276 72932 580277 72996
rect 580211 72931 580277 72932
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -7654 578414 -902
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -1306 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 691174 586890 705242
rect 586270 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 586890 691174
rect 586270 690854 586890 690938
rect 586270 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 586890 690854
rect 586270 655174 586890 690618
rect 586270 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 586890 655174
rect 586270 654854 586890 654938
rect 586270 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 586890 654854
rect 586270 619174 586890 654618
rect 586270 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 586890 619174
rect 586270 618854 586890 618938
rect 586270 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 586890 618854
rect 586270 583174 586890 618618
rect 586270 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 586890 583174
rect 586270 582854 586890 582938
rect 586270 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 586890 582854
rect 586270 547174 586890 582618
rect 586270 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 586890 547174
rect 586270 546854 586890 546938
rect 586270 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 586890 546854
rect 586270 511174 586890 546618
rect 586270 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 586890 511174
rect 586270 510854 586890 510938
rect 586270 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 586890 510854
rect 586270 475174 586890 510618
rect 586270 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 586890 475174
rect 586270 474854 586890 474938
rect 586270 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 586890 474854
rect 586270 439174 586890 474618
rect 586270 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 586890 439174
rect 586270 438854 586890 438938
rect 586270 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 586890 438854
rect 586270 403174 586890 438618
rect 586270 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 586890 403174
rect 586270 402854 586890 402938
rect 586270 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 586890 402854
rect 586270 367174 586890 402618
rect 586270 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 586890 367174
rect 586270 366854 586890 366938
rect 586270 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 586890 366854
rect 586270 331174 586890 366618
rect 586270 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 586890 331174
rect 586270 330854 586890 330938
rect 586270 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 586890 330854
rect 586270 295174 586890 330618
rect 586270 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 586890 295174
rect 586270 294854 586890 294938
rect 586270 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 586890 294854
rect 586270 259174 586890 294618
rect 586270 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 586890 259174
rect 586270 258854 586890 258938
rect 586270 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 586890 258854
rect 586270 223174 586890 258618
rect 586270 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 586890 223174
rect 586270 222854 586890 222938
rect 586270 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 586890 222854
rect 586270 187174 586890 222618
rect 586270 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 586890 187174
rect 586270 186854 586890 186938
rect 586270 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 586890 186854
rect 586270 151174 586890 186618
rect 586270 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 586890 151174
rect 586270 150854 586890 150938
rect 586270 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 586890 150854
rect 586270 115174 586890 150618
rect 586270 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 586890 115174
rect 586270 114854 586890 114938
rect 586270 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 586890 114854
rect 586270 79174 586890 114618
rect 586270 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 586890 79174
rect 586270 78854 586890 78938
rect 586270 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 586890 78854
rect 586270 43174 586890 78618
rect 586270 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 586890 43174
rect 586270 42854 586890 42938
rect 586270 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 586890 42854
rect 586270 7174 586890 42618
rect 586270 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 586890 7174
rect 586270 6854 586890 6938
rect 586270 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 586890 6854
rect 581514 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 582134 -1306
rect 581514 -1626 582134 -1542
rect 581514 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 582134 -1626
rect 581514 -7654 582134 -1862
rect 586270 -1306 586890 6618
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 694894 587850 706202
rect 587230 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 587850 694894
rect 587230 694574 587850 694658
rect 587230 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 587850 694574
rect 587230 658894 587850 694338
rect 587230 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 587850 658894
rect 587230 658574 587850 658658
rect 587230 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 587850 658574
rect 587230 622894 587850 658338
rect 587230 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 587850 622894
rect 587230 622574 587850 622658
rect 587230 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 587850 622574
rect 587230 586894 587850 622338
rect 587230 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 587850 586894
rect 587230 586574 587850 586658
rect 587230 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 587850 586574
rect 587230 550894 587850 586338
rect 587230 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 587850 550894
rect 587230 550574 587850 550658
rect 587230 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 587850 550574
rect 587230 514894 587850 550338
rect 587230 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 587850 514894
rect 587230 514574 587850 514658
rect 587230 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 587850 514574
rect 587230 478894 587850 514338
rect 587230 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 587850 478894
rect 587230 478574 587850 478658
rect 587230 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 587850 478574
rect 587230 442894 587850 478338
rect 587230 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 587850 442894
rect 587230 442574 587850 442658
rect 587230 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 587850 442574
rect 587230 406894 587850 442338
rect 587230 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 587850 406894
rect 587230 406574 587850 406658
rect 587230 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 587850 406574
rect 587230 370894 587850 406338
rect 587230 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 587850 370894
rect 587230 370574 587850 370658
rect 587230 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 587850 370574
rect 587230 334894 587850 370338
rect 587230 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 587850 334894
rect 587230 334574 587850 334658
rect 587230 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 587850 334574
rect 587230 298894 587850 334338
rect 587230 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 587850 298894
rect 587230 298574 587850 298658
rect 587230 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 587850 298574
rect 587230 262894 587850 298338
rect 587230 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 587850 262894
rect 587230 262574 587850 262658
rect 587230 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 587850 262574
rect 587230 226894 587850 262338
rect 587230 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 587850 226894
rect 587230 226574 587850 226658
rect 587230 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 587850 226574
rect 587230 190894 587850 226338
rect 587230 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 587850 190894
rect 587230 190574 587850 190658
rect 587230 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 587850 190574
rect 587230 154894 587850 190338
rect 587230 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 587850 154894
rect 587230 154574 587850 154658
rect 587230 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 587850 154574
rect 587230 118894 587850 154338
rect 587230 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 587850 118894
rect 587230 118574 587850 118658
rect 587230 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 587850 118574
rect 587230 82894 587850 118338
rect 587230 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 587850 82894
rect 587230 82574 587850 82658
rect 587230 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 587850 82574
rect 587230 46894 587850 82338
rect 587230 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 587850 46894
rect 587230 46574 587850 46658
rect 587230 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 587850 46574
rect 587230 10894 587850 46338
rect 587230 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 587850 10894
rect 587230 10574 587850 10658
rect 587230 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 587850 10574
rect 587230 -2266 587850 10338
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 698614 588810 707162
rect 588190 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 588810 698614
rect 588190 698294 588810 698378
rect 588190 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 588810 698294
rect 588190 662614 588810 698058
rect 588190 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 588810 662614
rect 588190 662294 588810 662378
rect 588190 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 588810 662294
rect 588190 626614 588810 662058
rect 588190 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 588810 626614
rect 588190 626294 588810 626378
rect 588190 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 588810 626294
rect 588190 590614 588810 626058
rect 588190 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 588810 590614
rect 588190 590294 588810 590378
rect 588190 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 588810 590294
rect 588190 554614 588810 590058
rect 588190 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 588810 554614
rect 588190 554294 588810 554378
rect 588190 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 588810 554294
rect 588190 518614 588810 554058
rect 588190 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 588810 518614
rect 588190 518294 588810 518378
rect 588190 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 588810 518294
rect 588190 482614 588810 518058
rect 588190 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 588810 482614
rect 588190 482294 588810 482378
rect 588190 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 588810 482294
rect 588190 446614 588810 482058
rect 588190 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 588810 446614
rect 588190 446294 588810 446378
rect 588190 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 588810 446294
rect 588190 410614 588810 446058
rect 588190 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 588810 410614
rect 588190 410294 588810 410378
rect 588190 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 588810 410294
rect 588190 374614 588810 410058
rect 588190 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 588810 374614
rect 588190 374294 588810 374378
rect 588190 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 588810 374294
rect 588190 338614 588810 374058
rect 588190 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 588810 338614
rect 588190 338294 588810 338378
rect 588190 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 588810 338294
rect 588190 302614 588810 338058
rect 588190 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 588810 302614
rect 588190 302294 588810 302378
rect 588190 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 588810 302294
rect 588190 266614 588810 302058
rect 588190 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 588810 266614
rect 588190 266294 588810 266378
rect 588190 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 588810 266294
rect 588190 230614 588810 266058
rect 588190 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 588810 230614
rect 588190 230294 588810 230378
rect 588190 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 588810 230294
rect 588190 194614 588810 230058
rect 588190 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 588810 194614
rect 588190 194294 588810 194378
rect 588190 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 588810 194294
rect 588190 158614 588810 194058
rect 588190 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 588810 158614
rect 588190 158294 588810 158378
rect 588190 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 588810 158294
rect 588190 122614 588810 158058
rect 588190 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 588810 122614
rect 588190 122294 588810 122378
rect 588190 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 588810 122294
rect 588190 86614 588810 122058
rect 588190 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 588810 86614
rect 588190 86294 588810 86378
rect 588190 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 588810 86294
rect 588190 50614 588810 86058
rect 588190 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 588810 50614
rect 588190 50294 588810 50378
rect 588190 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 588810 50294
rect 588190 14614 588810 50058
rect 588190 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 588810 14614
rect 588190 14294 588810 14378
rect 588190 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 588810 14294
rect 588190 -3226 588810 14058
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 666334 589770 708122
rect 589150 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 589770 666334
rect 589150 666014 589770 666098
rect 589150 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 589770 666014
rect 589150 630334 589770 665778
rect 589150 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 589770 630334
rect 589150 630014 589770 630098
rect 589150 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 589770 630014
rect 589150 594334 589770 629778
rect 589150 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 589770 594334
rect 589150 594014 589770 594098
rect 589150 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 589770 594014
rect 589150 558334 589770 593778
rect 589150 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 589770 558334
rect 589150 558014 589770 558098
rect 589150 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 589770 558014
rect 589150 522334 589770 557778
rect 589150 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 589770 522334
rect 589150 522014 589770 522098
rect 589150 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 589770 522014
rect 589150 486334 589770 521778
rect 589150 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 589770 486334
rect 589150 486014 589770 486098
rect 589150 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 589770 486014
rect 589150 450334 589770 485778
rect 589150 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 589770 450334
rect 589150 450014 589770 450098
rect 589150 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 589770 450014
rect 589150 414334 589770 449778
rect 589150 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 589770 414334
rect 589150 414014 589770 414098
rect 589150 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 589770 414014
rect 589150 378334 589770 413778
rect 589150 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 589770 378334
rect 589150 378014 589770 378098
rect 589150 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 589770 378014
rect 589150 342334 589770 377778
rect 589150 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 589770 342334
rect 589150 342014 589770 342098
rect 589150 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 589770 342014
rect 589150 306334 589770 341778
rect 589150 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 589770 306334
rect 589150 306014 589770 306098
rect 589150 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 589770 306014
rect 589150 270334 589770 305778
rect 589150 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 589770 270334
rect 589150 270014 589770 270098
rect 589150 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 589770 270014
rect 589150 234334 589770 269778
rect 589150 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 589770 234334
rect 589150 234014 589770 234098
rect 589150 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 589770 234014
rect 589150 198334 589770 233778
rect 589150 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 589770 198334
rect 589150 198014 589770 198098
rect 589150 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 589770 198014
rect 589150 162334 589770 197778
rect 589150 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 589770 162334
rect 589150 162014 589770 162098
rect 589150 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 589770 162014
rect 589150 126334 589770 161778
rect 589150 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 589770 126334
rect 589150 126014 589770 126098
rect 589150 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 589770 126014
rect 589150 90334 589770 125778
rect 589150 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 589770 90334
rect 589150 90014 589770 90098
rect 589150 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 589770 90014
rect 589150 54334 589770 89778
rect 589150 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 589770 54334
rect 589150 54014 589770 54098
rect 589150 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 589770 54014
rect 589150 18334 589770 53778
rect 589150 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 589770 18334
rect 589150 18014 589770 18098
rect 589150 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 589770 18014
rect 589150 -4186 589770 17778
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 670054 590730 709082
rect 590110 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 590730 670054
rect 590110 669734 590730 669818
rect 590110 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 590730 669734
rect 590110 634054 590730 669498
rect 590110 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 590730 634054
rect 590110 633734 590730 633818
rect 590110 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 590730 633734
rect 590110 598054 590730 633498
rect 590110 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 590730 598054
rect 590110 597734 590730 597818
rect 590110 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 590730 597734
rect 590110 562054 590730 597498
rect 590110 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 590730 562054
rect 590110 561734 590730 561818
rect 590110 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 590730 561734
rect 590110 526054 590730 561498
rect 590110 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 590730 526054
rect 590110 525734 590730 525818
rect 590110 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 590730 525734
rect 590110 490054 590730 525498
rect 590110 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 590730 490054
rect 590110 489734 590730 489818
rect 590110 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 590730 489734
rect 590110 454054 590730 489498
rect 590110 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 590730 454054
rect 590110 453734 590730 453818
rect 590110 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 590730 453734
rect 590110 418054 590730 453498
rect 590110 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 590730 418054
rect 590110 417734 590730 417818
rect 590110 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 590730 417734
rect 590110 382054 590730 417498
rect 590110 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 590730 382054
rect 590110 381734 590730 381818
rect 590110 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 590730 381734
rect 590110 346054 590730 381498
rect 590110 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 590730 346054
rect 590110 345734 590730 345818
rect 590110 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 590730 345734
rect 590110 310054 590730 345498
rect 590110 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 590730 310054
rect 590110 309734 590730 309818
rect 590110 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 590730 309734
rect 590110 274054 590730 309498
rect 590110 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 590730 274054
rect 590110 273734 590730 273818
rect 590110 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 590730 273734
rect 590110 238054 590730 273498
rect 590110 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 590730 238054
rect 590110 237734 590730 237818
rect 590110 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 590730 237734
rect 590110 202054 590730 237498
rect 590110 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 590730 202054
rect 590110 201734 590730 201818
rect 590110 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 590730 201734
rect 590110 166054 590730 201498
rect 590110 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 590730 166054
rect 590110 165734 590730 165818
rect 590110 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 590730 165734
rect 590110 130054 590730 165498
rect 590110 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 590730 130054
rect 590110 129734 590730 129818
rect 590110 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 590730 129734
rect 590110 94054 590730 129498
rect 590110 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 590730 94054
rect 590110 93734 590730 93818
rect 590110 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 590730 93734
rect 590110 58054 590730 93498
rect 590110 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 590730 58054
rect 590110 57734 590730 57818
rect 590110 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 590730 57734
rect 590110 22054 590730 57498
rect 590110 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 590730 22054
rect 590110 21734 590730 21818
rect 590110 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 590730 21734
rect 590110 -5146 590730 21498
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 673774 591690 710042
rect 591070 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 591690 673774
rect 591070 673454 591690 673538
rect 591070 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 591690 673454
rect 591070 637774 591690 673218
rect 591070 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 591690 637774
rect 591070 637454 591690 637538
rect 591070 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 591690 637454
rect 591070 601774 591690 637218
rect 591070 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 591690 601774
rect 591070 601454 591690 601538
rect 591070 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 591690 601454
rect 591070 565774 591690 601218
rect 591070 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 591690 565774
rect 591070 565454 591690 565538
rect 591070 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 591690 565454
rect 591070 529774 591690 565218
rect 591070 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 591690 529774
rect 591070 529454 591690 529538
rect 591070 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 591690 529454
rect 591070 493774 591690 529218
rect 591070 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 591690 493774
rect 591070 493454 591690 493538
rect 591070 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 591690 493454
rect 591070 457774 591690 493218
rect 591070 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 591690 457774
rect 591070 457454 591690 457538
rect 591070 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 591690 457454
rect 591070 421774 591690 457218
rect 591070 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 591690 421774
rect 591070 421454 591690 421538
rect 591070 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 591690 421454
rect 591070 385774 591690 421218
rect 591070 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 591690 385774
rect 591070 385454 591690 385538
rect 591070 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 591690 385454
rect 591070 349774 591690 385218
rect 591070 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 591690 349774
rect 591070 349454 591690 349538
rect 591070 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 591690 349454
rect 591070 313774 591690 349218
rect 591070 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 591690 313774
rect 591070 313454 591690 313538
rect 591070 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 591690 313454
rect 591070 277774 591690 313218
rect 591070 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 591690 277774
rect 591070 277454 591690 277538
rect 591070 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 591690 277454
rect 591070 241774 591690 277218
rect 591070 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 591690 241774
rect 591070 241454 591690 241538
rect 591070 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 591690 241454
rect 591070 205774 591690 241218
rect 591070 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 591690 205774
rect 591070 205454 591690 205538
rect 591070 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 591690 205454
rect 591070 169774 591690 205218
rect 591070 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 591690 169774
rect 591070 169454 591690 169538
rect 591070 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 591690 169454
rect 591070 133774 591690 169218
rect 591070 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 591690 133774
rect 591070 133454 591690 133538
rect 591070 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 591690 133454
rect 591070 97774 591690 133218
rect 591070 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 591690 97774
rect 591070 97454 591690 97538
rect 591070 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 591690 97454
rect 591070 61774 591690 97218
rect 591070 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 591690 61774
rect 591070 61454 591690 61538
rect 591070 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 591690 61454
rect 591070 25774 591690 61218
rect 591070 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 591690 25774
rect 591070 25454 591690 25538
rect 591070 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 591690 25454
rect 591070 -6106 591690 25218
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 677494 592650 711002
rect 592030 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect 592030 677174 592650 677258
rect 592030 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect 592030 641494 592650 676938
rect 592030 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect 592030 641174 592650 641258
rect 592030 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect 592030 605494 592650 640938
rect 592030 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect 592030 605174 592650 605258
rect 592030 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect 592030 569494 592650 604938
rect 592030 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect 592030 569174 592650 569258
rect 592030 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect 592030 533494 592650 568938
rect 592030 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect 592030 533174 592650 533258
rect 592030 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect 592030 497494 592650 532938
rect 592030 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect 592030 497174 592650 497258
rect 592030 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect 592030 461494 592650 496938
rect 592030 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect 592030 461174 592650 461258
rect 592030 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect 592030 425494 592650 460938
rect 592030 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect 592030 425174 592650 425258
rect 592030 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect 592030 389494 592650 424938
rect 592030 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect 592030 389174 592650 389258
rect 592030 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect 592030 353494 592650 388938
rect 592030 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect 592030 353174 592650 353258
rect 592030 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect 592030 317494 592650 352938
rect 592030 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect 592030 317174 592650 317258
rect 592030 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect 592030 281494 592650 316938
rect 592030 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect 592030 281174 592650 281258
rect 592030 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect 592030 245494 592650 280938
rect 592030 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect 592030 245174 592650 245258
rect 592030 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect 592030 209494 592650 244938
rect 592030 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect 592030 209174 592650 209258
rect 592030 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect 592030 173494 592650 208938
rect 592030 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect 592030 173174 592650 173258
rect 592030 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect 592030 137494 592650 172938
rect 592030 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect 592030 137174 592650 137258
rect 592030 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect 592030 101494 592650 136938
rect 592030 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect 592030 101174 592650 101258
rect 592030 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect 592030 65494 592650 100938
rect 592030 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect 592030 65174 592650 65258
rect 592030 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect 592030 29494 592650 64938
rect 592030 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect 592030 29174 592650 29258
rect 592030 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect 592030 -7066 592650 28938
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 677258 -8458 677494
rect -8374 677258 -8138 677494
rect -8694 676938 -8458 677174
rect -8374 676938 -8138 677174
rect -8694 641258 -8458 641494
rect -8374 641258 -8138 641494
rect -8694 640938 -8458 641174
rect -8374 640938 -8138 641174
rect -8694 605258 -8458 605494
rect -8374 605258 -8138 605494
rect -8694 604938 -8458 605174
rect -8374 604938 -8138 605174
rect -8694 569258 -8458 569494
rect -8374 569258 -8138 569494
rect -8694 568938 -8458 569174
rect -8374 568938 -8138 569174
rect -8694 533258 -8458 533494
rect -8374 533258 -8138 533494
rect -8694 532938 -8458 533174
rect -8374 532938 -8138 533174
rect -8694 497258 -8458 497494
rect -8374 497258 -8138 497494
rect -8694 496938 -8458 497174
rect -8374 496938 -8138 497174
rect -8694 461258 -8458 461494
rect -8374 461258 -8138 461494
rect -8694 460938 -8458 461174
rect -8374 460938 -8138 461174
rect -8694 425258 -8458 425494
rect -8374 425258 -8138 425494
rect -8694 424938 -8458 425174
rect -8374 424938 -8138 425174
rect -8694 389258 -8458 389494
rect -8374 389258 -8138 389494
rect -8694 388938 -8458 389174
rect -8374 388938 -8138 389174
rect -8694 353258 -8458 353494
rect -8374 353258 -8138 353494
rect -8694 352938 -8458 353174
rect -8374 352938 -8138 353174
rect -8694 317258 -8458 317494
rect -8374 317258 -8138 317494
rect -8694 316938 -8458 317174
rect -8374 316938 -8138 317174
rect -8694 281258 -8458 281494
rect -8374 281258 -8138 281494
rect -8694 280938 -8458 281174
rect -8374 280938 -8138 281174
rect -8694 245258 -8458 245494
rect -8374 245258 -8138 245494
rect -8694 244938 -8458 245174
rect -8374 244938 -8138 245174
rect -8694 209258 -8458 209494
rect -8374 209258 -8138 209494
rect -8694 208938 -8458 209174
rect -8374 208938 -8138 209174
rect -8694 173258 -8458 173494
rect -8374 173258 -8138 173494
rect -8694 172938 -8458 173174
rect -8374 172938 -8138 173174
rect -8694 137258 -8458 137494
rect -8374 137258 -8138 137494
rect -8694 136938 -8458 137174
rect -8374 136938 -8138 137174
rect -8694 101258 -8458 101494
rect -8374 101258 -8138 101494
rect -8694 100938 -8458 101174
rect -8374 100938 -8138 101174
rect -8694 65258 -8458 65494
rect -8374 65258 -8138 65494
rect -8694 64938 -8458 65174
rect -8374 64938 -8138 65174
rect -8694 29258 -8458 29494
rect -8374 29258 -8138 29494
rect -8694 28938 -8458 29174
rect -8374 28938 -8138 29174
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -7734 673538 -7498 673774
rect -7414 673538 -7178 673774
rect -7734 673218 -7498 673454
rect -7414 673218 -7178 673454
rect -7734 637538 -7498 637774
rect -7414 637538 -7178 637774
rect -7734 637218 -7498 637454
rect -7414 637218 -7178 637454
rect -7734 601538 -7498 601774
rect -7414 601538 -7178 601774
rect -7734 601218 -7498 601454
rect -7414 601218 -7178 601454
rect -7734 565538 -7498 565774
rect -7414 565538 -7178 565774
rect -7734 565218 -7498 565454
rect -7414 565218 -7178 565454
rect -7734 529538 -7498 529774
rect -7414 529538 -7178 529774
rect -7734 529218 -7498 529454
rect -7414 529218 -7178 529454
rect -7734 493538 -7498 493774
rect -7414 493538 -7178 493774
rect -7734 493218 -7498 493454
rect -7414 493218 -7178 493454
rect -7734 457538 -7498 457774
rect -7414 457538 -7178 457774
rect -7734 457218 -7498 457454
rect -7414 457218 -7178 457454
rect -7734 421538 -7498 421774
rect -7414 421538 -7178 421774
rect -7734 421218 -7498 421454
rect -7414 421218 -7178 421454
rect -7734 385538 -7498 385774
rect -7414 385538 -7178 385774
rect -7734 385218 -7498 385454
rect -7414 385218 -7178 385454
rect -7734 349538 -7498 349774
rect -7414 349538 -7178 349774
rect -7734 349218 -7498 349454
rect -7414 349218 -7178 349454
rect -7734 313538 -7498 313774
rect -7414 313538 -7178 313774
rect -7734 313218 -7498 313454
rect -7414 313218 -7178 313454
rect -7734 277538 -7498 277774
rect -7414 277538 -7178 277774
rect -7734 277218 -7498 277454
rect -7414 277218 -7178 277454
rect -7734 241538 -7498 241774
rect -7414 241538 -7178 241774
rect -7734 241218 -7498 241454
rect -7414 241218 -7178 241454
rect -7734 205538 -7498 205774
rect -7414 205538 -7178 205774
rect -7734 205218 -7498 205454
rect -7414 205218 -7178 205454
rect -7734 169538 -7498 169774
rect -7414 169538 -7178 169774
rect -7734 169218 -7498 169454
rect -7414 169218 -7178 169454
rect -7734 133538 -7498 133774
rect -7414 133538 -7178 133774
rect -7734 133218 -7498 133454
rect -7414 133218 -7178 133454
rect -7734 97538 -7498 97774
rect -7414 97538 -7178 97774
rect -7734 97218 -7498 97454
rect -7414 97218 -7178 97454
rect -7734 61538 -7498 61774
rect -7414 61538 -7178 61774
rect -7734 61218 -7498 61454
rect -7414 61218 -7178 61454
rect -7734 25538 -7498 25774
rect -7414 25538 -7178 25774
rect -7734 25218 -7498 25454
rect -7414 25218 -7178 25454
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 669818 -6538 670054
rect -6454 669818 -6218 670054
rect -6774 669498 -6538 669734
rect -6454 669498 -6218 669734
rect -6774 633818 -6538 634054
rect -6454 633818 -6218 634054
rect -6774 633498 -6538 633734
rect -6454 633498 -6218 633734
rect -6774 597818 -6538 598054
rect -6454 597818 -6218 598054
rect -6774 597498 -6538 597734
rect -6454 597498 -6218 597734
rect -6774 561818 -6538 562054
rect -6454 561818 -6218 562054
rect -6774 561498 -6538 561734
rect -6454 561498 -6218 561734
rect -6774 525818 -6538 526054
rect -6454 525818 -6218 526054
rect -6774 525498 -6538 525734
rect -6454 525498 -6218 525734
rect -6774 489818 -6538 490054
rect -6454 489818 -6218 490054
rect -6774 489498 -6538 489734
rect -6454 489498 -6218 489734
rect -6774 453818 -6538 454054
rect -6454 453818 -6218 454054
rect -6774 453498 -6538 453734
rect -6454 453498 -6218 453734
rect -6774 417818 -6538 418054
rect -6454 417818 -6218 418054
rect -6774 417498 -6538 417734
rect -6454 417498 -6218 417734
rect -6774 381818 -6538 382054
rect -6454 381818 -6218 382054
rect -6774 381498 -6538 381734
rect -6454 381498 -6218 381734
rect -6774 345818 -6538 346054
rect -6454 345818 -6218 346054
rect -6774 345498 -6538 345734
rect -6454 345498 -6218 345734
rect -6774 309818 -6538 310054
rect -6454 309818 -6218 310054
rect -6774 309498 -6538 309734
rect -6454 309498 -6218 309734
rect -6774 273818 -6538 274054
rect -6454 273818 -6218 274054
rect -6774 273498 -6538 273734
rect -6454 273498 -6218 273734
rect -6774 237818 -6538 238054
rect -6454 237818 -6218 238054
rect -6774 237498 -6538 237734
rect -6454 237498 -6218 237734
rect -6774 201818 -6538 202054
rect -6454 201818 -6218 202054
rect -6774 201498 -6538 201734
rect -6454 201498 -6218 201734
rect -6774 165818 -6538 166054
rect -6454 165818 -6218 166054
rect -6774 165498 -6538 165734
rect -6454 165498 -6218 165734
rect -6774 129818 -6538 130054
rect -6454 129818 -6218 130054
rect -6774 129498 -6538 129734
rect -6454 129498 -6218 129734
rect -6774 93818 -6538 94054
rect -6454 93818 -6218 94054
rect -6774 93498 -6538 93734
rect -6454 93498 -6218 93734
rect -6774 57818 -6538 58054
rect -6454 57818 -6218 58054
rect -6774 57498 -6538 57734
rect -6454 57498 -6218 57734
rect -6774 21818 -6538 22054
rect -6454 21818 -6218 22054
rect -6774 21498 -6538 21734
rect -6454 21498 -6218 21734
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -5814 666098 -5578 666334
rect -5494 666098 -5258 666334
rect -5814 665778 -5578 666014
rect -5494 665778 -5258 666014
rect -5814 630098 -5578 630334
rect -5494 630098 -5258 630334
rect -5814 629778 -5578 630014
rect -5494 629778 -5258 630014
rect -5814 594098 -5578 594334
rect -5494 594098 -5258 594334
rect -5814 593778 -5578 594014
rect -5494 593778 -5258 594014
rect -5814 558098 -5578 558334
rect -5494 558098 -5258 558334
rect -5814 557778 -5578 558014
rect -5494 557778 -5258 558014
rect -5814 522098 -5578 522334
rect -5494 522098 -5258 522334
rect -5814 521778 -5578 522014
rect -5494 521778 -5258 522014
rect -5814 486098 -5578 486334
rect -5494 486098 -5258 486334
rect -5814 485778 -5578 486014
rect -5494 485778 -5258 486014
rect -5814 450098 -5578 450334
rect -5494 450098 -5258 450334
rect -5814 449778 -5578 450014
rect -5494 449778 -5258 450014
rect -5814 414098 -5578 414334
rect -5494 414098 -5258 414334
rect -5814 413778 -5578 414014
rect -5494 413778 -5258 414014
rect -5814 378098 -5578 378334
rect -5494 378098 -5258 378334
rect -5814 377778 -5578 378014
rect -5494 377778 -5258 378014
rect -5814 342098 -5578 342334
rect -5494 342098 -5258 342334
rect -5814 341778 -5578 342014
rect -5494 341778 -5258 342014
rect -5814 306098 -5578 306334
rect -5494 306098 -5258 306334
rect -5814 305778 -5578 306014
rect -5494 305778 -5258 306014
rect -5814 270098 -5578 270334
rect -5494 270098 -5258 270334
rect -5814 269778 -5578 270014
rect -5494 269778 -5258 270014
rect -5814 234098 -5578 234334
rect -5494 234098 -5258 234334
rect -5814 233778 -5578 234014
rect -5494 233778 -5258 234014
rect -5814 198098 -5578 198334
rect -5494 198098 -5258 198334
rect -5814 197778 -5578 198014
rect -5494 197778 -5258 198014
rect -5814 162098 -5578 162334
rect -5494 162098 -5258 162334
rect -5814 161778 -5578 162014
rect -5494 161778 -5258 162014
rect -5814 126098 -5578 126334
rect -5494 126098 -5258 126334
rect -5814 125778 -5578 126014
rect -5494 125778 -5258 126014
rect -5814 90098 -5578 90334
rect -5494 90098 -5258 90334
rect -5814 89778 -5578 90014
rect -5494 89778 -5258 90014
rect -5814 54098 -5578 54334
rect -5494 54098 -5258 54334
rect -5814 53778 -5578 54014
rect -5494 53778 -5258 54014
rect -5814 18098 -5578 18334
rect -5494 18098 -5258 18334
rect -5814 17778 -5578 18014
rect -5494 17778 -5258 18014
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 698378 -4618 698614
rect -4534 698378 -4298 698614
rect -4854 698058 -4618 698294
rect -4534 698058 -4298 698294
rect -4854 662378 -4618 662614
rect -4534 662378 -4298 662614
rect -4854 662058 -4618 662294
rect -4534 662058 -4298 662294
rect -4854 626378 -4618 626614
rect -4534 626378 -4298 626614
rect -4854 626058 -4618 626294
rect -4534 626058 -4298 626294
rect -4854 590378 -4618 590614
rect -4534 590378 -4298 590614
rect -4854 590058 -4618 590294
rect -4534 590058 -4298 590294
rect -4854 554378 -4618 554614
rect -4534 554378 -4298 554614
rect -4854 554058 -4618 554294
rect -4534 554058 -4298 554294
rect -4854 518378 -4618 518614
rect -4534 518378 -4298 518614
rect -4854 518058 -4618 518294
rect -4534 518058 -4298 518294
rect -4854 482378 -4618 482614
rect -4534 482378 -4298 482614
rect -4854 482058 -4618 482294
rect -4534 482058 -4298 482294
rect -4854 446378 -4618 446614
rect -4534 446378 -4298 446614
rect -4854 446058 -4618 446294
rect -4534 446058 -4298 446294
rect -4854 410378 -4618 410614
rect -4534 410378 -4298 410614
rect -4854 410058 -4618 410294
rect -4534 410058 -4298 410294
rect -4854 374378 -4618 374614
rect -4534 374378 -4298 374614
rect -4854 374058 -4618 374294
rect -4534 374058 -4298 374294
rect -4854 338378 -4618 338614
rect -4534 338378 -4298 338614
rect -4854 338058 -4618 338294
rect -4534 338058 -4298 338294
rect -4854 302378 -4618 302614
rect -4534 302378 -4298 302614
rect -4854 302058 -4618 302294
rect -4534 302058 -4298 302294
rect -4854 266378 -4618 266614
rect -4534 266378 -4298 266614
rect -4854 266058 -4618 266294
rect -4534 266058 -4298 266294
rect -4854 230378 -4618 230614
rect -4534 230378 -4298 230614
rect -4854 230058 -4618 230294
rect -4534 230058 -4298 230294
rect -4854 194378 -4618 194614
rect -4534 194378 -4298 194614
rect -4854 194058 -4618 194294
rect -4534 194058 -4298 194294
rect -4854 158378 -4618 158614
rect -4534 158378 -4298 158614
rect -4854 158058 -4618 158294
rect -4534 158058 -4298 158294
rect -4854 122378 -4618 122614
rect -4534 122378 -4298 122614
rect -4854 122058 -4618 122294
rect -4534 122058 -4298 122294
rect -4854 86378 -4618 86614
rect -4534 86378 -4298 86614
rect -4854 86058 -4618 86294
rect -4534 86058 -4298 86294
rect -4854 50378 -4618 50614
rect -4534 50378 -4298 50614
rect -4854 50058 -4618 50294
rect -4534 50058 -4298 50294
rect -4854 14378 -4618 14614
rect -4534 14378 -4298 14614
rect -4854 14058 -4618 14294
rect -4534 14058 -4298 14294
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -3894 694658 -3658 694894
rect -3574 694658 -3338 694894
rect -3894 694338 -3658 694574
rect -3574 694338 -3338 694574
rect -3894 658658 -3658 658894
rect -3574 658658 -3338 658894
rect -3894 658338 -3658 658574
rect -3574 658338 -3338 658574
rect -3894 622658 -3658 622894
rect -3574 622658 -3338 622894
rect -3894 622338 -3658 622574
rect -3574 622338 -3338 622574
rect -3894 586658 -3658 586894
rect -3574 586658 -3338 586894
rect -3894 586338 -3658 586574
rect -3574 586338 -3338 586574
rect -3894 550658 -3658 550894
rect -3574 550658 -3338 550894
rect -3894 550338 -3658 550574
rect -3574 550338 -3338 550574
rect -3894 514658 -3658 514894
rect -3574 514658 -3338 514894
rect -3894 514338 -3658 514574
rect -3574 514338 -3338 514574
rect -3894 478658 -3658 478894
rect -3574 478658 -3338 478894
rect -3894 478338 -3658 478574
rect -3574 478338 -3338 478574
rect -3894 442658 -3658 442894
rect -3574 442658 -3338 442894
rect -3894 442338 -3658 442574
rect -3574 442338 -3338 442574
rect -3894 406658 -3658 406894
rect -3574 406658 -3338 406894
rect -3894 406338 -3658 406574
rect -3574 406338 -3338 406574
rect -3894 370658 -3658 370894
rect -3574 370658 -3338 370894
rect -3894 370338 -3658 370574
rect -3574 370338 -3338 370574
rect -3894 334658 -3658 334894
rect -3574 334658 -3338 334894
rect -3894 334338 -3658 334574
rect -3574 334338 -3338 334574
rect -3894 298658 -3658 298894
rect -3574 298658 -3338 298894
rect -3894 298338 -3658 298574
rect -3574 298338 -3338 298574
rect -3894 262658 -3658 262894
rect -3574 262658 -3338 262894
rect -3894 262338 -3658 262574
rect -3574 262338 -3338 262574
rect -3894 226658 -3658 226894
rect -3574 226658 -3338 226894
rect -3894 226338 -3658 226574
rect -3574 226338 -3338 226574
rect -3894 190658 -3658 190894
rect -3574 190658 -3338 190894
rect -3894 190338 -3658 190574
rect -3574 190338 -3338 190574
rect -3894 154658 -3658 154894
rect -3574 154658 -3338 154894
rect -3894 154338 -3658 154574
rect -3574 154338 -3338 154574
rect -3894 118658 -3658 118894
rect -3574 118658 -3338 118894
rect -3894 118338 -3658 118574
rect -3574 118338 -3338 118574
rect -3894 82658 -3658 82894
rect -3574 82658 -3338 82894
rect -3894 82338 -3658 82574
rect -3574 82338 -3338 82574
rect -3894 46658 -3658 46894
rect -3574 46658 -3338 46894
rect -3894 46338 -3658 46574
rect -3574 46338 -3338 46574
rect -3894 10658 -3658 10894
rect -3574 10658 -3338 10894
rect -3894 10338 -3658 10574
rect -3574 10338 -3338 10574
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 690938 -2698 691174
rect -2614 690938 -2378 691174
rect -2934 690618 -2698 690854
rect -2614 690618 -2378 690854
rect -2934 654938 -2698 655174
rect -2614 654938 -2378 655174
rect -2934 654618 -2698 654854
rect -2614 654618 -2378 654854
rect -2934 618938 -2698 619174
rect -2614 618938 -2378 619174
rect -2934 618618 -2698 618854
rect -2614 618618 -2378 618854
rect -2934 582938 -2698 583174
rect -2614 582938 -2378 583174
rect -2934 582618 -2698 582854
rect -2614 582618 -2378 582854
rect -2934 546938 -2698 547174
rect -2614 546938 -2378 547174
rect -2934 546618 -2698 546854
rect -2614 546618 -2378 546854
rect -2934 510938 -2698 511174
rect -2614 510938 -2378 511174
rect -2934 510618 -2698 510854
rect -2614 510618 -2378 510854
rect -2934 474938 -2698 475174
rect -2614 474938 -2378 475174
rect -2934 474618 -2698 474854
rect -2614 474618 -2378 474854
rect -2934 438938 -2698 439174
rect -2614 438938 -2378 439174
rect -2934 438618 -2698 438854
rect -2614 438618 -2378 438854
rect -2934 402938 -2698 403174
rect -2614 402938 -2378 403174
rect -2934 402618 -2698 402854
rect -2614 402618 -2378 402854
rect -2934 366938 -2698 367174
rect -2614 366938 -2378 367174
rect -2934 366618 -2698 366854
rect -2614 366618 -2378 366854
rect -2934 330938 -2698 331174
rect -2614 330938 -2378 331174
rect -2934 330618 -2698 330854
rect -2614 330618 -2378 330854
rect -2934 294938 -2698 295174
rect -2614 294938 -2378 295174
rect -2934 294618 -2698 294854
rect -2614 294618 -2378 294854
rect -2934 258938 -2698 259174
rect -2614 258938 -2378 259174
rect -2934 258618 -2698 258854
rect -2614 258618 -2378 258854
rect -2934 222938 -2698 223174
rect -2614 222938 -2378 223174
rect -2934 222618 -2698 222854
rect -2614 222618 -2378 222854
rect -2934 186938 -2698 187174
rect -2614 186938 -2378 187174
rect -2934 186618 -2698 186854
rect -2614 186618 -2378 186854
rect -2934 150938 -2698 151174
rect -2614 150938 -2378 151174
rect -2934 150618 -2698 150854
rect -2614 150618 -2378 150854
rect -2934 114938 -2698 115174
rect -2614 114938 -2378 115174
rect -2934 114618 -2698 114854
rect -2614 114618 -2378 114854
rect -2934 78938 -2698 79174
rect -2614 78938 -2378 79174
rect -2934 78618 -2698 78854
rect -2614 78618 -2378 78854
rect -2934 42938 -2698 43174
rect -2614 42938 -2378 43174
rect -2934 42618 -2698 42854
rect -2614 42618 -2378 42854
rect -2934 6938 -2698 7174
rect -2614 6938 -2378 7174
rect -2934 6618 -2698 6854
rect -2614 6618 -2378 6854
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 5546 705562 5782 705798
rect 5866 705562 6102 705798
rect 5546 705242 5782 705478
rect 5866 705242 6102 705478
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 5546 -1542 5782 -1306
rect 5866 -1542 6102 -1306
rect 5546 -1862 5782 -1626
rect 5866 -1862 6102 -1626
rect 9266 706522 9502 706758
rect 9586 706522 9822 706758
rect 9266 706202 9502 706438
rect 9586 706202 9822 706438
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 9266 -2502 9502 -2266
rect 9586 -2502 9822 -2266
rect 9266 -2822 9502 -2586
rect 9586 -2822 9822 -2586
rect 12986 707482 13222 707718
rect 13306 707482 13542 707718
rect 12986 707162 13222 707398
rect 13306 707162 13542 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 16706 708442 16942 708678
rect 17026 708442 17262 708678
rect 16706 708122 16942 708358
rect 17026 708122 17262 708358
rect 16706 666098 16942 666334
rect 17026 666098 17262 666334
rect 16706 665778 16942 666014
rect 17026 665778 17262 666014
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 16706 630098 16942 630334
rect 17026 630098 17262 630334
rect 16706 629778 16942 630014
rect 17026 629778 17262 630014
rect 16706 594098 16942 594334
rect 17026 594098 17262 594334
rect 16706 593778 16942 594014
rect 17026 593778 17262 594014
rect 16706 558098 16942 558334
rect 17026 558098 17262 558334
rect 16706 557778 16942 558014
rect 17026 557778 17262 558014
rect 20426 709402 20662 709638
rect 20746 709402 20982 709638
rect 20426 709082 20662 709318
rect 20746 709082 20982 709318
rect 20426 669818 20662 670054
rect 20746 669818 20982 670054
rect 20426 669498 20662 669734
rect 20746 669498 20982 669734
rect 20426 633818 20662 634054
rect 20746 633818 20982 634054
rect 20426 633498 20662 633734
rect 20746 633498 20982 633734
rect 20426 597818 20662 598054
rect 20746 597818 20982 598054
rect 20426 597498 20662 597734
rect 20746 597498 20982 597734
rect 20426 561818 20662 562054
rect 20746 561818 20982 562054
rect 20426 561498 20662 561734
rect 20746 561498 20982 561734
rect 16706 522098 16942 522334
rect 17026 522098 17262 522334
rect 16706 521778 16942 522014
rect 17026 521778 17262 522014
rect 16706 486098 16942 486334
rect 17026 486098 17262 486334
rect 16706 485778 16942 486014
rect 17026 485778 17262 486014
rect 16706 450098 16942 450334
rect 17026 450098 17262 450334
rect 16706 449778 16942 450014
rect 17026 449778 17262 450014
rect 16706 414098 16942 414334
rect 17026 414098 17262 414334
rect 16706 413778 16942 414014
rect 17026 413778 17262 414014
rect 16706 378098 16942 378334
rect 17026 378098 17262 378334
rect 16706 377778 16942 378014
rect 17026 377778 17262 378014
rect 16706 342098 16942 342334
rect 17026 342098 17262 342334
rect 16706 341778 16942 342014
rect 17026 341778 17262 342014
rect 16706 306098 16942 306334
rect 17026 306098 17262 306334
rect 16706 305778 16942 306014
rect 17026 305778 17262 306014
rect 16706 270098 16942 270334
rect 17026 270098 17262 270334
rect 16706 269778 16942 270014
rect 17026 269778 17262 270014
rect 16706 234098 16942 234334
rect 17026 234098 17262 234334
rect 16706 233778 16942 234014
rect 17026 233778 17262 234014
rect 16706 198098 16942 198334
rect 17026 198098 17262 198334
rect 16706 197778 16942 198014
rect 17026 197778 17262 198014
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 12986 -3462 13222 -3226
rect 13306 -3462 13542 -3226
rect 12986 -3782 13222 -3546
rect 13306 -3782 13542 -3546
rect 20426 525818 20662 526054
rect 20746 525818 20982 526054
rect 20426 525498 20662 525734
rect 20746 525498 20982 525734
rect 24146 710362 24382 710598
rect 24466 710362 24702 710598
rect 24146 710042 24382 710278
rect 24466 710042 24702 710278
rect 24146 673538 24382 673774
rect 24466 673538 24702 673774
rect 24146 673218 24382 673454
rect 24466 673218 24702 673454
rect 24146 637538 24382 637774
rect 24466 637538 24702 637774
rect 24146 637218 24382 637454
rect 24466 637218 24702 637454
rect 27866 711322 28102 711558
rect 28186 711322 28422 711558
rect 27866 711002 28102 711238
rect 28186 711002 28422 711238
rect 27866 677258 28102 677494
rect 28186 677258 28422 677494
rect 27866 676938 28102 677174
rect 28186 676938 28422 677174
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 27866 641258 28102 641494
rect 28186 641258 28422 641494
rect 27866 640938 28102 641174
rect 28186 640938 28422 641174
rect 24146 601538 24382 601774
rect 24466 601538 24702 601774
rect 24146 601218 24382 601454
rect 24466 601218 24702 601454
rect 24146 565538 24382 565774
rect 24466 565538 24702 565774
rect 24146 565218 24382 565454
rect 24466 565218 24702 565454
rect 24146 529538 24382 529774
rect 24466 529538 24702 529774
rect 24146 529218 24382 529454
rect 24466 529218 24702 529454
rect 20426 489818 20662 490054
rect 20746 489818 20982 490054
rect 20426 489498 20662 489734
rect 20746 489498 20982 489734
rect 20426 453818 20662 454054
rect 20746 453818 20982 454054
rect 20426 453498 20662 453734
rect 20746 453498 20982 453734
rect 20426 417818 20662 418054
rect 20746 417818 20982 418054
rect 20426 417498 20662 417734
rect 20746 417498 20982 417734
rect 20426 381818 20662 382054
rect 20746 381818 20982 382054
rect 20426 381498 20662 381734
rect 20746 381498 20982 381734
rect 20426 345818 20662 346054
rect 20746 345818 20982 346054
rect 20426 345498 20662 345734
rect 20746 345498 20982 345734
rect 20426 309818 20662 310054
rect 20746 309818 20982 310054
rect 20426 309498 20662 309734
rect 20746 309498 20982 309734
rect 20426 273818 20662 274054
rect 20746 273818 20982 274054
rect 20426 273498 20662 273734
rect 20746 273498 20982 273734
rect 20426 237818 20662 238054
rect 20746 237818 20982 238054
rect 20426 237498 20662 237734
rect 20746 237498 20982 237734
rect 20426 201818 20662 202054
rect 20746 201818 20982 202054
rect 20426 201498 20662 201734
rect 20746 201498 20982 201734
rect 16706 162098 16942 162334
rect 17026 162098 17262 162334
rect 16706 161778 16942 162014
rect 17026 161778 17262 162014
rect 16706 126098 16942 126334
rect 17026 126098 17262 126334
rect 16706 125778 16942 126014
rect 17026 125778 17262 126014
rect 16706 90098 16942 90334
rect 17026 90098 17262 90334
rect 16706 89778 16942 90014
rect 17026 89778 17262 90014
rect 16706 54098 16942 54334
rect 17026 54098 17262 54334
rect 16706 53778 16942 54014
rect 17026 53778 17262 54014
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 16706 -4422 16942 -4186
rect 17026 -4422 17262 -4186
rect 16706 -4742 16942 -4506
rect 17026 -4742 17262 -4506
rect 24146 493538 24382 493774
rect 24466 493538 24702 493774
rect 24146 493218 24382 493454
rect 24466 493218 24702 493454
rect 24146 457538 24382 457774
rect 24466 457538 24702 457774
rect 24146 457218 24382 457454
rect 24466 457218 24702 457454
rect 24146 421538 24382 421774
rect 24466 421538 24702 421774
rect 24146 421218 24382 421454
rect 24466 421218 24702 421454
rect 24146 385538 24382 385774
rect 24466 385538 24702 385774
rect 24146 385218 24382 385454
rect 24466 385218 24702 385454
rect 24146 349538 24382 349774
rect 24466 349538 24702 349774
rect 24146 349218 24382 349454
rect 24466 349218 24702 349454
rect 24146 313538 24382 313774
rect 24466 313538 24702 313774
rect 24146 313218 24382 313454
rect 24466 313218 24702 313454
rect 24146 277538 24382 277774
rect 24466 277538 24702 277774
rect 24146 277218 24382 277454
rect 24466 277218 24702 277454
rect 24146 241538 24382 241774
rect 24466 241538 24702 241774
rect 24146 241218 24382 241454
rect 24466 241218 24702 241454
rect 24146 205538 24382 205774
rect 24466 205538 24702 205774
rect 24146 205218 24382 205454
rect 24466 205218 24702 205454
rect 20426 165818 20662 166054
rect 20746 165818 20982 166054
rect 20426 165498 20662 165734
rect 20746 165498 20982 165734
rect 20426 129818 20662 130054
rect 20746 129818 20982 130054
rect 20426 129498 20662 129734
rect 20746 129498 20982 129734
rect 20426 93818 20662 94054
rect 20746 93818 20982 94054
rect 20426 93498 20662 93734
rect 20746 93498 20982 93734
rect 20426 57818 20662 58054
rect 20746 57818 20982 58054
rect 20426 57498 20662 57734
rect 20746 57498 20982 57734
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 20426 -5382 20662 -5146
rect 20746 -5382 20982 -5146
rect 20426 -5702 20662 -5466
rect 20746 -5702 20982 -5466
rect 27866 605258 28102 605494
rect 28186 605258 28422 605494
rect 27866 604938 28102 605174
rect 28186 604938 28422 605174
rect 27866 569258 28102 569494
rect 28186 569258 28422 569494
rect 27866 568938 28102 569174
rect 28186 568938 28422 569174
rect 27866 533258 28102 533494
rect 28186 533258 28422 533494
rect 27866 532938 28102 533174
rect 28186 532938 28422 533174
rect 27866 497258 28102 497494
rect 28186 497258 28422 497494
rect 27866 496938 28102 497174
rect 28186 496938 28422 497174
rect 27866 461258 28102 461494
rect 28186 461258 28422 461494
rect 27866 460938 28102 461174
rect 28186 460938 28422 461174
rect 27866 425258 28102 425494
rect 28186 425258 28422 425494
rect 27866 424938 28102 425174
rect 28186 424938 28422 425174
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 27866 389258 28102 389494
rect 28186 389258 28422 389494
rect 27866 388938 28102 389174
rect 28186 388938 28422 389174
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 41546 705562 41782 705798
rect 41866 705562 42102 705798
rect 41546 705242 41782 705478
rect 41866 705242 42102 705478
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 45266 706522 45502 706758
rect 45586 706522 45822 706758
rect 45266 706202 45502 706438
rect 45586 706202 45822 706438
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 27866 353258 28102 353494
rect 28186 353258 28422 353494
rect 27866 352938 28102 353174
rect 28186 352938 28422 353174
rect 27866 317258 28102 317494
rect 28186 317258 28422 317494
rect 27866 316938 28102 317174
rect 28186 316938 28422 317174
rect 27866 281258 28102 281494
rect 28186 281258 28422 281494
rect 27866 280938 28102 281174
rect 28186 280938 28422 281174
rect 27866 245258 28102 245494
rect 28186 245258 28422 245494
rect 27866 244938 28102 245174
rect 28186 244938 28422 245174
rect 27866 209258 28102 209494
rect 28186 209258 28422 209494
rect 27866 208938 28102 209174
rect 28186 208938 28422 209174
rect 24146 169538 24382 169774
rect 24466 169538 24702 169774
rect 24146 169218 24382 169454
rect 24466 169218 24702 169454
rect 24146 133538 24382 133774
rect 24466 133538 24702 133774
rect 24146 133218 24382 133454
rect 24466 133218 24702 133454
rect 24146 97538 24382 97774
rect 24466 97538 24702 97774
rect 24146 97218 24382 97454
rect 24466 97218 24702 97454
rect 24146 61538 24382 61774
rect 24466 61538 24702 61774
rect 24146 61218 24382 61454
rect 24466 61218 24702 61454
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 24146 -6342 24382 -6106
rect 24466 -6342 24702 -6106
rect 24146 -6662 24382 -6426
rect 24466 -6662 24702 -6426
rect 27866 173258 28102 173494
rect 28186 173258 28422 173494
rect 27866 172938 28102 173174
rect 28186 172938 28422 173174
rect 27866 137258 28102 137494
rect 28186 137258 28422 137494
rect 27866 136938 28102 137174
rect 28186 136938 28422 137174
rect 27866 101258 28102 101494
rect 28186 101258 28422 101494
rect 27866 100938 28102 101174
rect 28186 100938 28422 101174
rect 27866 65258 28102 65494
rect 28186 65258 28422 65494
rect 27866 64938 28102 65174
rect 28186 64938 28422 65174
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 27866 -7302 28102 -7066
rect 28186 -7302 28422 -7066
rect 27866 -7622 28102 -7386
rect 28186 -7622 28422 -7386
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 48986 707482 49222 707718
rect 49306 707482 49542 707718
rect 48986 707162 49222 707398
rect 49306 707162 49542 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 52706 708442 52942 708678
rect 53026 708442 53262 708678
rect 52706 708122 52942 708358
rect 53026 708122 53262 708358
rect 52706 666098 52942 666334
rect 53026 666098 53262 666334
rect 52706 665778 52942 666014
rect 53026 665778 53262 666014
rect 56426 709402 56662 709638
rect 56746 709402 56982 709638
rect 56426 709082 56662 709318
rect 56746 709082 56982 709318
rect 56426 669818 56662 670054
rect 56746 669818 56982 670054
rect 56426 669498 56662 669734
rect 56746 669498 56982 669734
rect 52706 630098 52942 630334
rect 53026 630098 53262 630334
rect 52706 629778 52942 630014
rect 53026 629778 53262 630014
rect 52706 594098 52942 594334
rect 53026 594098 53262 594334
rect 52706 593778 52942 594014
rect 53026 593778 53262 594014
rect 52706 558098 52942 558334
rect 53026 558098 53262 558334
rect 52706 557778 52942 558014
rect 53026 557778 53262 558014
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -1542 41782 -1306
rect 41866 -1542 42102 -1306
rect 41546 -1862 41782 -1626
rect 41866 -1862 42102 -1626
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 52706 522098 52942 522334
rect 53026 522098 53262 522334
rect 52706 521778 52942 522014
rect 53026 521778 53262 522014
rect 52706 486098 52942 486334
rect 53026 486098 53262 486334
rect 52706 485778 52942 486014
rect 53026 485778 53262 486014
rect 52706 450098 52942 450334
rect 53026 450098 53262 450334
rect 52706 449778 52942 450014
rect 53026 449778 53262 450014
rect 52706 414098 52942 414334
rect 53026 414098 53262 414334
rect 52706 413778 52942 414014
rect 53026 413778 53262 414014
rect 52706 378098 52942 378334
rect 53026 378098 53262 378334
rect 52706 377778 52942 378014
rect 53026 377778 53262 378014
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -2502 45502 -2266
rect 45586 -2502 45822 -2266
rect 45266 -2822 45502 -2586
rect 45586 -2822 45822 -2586
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 48986 -3462 49222 -3226
rect 49306 -3462 49542 -3226
rect 48986 -3782 49222 -3546
rect 49306 -3782 49542 -3546
rect 52706 342098 52942 342334
rect 53026 342098 53262 342334
rect 52706 341778 52942 342014
rect 53026 341778 53262 342014
rect 52706 306098 52942 306334
rect 53026 306098 53262 306334
rect 52706 305778 52942 306014
rect 53026 305778 53262 306014
rect 56426 633818 56662 634054
rect 56746 633818 56982 634054
rect 56426 633498 56662 633734
rect 56746 633498 56982 633734
rect 60146 710362 60382 710598
rect 60466 710362 60702 710598
rect 60146 710042 60382 710278
rect 60466 710042 60702 710278
rect 60146 673538 60382 673774
rect 60466 673538 60702 673774
rect 60146 673218 60382 673454
rect 60466 673218 60702 673454
rect 60146 637538 60382 637774
rect 60466 637538 60702 637774
rect 60146 637218 60382 637454
rect 60466 637218 60702 637454
rect 63866 711322 64102 711558
rect 64186 711322 64422 711558
rect 63866 711002 64102 711238
rect 64186 711002 64422 711238
rect 63866 677258 64102 677494
rect 64186 677258 64422 677494
rect 63866 676938 64102 677174
rect 64186 676938 64422 677174
rect 63866 641258 64102 641494
rect 64186 641258 64422 641494
rect 63866 640938 64102 641174
rect 64186 640938 64422 641174
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 705562 77782 705798
rect 77866 705562 78102 705798
rect 77546 705242 77782 705478
rect 77866 705242 78102 705478
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 706522 81502 706758
rect 81586 706522 81822 706758
rect 81266 706202 81502 706438
rect 81586 706202 81822 706438
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 84986 707482 85222 707718
rect 85306 707482 85542 707718
rect 84986 707162 85222 707398
rect 85306 707162 85542 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 88706 708442 88942 708678
rect 89026 708442 89262 708678
rect 88706 708122 88942 708358
rect 89026 708122 89262 708358
rect 88706 666098 88942 666334
rect 89026 666098 89262 666334
rect 88706 665778 88942 666014
rect 89026 665778 89262 666014
rect 92426 709402 92662 709638
rect 92746 709402 92982 709638
rect 92426 709082 92662 709318
rect 92746 709082 92982 709318
rect 92426 669818 92662 670054
rect 92746 669818 92982 670054
rect 92426 669498 92662 669734
rect 92746 669498 92982 669734
rect 92426 633818 92662 634054
rect 92746 633818 92982 634054
rect 92426 633498 92662 633734
rect 92746 633498 92982 633734
rect 96146 710362 96382 710598
rect 96466 710362 96702 710598
rect 96146 710042 96382 710278
rect 96466 710042 96702 710278
rect 96146 673538 96382 673774
rect 96466 673538 96702 673774
rect 96146 673218 96382 673454
rect 96466 673218 96702 673454
rect 96146 637538 96382 637774
rect 96466 637538 96702 637774
rect 96146 637218 96382 637454
rect 96466 637218 96702 637454
rect 99866 711322 100102 711558
rect 100186 711322 100422 711558
rect 99866 711002 100102 711238
rect 100186 711002 100422 711238
rect 99866 677258 100102 677494
rect 100186 677258 100422 677494
rect 99866 676938 100102 677174
rect 100186 676938 100422 677174
rect 99866 641258 100102 641494
rect 100186 641258 100422 641494
rect 99866 640938 100102 641174
rect 100186 640938 100422 641174
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 705562 113782 705798
rect 113866 705562 114102 705798
rect 113546 705242 113782 705478
rect 113866 705242 114102 705478
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 706522 117502 706758
rect 117586 706522 117822 706758
rect 117266 706202 117502 706438
rect 117586 706202 117822 706438
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 120986 707482 121222 707718
rect 121306 707482 121542 707718
rect 120986 707162 121222 707398
rect 121306 707162 121542 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 124706 708442 124942 708678
rect 125026 708442 125262 708678
rect 124706 708122 124942 708358
rect 125026 708122 125262 708358
rect 124706 666098 124942 666334
rect 125026 666098 125262 666334
rect 124706 665778 124942 666014
rect 125026 665778 125262 666014
rect 128426 709402 128662 709638
rect 128746 709402 128982 709638
rect 128426 709082 128662 709318
rect 128746 709082 128982 709318
rect 128426 669818 128662 670054
rect 128746 669818 128982 670054
rect 128426 669498 128662 669734
rect 128746 669498 128982 669734
rect 128426 633818 128662 634054
rect 128746 633818 128982 634054
rect 128426 633498 128662 633734
rect 128746 633498 128982 633734
rect 132146 710362 132382 710598
rect 132466 710362 132702 710598
rect 132146 710042 132382 710278
rect 132466 710042 132702 710278
rect 132146 673538 132382 673774
rect 132466 673538 132702 673774
rect 132146 673218 132382 673454
rect 132466 673218 132702 673454
rect 132146 637538 132382 637774
rect 132466 637538 132702 637774
rect 132146 637218 132382 637454
rect 132466 637218 132702 637454
rect 135866 711322 136102 711558
rect 136186 711322 136422 711558
rect 135866 711002 136102 711238
rect 136186 711002 136422 711238
rect 135866 677258 136102 677494
rect 136186 677258 136422 677494
rect 135866 676938 136102 677174
rect 136186 676938 136422 677174
rect 135866 641258 136102 641494
rect 136186 641258 136422 641494
rect 135866 640938 136102 641174
rect 136186 640938 136422 641174
rect 56426 597818 56662 598054
rect 56746 597818 56982 598054
rect 56426 597498 56662 597734
rect 56746 597498 56982 597734
rect 56426 561818 56662 562054
rect 56746 561818 56982 562054
rect 56426 561498 56662 561734
rect 56746 561498 56982 561734
rect 56426 525818 56662 526054
rect 56746 525818 56982 526054
rect 56426 525498 56662 525734
rect 56746 525498 56982 525734
rect 56426 489818 56662 490054
rect 56746 489818 56982 490054
rect 56426 489498 56662 489734
rect 56746 489498 56982 489734
rect 56426 453818 56662 454054
rect 56746 453818 56982 454054
rect 56426 453498 56662 453734
rect 56746 453498 56982 453734
rect 79610 618938 79846 619174
rect 79610 618618 79846 618854
rect 110330 618938 110566 619174
rect 110330 618618 110566 618854
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 125690 615218 125926 615454
rect 125690 614898 125926 615134
rect 135866 605258 136102 605494
rect 136186 605258 136422 605494
rect 135866 604938 136102 605174
rect 136186 604938 136422 605174
rect 79610 582938 79846 583174
rect 79610 582618 79846 582854
rect 110330 582938 110566 583174
rect 110330 582618 110566 582854
rect 64250 579218 64486 579454
rect 64250 578898 64486 579134
rect 94970 579218 95206 579454
rect 94970 578898 95206 579134
rect 125690 579218 125926 579454
rect 125690 578898 125926 579134
rect 135866 569258 136102 569494
rect 136186 569258 136422 569494
rect 135866 568938 136102 569174
rect 136186 568938 136422 569174
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 60146 529538 60382 529774
rect 60466 529538 60702 529774
rect 60146 529218 60382 529454
rect 60466 529218 60702 529454
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 60146 493538 60382 493774
rect 60466 493538 60702 493774
rect 60146 493218 60382 493454
rect 60466 493218 60702 493454
rect 64250 471218 64486 471454
rect 64250 470898 64486 471134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 60146 457538 60382 457774
rect 60466 457538 60702 457774
rect 60146 457218 60382 457454
rect 60466 457218 60702 457454
rect 56426 417818 56662 418054
rect 56746 417818 56982 418054
rect 56426 417498 56662 417734
rect 56746 417498 56982 417734
rect 56426 381818 56662 382054
rect 56746 381818 56982 382054
rect 56426 381498 56662 381734
rect 56746 381498 56982 381734
rect 56426 345818 56662 346054
rect 56746 345818 56982 346054
rect 56426 345498 56662 345734
rect 56746 345498 56982 345734
rect 56426 309818 56662 310054
rect 56746 309818 56982 310054
rect 56426 309498 56662 309734
rect 56746 309498 56982 309734
rect 54250 291218 54486 291454
rect 54250 290898 54486 291134
rect 52706 270098 52942 270334
rect 53026 270098 53262 270334
rect 52706 269778 52942 270014
rect 53026 269778 53262 270014
rect 64250 435218 64486 435454
rect 64250 434898 64486 435134
rect 73826 435218 74062 435454
rect 74146 435218 74382 435454
rect 73826 434898 74062 435134
rect 74146 434898 74382 435134
rect 60146 421538 60382 421774
rect 60466 421538 60702 421774
rect 60146 421218 60382 421454
rect 60466 421218 60702 421454
rect 64250 399218 64486 399454
rect 64250 398898 64486 399134
rect 73826 399218 74062 399454
rect 74146 399218 74382 399454
rect 73826 398898 74062 399134
rect 74146 398898 74382 399134
rect 60146 385538 60382 385774
rect 60466 385538 60702 385774
rect 60146 385218 60382 385454
rect 60466 385218 60702 385454
rect 60146 349538 60382 349774
rect 60466 349538 60702 349774
rect 60146 349218 60382 349454
rect 60466 349218 60702 349454
rect 60146 313538 60382 313774
rect 60466 313538 60702 313774
rect 60146 313218 60382 313454
rect 60466 313218 60702 313454
rect 63866 389258 64102 389494
rect 64186 389258 64422 389494
rect 63866 388938 64102 389174
rect 64186 388938 64422 389174
rect 63866 353258 64102 353494
rect 64186 353258 64422 353494
rect 63866 352938 64102 353174
rect 64186 352938 64422 353174
rect 63866 317258 64102 317494
rect 64186 317258 64422 317494
rect 63866 316938 64102 317174
rect 64186 316938 64422 317174
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 79610 510938 79846 511174
rect 79610 510618 79846 510854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 79610 474938 79846 475174
rect 79610 474618 79846 474854
rect 81266 442658 81502 442894
rect 81586 442658 81822 442894
rect 81266 442338 81502 442574
rect 81586 442338 81822 442574
rect 77546 438938 77782 439174
rect 77866 438938 78102 439174
rect 77546 438618 77782 438854
rect 77866 438618 78102 438854
rect 79610 438938 79846 439174
rect 79610 438618 79846 438854
rect 81266 406658 81502 406894
rect 81586 406658 81822 406894
rect 81266 406338 81502 406574
rect 81586 406338 81822 406574
rect 77546 402938 77782 403174
rect 77866 402938 78102 403174
rect 77546 402618 77782 402854
rect 77866 402618 78102 402854
rect 79610 402938 79846 403174
rect 79610 402618 79846 402854
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 84986 446378 85222 446614
rect 85306 446378 85542 446614
rect 84986 446058 85222 446294
rect 85306 446058 85542 446294
rect 84986 410378 85222 410614
rect 85306 410378 85542 410614
rect 84986 410058 85222 410294
rect 85306 410058 85542 410294
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 88706 558098 88942 558334
rect 89026 558098 89262 558334
rect 88706 557778 88942 558014
rect 89026 557778 89262 558014
rect 88706 522098 88942 522334
rect 89026 522098 89262 522334
rect 88706 521778 88942 522014
rect 89026 521778 89262 522014
rect 88706 486098 88942 486334
rect 89026 486098 89262 486334
rect 88706 485778 88942 486014
rect 89026 485778 89262 486014
rect 88706 450098 88942 450334
rect 89026 450098 89262 450334
rect 88706 449778 88942 450014
rect 89026 449778 89262 450014
rect 88706 414098 88942 414334
rect 89026 414098 89262 414334
rect 88706 413778 88942 414014
rect 89026 413778 89262 414014
rect 88706 378098 88942 378334
rect 89026 378098 89262 378334
rect 88706 377778 88942 378014
rect 89026 377778 89262 378014
rect 88706 342098 88942 342334
rect 89026 342098 89262 342334
rect 88706 341778 88942 342014
rect 89026 341778 89262 342014
rect 88706 306098 88942 306334
rect 89026 306098 89262 306334
rect 88706 305778 88942 306014
rect 89026 305778 89262 306014
rect 92426 525818 92662 526054
rect 92746 525818 92982 526054
rect 92426 525498 92662 525734
rect 92746 525498 92982 525734
rect 96146 529538 96382 529774
rect 96466 529538 96702 529774
rect 96146 529218 96382 529454
rect 96466 529218 96702 529454
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 92426 489818 92662 490054
rect 92746 489818 92982 490054
rect 92426 489498 92662 489734
rect 92746 489498 92982 489734
rect 96146 493538 96382 493774
rect 96466 493538 96702 493774
rect 96146 493218 96382 493454
rect 96466 493218 96702 493454
rect 94970 471218 95206 471454
rect 94970 470898 95206 471134
rect 92426 453818 92662 454054
rect 92746 453818 92982 454054
rect 92426 453498 92662 453734
rect 92746 453498 92982 453734
rect 96146 457538 96382 457774
rect 96466 457538 96702 457774
rect 96146 457218 96382 457454
rect 96466 457218 96702 457454
rect 94970 435218 95206 435454
rect 94970 434898 95206 435134
rect 92426 417818 92662 418054
rect 92746 417818 92982 418054
rect 92426 417498 92662 417734
rect 92746 417498 92982 417734
rect 96146 421538 96382 421774
rect 96466 421538 96702 421774
rect 96146 421218 96382 421454
rect 96466 421218 96702 421454
rect 94970 399218 95206 399454
rect 94970 398898 95206 399134
rect 92426 381818 92662 382054
rect 92746 381818 92982 382054
rect 92426 381498 92662 381734
rect 92746 381498 92982 381734
rect 92426 345818 92662 346054
rect 92746 345818 92982 346054
rect 92426 345498 92662 345734
rect 92746 345498 92982 345734
rect 92426 309818 92662 310054
rect 92746 309818 92982 310054
rect 92426 309498 92662 309734
rect 92746 309498 92982 309734
rect 96146 385538 96382 385774
rect 96466 385538 96702 385774
rect 96146 385218 96382 385454
rect 96466 385218 96702 385454
rect 96146 349538 96382 349774
rect 96466 349538 96702 349774
rect 96146 349218 96382 349454
rect 96466 349218 96702 349454
rect 96146 313538 96382 313774
rect 96466 313538 96702 313774
rect 96146 313218 96382 313454
rect 96466 313218 96702 313454
rect 99866 533258 100102 533494
rect 100186 533258 100422 533494
rect 99866 532938 100102 533174
rect 100186 532938 100422 533174
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 110330 510938 110566 511174
rect 110330 510618 110566 510854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 99866 497258 100102 497494
rect 100186 497258 100422 497494
rect 99866 496938 100102 497174
rect 100186 496938 100422 497174
rect 110330 474938 110566 475174
rect 110330 474618 110566 474854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 99866 461258 100102 461494
rect 100186 461258 100422 461494
rect 99866 460938 100102 461174
rect 100186 460938 100422 461174
rect 110330 438938 110566 439174
rect 110330 438618 110566 438854
rect 113546 438938 113782 439174
rect 113866 438938 114102 439174
rect 113546 438618 113782 438854
rect 113866 438618 114102 438854
rect 99866 425258 100102 425494
rect 100186 425258 100422 425494
rect 99866 424938 100102 425174
rect 100186 424938 100422 425174
rect 110330 402938 110566 403174
rect 110330 402618 110566 402854
rect 113546 402938 113782 403174
rect 113866 402938 114102 403174
rect 113546 402618 113782 402854
rect 113866 402618 114102 402854
rect 99866 389258 100102 389494
rect 100186 389258 100422 389494
rect 99866 388938 100102 389174
rect 100186 388938 100422 389174
rect 99866 353258 100102 353494
rect 100186 353258 100422 353494
rect 99866 352938 100102 353174
rect 100186 352938 100422 353174
rect 99866 317258 100102 317494
rect 100186 317258 100422 317494
rect 99866 316938 100102 317174
rect 100186 316938 100422 317174
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 69610 294938 69846 295174
rect 69610 294618 69846 294854
rect 100330 294938 100566 295174
rect 100330 294618 100566 294854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 84970 291218 85206 291454
rect 84970 290898 85206 291134
rect 56426 273818 56662 274054
rect 56746 273818 56982 274054
rect 56426 273498 56662 273734
rect 56746 273498 56982 273734
rect 54250 255218 54486 255454
rect 54250 254898 54486 255134
rect 52706 234098 52942 234334
rect 53026 234098 53262 234334
rect 52706 233778 52942 234014
rect 53026 233778 53262 234014
rect 52706 198098 52942 198334
rect 53026 198098 53262 198334
rect 52706 197778 52942 198014
rect 53026 197778 53262 198014
rect 52706 162098 52942 162334
rect 53026 162098 53262 162334
rect 52706 161778 52942 162014
rect 53026 161778 53262 162014
rect 69610 258938 69846 259174
rect 69610 258618 69846 258854
rect 100330 258938 100566 259174
rect 100330 258618 100566 258854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 84970 255218 85206 255454
rect 84970 254898 85206 255134
rect 56426 237818 56662 238054
rect 56746 237818 56982 238054
rect 56426 237498 56662 237734
rect 56746 237498 56982 237734
rect 56426 201818 56662 202054
rect 56746 201818 56982 202054
rect 56426 201498 56662 201734
rect 56746 201498 56982 201734
rect 56426 165818 56662 166054
rect 56746 165818 56982 166054
rect 56426 165498 56662 165734
rect 56746 165498 56982 165734
rect 52706 126098 52942 126334
rect 53026 126098 53262 126334
rect 52706 125778 52942 126014
rect 53026 125778 53262 126014
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 88706 234098 88942 234334
rect 89026 234098 89262 234334
rect 88706 233778 88942 234014
rect 89026 233778 89262 234014
rect 88706 198098 88942 198334
rect 89026 198098 89262 198334
rect 88706 197778 88942 198014
rect 89026 197778 89262 198014
rect 92426 237818 92662 238054
rect 92746 237818 92982 238054
rect 92426 237498 92662 237734
rect 92746 237498 92982 237734
rect 92426 201818 92662 202054
rect 92746 201818 92982 202054
rect 92426 201498 92662 201734
rect 92746 201498 92982 201734
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 442658 117502 442894
rect 117586 442658 117822 442894
rect 117266 442338 117502 442574
rect 117586 442338 117822 442574
rect 117266 406658 117502 406894
rect 117586 406658 117822 406894
rect 117266 406338 117502 406574
rect 117586 406338 117822 406574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 79610 150938 79846 151174
rect 79610 150618 79846 150854
rect 110330 150938 110566 151174
rect 110330 150618 110566 150854
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 56426 129818 56662 130054
rect 56746 129818 56982 130054
rect 56426 129498 56662 129734
rect 56746 129498 56982 129734
rect 52706 90098 52942 90334
rect 53026 90098 53262 90334
rect 52706 89778 52942 90014
rect 53026 89778 53262 90014
rect 56426 93818 56662 94054
rect 56746 93818 56982 94054
rect 56426 93498 56662 93734
rect 56746 93498 56982 93734
rect 55080 75218 55316 75454
rect 55080 74898 55316 75134
rect 52706 54098 52942 54334
rect 53026 54098 53262 54334
rect 52706 53778 52942 54014
rect 53026 53778 53262 54014
rect 52706 18098 52942 18334
rect 53026 18098 53262 18334
rect 52706 17778 52942 18014
rect 53026 17778 53262 18014
rect 52706 -4422 52942 -4186
rect 53026 -4422 53262 -4186
rect 52706 -4742 52942 -4506
rect 53026 -4742 53262 -4506
rect 56426 57818 56662 58054
rect 56746 57818 56982 58054
rect 56426 57498 56662 57734
rect 56746 57498 56982 57734
rect 60146 97538 60382 97774
rect 60466 97538 60702 97774
rect 60146 97218 60382 97454
rect 60466 97218 60702 97454
rect 59174 78938 59410 79174
rect 59174 78618 59410 78854
rect 63866 101258 64102 101494
rect 64186 101258 64422 101494
rect 63866 100938 64102 101174
rect 64186 100938 64422 101174
rect 63268 75218 63504 75454
rect 63268 74898 63504 75134
rect 60146 61538 60382 61774
rect 60466 61538 60702 61774
rect 60146 61218 60382 61454
rect 60466 61218 60702 61454
rect 56426 21818 56662 22054
rect 56746 21818 56982 22054
rect 56426 21498 56662 21734
rect 56746 21498 56982 21734
rect 56426 -5382 56662 -5146
rect 56746 -5382 56982 -5146
rect 56426 -5702 56662 -5466
rect 56746 -5702 56982 -5466
rect 60146 25538 60382 25774
rect 60466 25538 60702 25774
rect 60146 25218 60382 25454
rect 60466 25218 60702 25454
rect 60146 -6342 60382 -6106
rect 60466 -6342 60702 -6106
rect 60146 -6662 60382 -6426
rect 60466 -6662 60702 -6426
rect 73826 111218 74062 111454
rect 74146 111218 74382 111454
rect 73826 110898 74062 111134
rect 74146 110898 74382 111134
rect 67362 78938 67598 79174
rect 67362 78618 67598 78854
rect 71456 75218 71692 75454
rect 71456 74898 71692 75134
rect 77546 114938 77782 115174
rect 77866 114938 78102 115174
rect 77546 114618 77782 114854
rect 77866 114618 78102 114854
rect 75550 78938 75786 79174
rect 75550 78618 75786 78854
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 63866 65258 64102 65494
rect 64186 65258 64422 65494
rect 63866 64938 64102 65174
rect 64186 64938 64422 65174
rect 63866 29258 64102 29494
rect 64186 29258 64422 29494
rect 63866 28938 64102 29174
rect 64186 28938 64422 29174
rect 63866 -7302 64102 -7066
rect 64186 -7302 64422 -7066
rect 63866 -7622 64102 -7386
rect 64186 -7622 64422 -7386
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 81266 118658 81502 118894
rect 81586 118658 81822 118894
rect 81266 118338 81502 118574
rect 81586 118338 81822 118574
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 79644 75218 79880 75454
rect 79644 74898 79880 75134
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -1542 77782 -1306
rect 77866 -1542 78102 -1306
rect 77546 -1862 77782 -1626
rect 77866 -1862 78102 -1626
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 83738 78938 83974 79174
rect 83738 78618 83974 78854
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -2502 81502 -2266
rect 81586 -2502 81822 -2266
rect 81266 -2822 81502 -2586
rect 81586 -2822 81822 -2586
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 84986 -3462 85222 -3226
rect 85306 -3462 85542 -3226
rect 84986 -3782 85222 -3546
rect 85306 -3782 85542 -3546
rect 88706 90098 88942 90334
rect 89026 90098 89262 90334
rect 88706 89778 88942 90014
rect 89026 89778 89262 90014
rect 88706 54098 88942 54334
rect 89026 54098 89262 54334
rect 88706 53778 88942 54014
rect 89026 53778 89262 54014
rect 88706 18098 88942 18334
rect 89026 18098 89262 18334
rect 88706 17778 88942 18014
rect 89026 17778 89262 18014
rect 88706 -4422 88942 -4186
rect 89026 -4422 89262 -4186
rect 88706 -4742 88942 -4506
rect 89026 -4742 89262 -4506
rect 92426 93818 92662 94054
rect 92746 93818 92982 94054
rect 92426 93498 92662 93734
rect 92746 93498 92982 93734
rect 92426 57818 92662 58054
rect 92746 57818 92982 58054
rect 92426 57498 92662 57734
rect 92746 57498 92982 57734
rect 92426 21818 92662 22054
rect 92746 21818 92982 22054
rect 92426 21498 92662 21734
rect 92746 21498 92982 21734
rect 92426 -5382 92662 -5146
rect 92746 -5382 92982 -5146
rect 92426 -5702 92662 -5466
rect 92746 -5702 92982 -5466
rect 96146 97538 96382 97774
rect 96466 97538 96702 97774
rect 96146 97218 96382 97454
rect 96466 97218 96702 97454
rect 96146 61538 96382 61774
rect 96466 61538 96702 61774
rect 96146 61218 96382 61454
rect 96466 61218 96702 61454
rect 96146 25538 96382 25774
rect 96466 25538 96702 25774
rect 96146 25218 96382 25454
rect 96466 25218 96702 25454
rect 96146 -6342 96382 -6106
rect 96466 -6342 96702 -6106
rect 96146 -6662 96382 -6426
rect 96466 -6662 96702 -6426
rect 99866 101258 100102 101494
rect 100186 101258 100422 101494
rect 99866 100938 100102 101174
rect 100186 100938 100422 101174
rect 99866 65258 100102 65494
rect 100186 65258 100422 65494
rect 99866 64938 100102 65174
rect 100186 64938 100422 65174
rect 99866 29258 100102 29494
rect 100186 29258 100422 29494
rect 99866 28938 100102 29174
rect 100186 28938 100422 29174
rect 99866 -7302 100102 -7066
rect 100186 -7302 100422 -7066
rect 99866 -7622 100102 -7386
rect 100186 -7622 100422 -7386
rect 109826 111218 110062 111454
rect 110146 111218 110382 111454
rect 109826 110898 110062 111134
rect 110146 110898 110382 111134
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 114938 113782 115174
rect 113866 114938 114102 115174
rect 113546 114618 113782 114854
rect 113866 114618 114102 114854
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -1542 113782 -1306
rect 113866 -1542 114102 -1306
rect 113546 -1862 113782 -1626
rect 113866 -1862 114102 -1626
rect 117266 118658 117502 118894
rect 117586 118658 117822 118894
rect 117266 118338 117502 118574
rect 117586 118338 117822 118574
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -2502 117502 -2266
rect 117586 -2502 117822 -2266
rect 117266 -2822 117502 -2586
rect 117586 -2822 117822 -2586
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 120986 446378 121222 446614
rect 121306 446378 121542 446614
rect 120986 446058 121222 446294
rect 121306 446058 121542 446294
rect 120986 410378 121222 410614
rect 121306 410378 121542 410614
rect 120986 410058 121222 410294
rect 121306 410058 121542 410294
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 120986 122378 121222 122614
rect 121306 122378 121542 122614
rect 120986 122058 121222 122294
rect 121306 122058 121542 122294
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 120986 -3462 121222 -3226
rect 121306 -3462 121542 -3226
rect 120986 -3782 121222 -3546
rect 121306 -3782 121542 -3546
rect 124706 558098 124942 558334
rect 125026 558098 125262 558334
rect 124706 557778 124942 558014
rect 125026 557778 125262 558014
rect 124706 522098 124942 522334
rect 125026 522098 125262 522334
rect 124706 521778 124942 522014
rect 125026 521778 125262 522014
rect 128426 525818 128662 526054
rect 128746 525818 128982 526054
rect 128426 525498 128662 525734
rect 128746 525498 128982 525734
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 124706 486098 124942 486334
rect 125026 486098 125262 486334
rect 124706 485778 124942 486014
rect 125026 485778 125262 486014
rect 128426 489818 128662 490054
rect 128746 489818 128982 490054
rect 128426 489498 128662 489734
rect 128746 489498 128982 489734
rect 125690 471218 125926 471454
rect 125690 470898 125926 471134
rect 124706 450098 124942 450334
rect 125026 450098 125262 450334
rect 124706 449778 124942 450014
rect 125026 449778 125262 450014
rect 128426 453818 128662 454054
rect 128746 453818 128982 454054
rect 128426 453498 128662 453734
rect 128746 453498 128982 453734
rect 125690 435218 125926 435454
rect 125690 434898 125926 435134
rect 124706 414098 124942 414334
rect 125026 414098 125262 414334
rect 124706 413778 124942 414014
rect 125026 413778 125262 414014
rect 128426 417818 128662 418054
rect 128746 417818 128982 418054
rect 128426 417498 128662 417734
rect 128746 417498 128982 417734
rect 125690 399218 125926 399454
rect 125690 398898 125926 399134
rect 124706 378098 124942 378334
rect 125026 378098 125262 378334
rect 124706 377778 124942 378014
rect 125026 377778 125262 378014
rect 124706 342098 124942 342334
rect 125026 342098 125262 342334
rect 124706 341778 124942 342014
rect 125026 341778 125262 342014
rect 124706 306098 124942 306334
rect 125026 306098 125262 306334
rect 124706 305778 124942 306014
rect 125026 305778 125262 306014
rect 124706 270098 124942 270334
rect 125026 270098 125262 270334
rect 124706 269778 124942 270014
rect 125026 269778 125262 270014
rect 124706 234098 124942 234334
rect 125026 234098 125262 234334
rect 124706 233778 124942 234014
rect 125026 233778 125262 234014
rect 124706 198098 124942 198334
rect 125026 198098 125262 198334
rect 124706 197778 124942 198014
rect 125026 197778 125262 198014
rect 124706 162098 124942 162334
rect 125026 162098 125262 162334
rect 124706 161778 124942 162014
rect 125026 161778 125262 162014
rect 128426 381818 128662 382054
rect 128746 381818 128982 382054
rect 128426 381498 128662 381734
rect 128746 381498 128982 381734
rect 128426 345818 128662 346054
rect 128746 345818 128982 346054
rect 128426 345498 128662 345734
rect 128746 345498 128982 345734
rect 128426 309818 128662 310054
rect 128746 309818 128982 310054
rect 128426 309498 128662 309734
rect 128746 309498 128982 309734
rect 128426 273818 128662 274054
rect 128746 273818 128982 274054
rect 128426 273498 128662 273734
rect 128746 273498 128982 273734
rect 128426 237818 128662 238054
rect 128746 237818 128982 238054
rect 128426 237498 128662 237734
rect 128746 237498 128982 237734
rect 128426 201818 128662 202054
rect 128746 201818 128982 202054
rect 128426 201498 128662 201734
rect 128746 201498 128982 201734
rect 128426 165818 128662 166054
rect 128746 165818 128982 166054
rect 128426 165498 128662 165734
rect 128746 165498 128982 165734
rect 124706 126098 124942 126334
rect 125026 126098 125262 126334
rect 124706 125778 124942 126014
rect 125026 125778 125262 126014
rect 128426 129818 128662 130054
rect 128746 129818 128982 130054
rect 128426 129498 128662 129734
rect 128746 129498 128982 129734
rect 124706 90098 124942 90334
rect 125026 90098 125262 90334
rect 124706 89778 124942 90014
rect 125026 89778 125262 90014
rect 124706 54098 124942 54334
rect 125026 54098 125262 54334
rect 124706 53778 124942 54014
rect 125026 53778 125262 54014
rect 124706 18098 124942 18334
rect 125026 18098 125262 18334
rect 124706 17778 124942 18014
rect 125026 17778 125262 18014
rect 124706 -4422 124942 -4186
rect 125026 -4422 125262 -4186
rect 124706 -4742 124942 -4506
rect 125026 -4742 125262 -4506
rect 128426 93818 128662 94054
rect 128746 93818 128982 94054
rect 128426 93498 128662 93734
rect 128746 93498 128982 93734
rect 128426 57818 128662 58054
rect 128746 57818 128982 58054
rect 128426 57498 128662 57734
rect 128746 57498 128982 57734
rect 128426 21818 128662 22054
rect 128746 21818 128982 22054
rect 128426 21498 128662 21734
rect 128746 21498 128982 21734
rect 128426 -5382 128662 -5146
rect 128746 -5382 128982 -5146
rect 128426 -5702 128662 -5466
rect 128746 -5702 128982 -5466
rect 132146 529538 132382 529774
rect 132466 529538 132702 529774
rect 132146 529218 132382 529454
rect 132466 529218 132702 529454
rect 132146 493538 132382 493774
rect 132466 493538 132702 493774
rect 132146 493218 132382 493454
rect 132466 493218 132702 493454
rect 132146 457538 132382 457774
rect 132466 457538 132702 457774
rect 132146 457218 132382 457454
rect 132466 457218 132702 457454
rect 132146 421538 132382 421774
rect 132466 421538 132702 421774
rect 132146 421218 132382 421454
rect 132466 421218 132702 421454
rect 132146 385538 132382 385774
rect 132466 385538 132702 385774
rect 132146 385218 132382 385454
rect 132466 385218 132702 385454
rect 132146 349538 132382 349774
rect 132466 349538 132702 349774
rect 132146 349218 132382 349454
rect 132466 349218 132702 349454
rect 132146 313538 132382 313774
rect 132466 313538 132702 313774
rect 132146 313218 132382 313454
rect 132466 313218 132702 313454
rect 132146 277538 132382 277774
rect 132466 277538 132702 277774
rect 132146 277218 132382 277454
rect 132466 277218 132702 277454
rect 132146 241538 132382 241774
rect 132466 241538 132702 241774
rect 132146 241218 132382 241454
rect 132466 241218 132702 241454
rect 132146 205538 132382 205774
rect 132466 205538 132702 205774
rect 132146 205218 132382 205454
rect 132466 205218 132702 205454
rect 135866 533258 136102 533494
rect 136186 533258 136422 533494
rect 135866 532938 136102 533174
rect 136186 532938 136422 533174
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 141050 510938 141286 511174
rect 141050 510618 141286 510854
rect 135866 497258 136102 497494
rect 136186 497258 136422 497494
rect 135866 496938 136102 497174
rect 136186 496938 136422 497174
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 141050 474938 141286 475174
rect 141050 474618 141286 474854
rect 135866 461258 136102 461494
rect 136186 461258 136422 461494
rect 135866 460938 136102 461174
rect 136186 460938 136422 461174
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 141050 438938 141286 439174
rect 141050 438618 141286 438854
rect 135866 425258 136102 425494
rect 136186 425258 136422 425494
rect 135866 424938 136102 425174
rect 136186 424938 136422 425174
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 141050 402938 141286 403174
rect 141050 402618 141286 402854
rect 135866 389258 136102 389494
rect 136186 389258 136422 389494
rect 135866 388938 136102 389174
rect 136186 388938 136422 389174
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 135866 353258 136102 353494
rect 136186 353258 136422 353494
rect 135866 352938 136102 353174
rect 136186 352938 136422 353174
rect 135866 317258 136102 317494
rect 136186 317258 136422 317494
rect 135866 316938 136102 317174
rect 136186 316938 136422 317174
rect 135866 281258 136102 281494
rect 136186 281258 136422 281494
rect 135866 280938 136102 281174
rect 136186 280938 136422 281174
rect 135866 245258 136102 245494
rect 136186 245258 136422 245494
rect 135866 244938 136102 245174
rect 136186 244938 136422 245174
rect 135866 209258 136102 209494
rect 136186 209258 136422 209494
rect 135866 208938 136102 209174
rect 136186 208938 136422 209174
rect 132146 169538 132382 169774
rect 132466 169538 132702 169774
rect 135866 173258 136102 173494
rect 136186 173258 136422 173494
rect 135866 172938 136102 173174
rect 136186 172938 136422 173174
rect 132146 169218 132382 169454
rect 132466 169218 132702 169454
rect 132146 133538 132382 133774
rect 132466 133538 132702 133774
rect 132146 133218 132382 133454
rect 132466 133218 132702 133454
rect 132146 97538 132382 97774
rect 132466 97538 132702 97774
rect 132146 97218 132382 97454
rect 132466 97218 132702 97454
rect 132146 61538 132382 61774
rect 132466 61538 132702 61774
rect 132146 61218 132382 61454
rect 132466 61218 132702 61454
rect 132146 25538 132382 25774
rect 132466 25538 132702 25774
rect 132146 25218 132382 25454
rect 132466 25218 132702 25454
rect 132146 -6342 132382 -6106
rect 132466 -6342 132702 -6106
rect 132146 -6662 132382 -6426
rect 132466 -6662 132702 -6426
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 135866 137258 136102 137494
rect 136186 137258 136422 137494
rect 135866 136938 136102 137174
rect 136186 136938 136422 137174
rect 135866 101258 136102 101494
rect 136186 101258 136422 101494
rect 135866 100938 136102 101174
rect 136186 100938 136422 101174
rect 135866 65258 136102 65494
rect 136186 65258 136422 65494
rect 135866 64938 136102 65174
rect 136186 64938 136422 65174
rect 135866 29258 136102 29494
rect 136186 29258 136422 29494
rect 135866 28938 136102 29174
rect 136186 28938 136422 29174
rect 135866 -7302 136102 -7066
rect 136186 -7302 136422 -7066
rect 135866 -7622 136102 -7386
rect 136186 -7622 136422 -7386
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 145826 111218 146062 111454
rect 146146 111218 146382 111454
rect 145826 110898 146062 111134
rect 146146 110898 146382 111134
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 705562 149782 705798
rect 149866 705562 150102 705798
rect 149546 705242 149782 705478
rect 149866 705242 150102 705478
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 149546 114938 149782 115174
rect 149866 114938 150102 115174
rect 149546 114618 149782 114854
rect 149866 114618 150102 114854
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -1542 149782 -1306
rect 149866 -1542 150102 -1306
rect 149546 -1862 149782 -1626
rect 149866 -1862 150102 -1626
rect 153266 706522 153502 706758
rect 153586 706522 153822 706758
rect 153266 706202 153502 706438
rect 153586 706202 153822 706438
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 156986 707482 157222 707718
rect 157306 707482 157542 707718
rect 156986 707162 157222 707398
rect 157306 707162 157542 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 156410 471218 156646 471454
rect 156410 470898 156646 471134
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156410 435218 156646 435454
rect 156410 434898 156646 435134
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156410 399218 156646 399454
rect 156410 398898 156646 399134
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 153266 118658 153502 118894
rect 153586 118658 153822 118894
rect 153266 118338 153502 118574
rect 153586 118338 153822 118574
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -2502 153502 -2266
rect 153586 -2502 153822 -2266
rect 153266 -2822 153502 -2586
rect 153586 -2822 153822 -2586
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 156986 122378 157222 122614
rect 157306 122378 157542 122614
rect 156986 122058 157222 122294
rect 157306 122058 157542 122294
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 156986 -3462 157222 -3226
rect 157306 -3462 157542 -3226
rect 156986 -3782 157222 -3546
rect 157306 -3782 157542 -3546
rect 160706 708442 160942 708678
rect 161026 708442 161262 708678
rect 160706 708122 160942 708358
rect 161026 708122 161262 708358
rect 160706 666098 160942 666334
rect 161026 666098 161262 666334
rect 160706 665778 160942 666014
rect 161026 665778 161262 666014
rect 160706 630098 160942 630334
rect 161026 630098 161262 630334
rect 160706 629778 160942 630014
rect 161026 629778 161262 630014
rect 160706 594098 160942 594334
rect 161026 594098 161262 594334
rect 160706 593778 160942 594014
rect 161026 593778 161262 594014
rect 160706 558098 160942 558334
rect 161026 558098 161262 558334
rect 160706 557778 160942 558014
rect 161026 557778 161262 558014
rect 160706 522098 160942 522334
rect 161026 522098 161262 522334
rect 160706 521778 160942 522014
rect 161026 521778 161262 522014
rect 160706 486098 160942 486334
rect 161026 486098 161262 486334
rect 160706 485778 160942 486014
rect 161026 485778 161262 486014
rect 160706 450098 160942 450334
rect 161026 450098 161262 450334
rect 160706 449778 160942 450014
rect 161026 449778 161262 450014
rect 160706 414098 160942 414334
rect 161026 414098 161262 414334
rect 160706 413778 160942 414014
rect 161026 413778 161262 414014
rect 160706 378098 160942 378334
rect 161026 378098 161262 378334
rect 160706 377778 160942 378014
rect 161026 377778 161262 378014
rect 160706 342098 160942 342334
rect 161026 342098 161262 342334
rect 160706 341778 160942 342014
rect 161026 341778 161262 342014
rect 160706 306098 160942 306334
rect 161026 306098 161262 306334
rect 160706 305778 160942 306014
rect 161026 305778 161262 306014
rect 160706 270098 160942 270334
rect 161026 270098 161262 270334
rect 160706 269778 160942 270014
rect 161026 269778 161262 270014
rect 160706 234098 160942 234334
rect 161026 234098 161262 234334
rect 160706 233778 160942 234014
rect 161026 233778 161262 234014
rect 160706 198098 160942 198334
rect 161026 198098 161262 198334
rect 160706 197778 160942 198014
rect 161026 197778 161262 198014
rect 160706 162098 160942 162334
rect 161026 162098 161262 162334
rect 160706 161778 160942 162014
rect 161026 161778 161262 162014
rect 160706 126098 160942 126334
rect 161026 126098 161262 126334
rect 160706 125778 160942 126014
rect 161026 125778 161262 126014
rect 160706 90098 160942 90334
rect 161026 90098 161262 90334
rect 160706 89778 160942 90014
rect 161026 89778 161262 90014
rect 160706 54098 160942 54334
rect 161026 54098 161262 54334
rect 160706 53778 160942 54014
rect 161026 53778 161262 54014
rect 160706 18098 160942 18334
rect 161026 18098 161262 18334
rect 160706 17778 160942 18014
rect 161026 17778 161262 18014
rect 160706 -4422 160942 -4186
rect 161026 -4422 161262 -4186
rect 160706 -4742 160942 -4506
rect 161026 -4742 161262 -4506
rect 164426 709402 164662 709638
rect 164746 709402 164982 709638
rect 164426 709082 164662 709318
rect 164746 709082 164982 709318
rect 164426 669818 164662 670054
rect 164746 669818 164982 670054
rect 164426 669498 164662 669734
rect 164746 669498 164982 669734
rect 164426 633818 164662 634054
rect 164746 633818 164982 634054
rect 164426 633498 164662 633734
rect 164746 633498 164982 633734
rect 168146 710362 168382 710598
rect 168466 710362 168702 710598
rect 168146 710042 168382 710278
rect 168466 710042 168702 710278
rect 168146 673538 168382 673774
rect 168466 673538 168702 673774
rect 168146 673218 168382 673454
rect 168466 673218 168702 673454
rect 168146 637538 168382 637774
rect 168466 637538 168702 637774
rect 168146 637218 168382 637454
rect 168466 637218 168702 637454
rect 164426 597818 164662 598054
rect 164746 597818 164982 598054
rect 164426 597498 164662 597734
rect 164746 597498 164982 597734
rect 164426 561818 164662 562054
rect 164746 561818 164982 562054
rect 164426 561498 164662 561734
rect 164746 561498 164982 561734
rect 168146 601538 168382 601774
rect 168466 601538 168702 601774
rect 168146 601218 168382 601454
rect 168466 601218 168702 601454
rect 171866 711322 172102 711558
rect 172186 711322 172422 711558
rect 171866 711002 172102 711238
rect 172186 711002 172422 711238
rect 171866 677258 172102 677494
rect 172186 677258 172422 677494
rect 171866 676938 172102 677174
rect 172186 676938 172422 677174
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 171866 641258 172102 641494
rect 172186 641258 172422 641494
rect 171866 640938 172102 641174
rect 172186 640938 172422 641174
rect 171866 605258 172102 605494
rect 172186 605258 172422 605494
rect 171866 604938 172102 605174
rect 172186 604938 172422 605174
rect 168146 565538 168382 565774
rect 168466 565538 168702 565774
rect 168146 565218 168382 565454
rect 168466 565218 168702 565454
rect 164426 525818 164662 526054
rect 164746 525818 164982 526054
rect 164426 525498 164662 525734
rect 164746 525498 164982 525734
rect 164426 489818 164662 490054
rect 164746 489818 164982 490054
rect 164426 489498 164662 489734
rect 164746 489498 164982 489734
rect 164426 453818 164662 454054
rect 164746 453818 164982 454054
rect 164426 453498 164662 453734
rect 164746 453498 164982 453734
rect 164426 417818 164662 418054
rect 164746 417818 164982 418054
rect 164426 417498 164662 417734
rect 164746 417498 164982 417734
rect 164426 381818 164662 382054
rect 164746 381818 164982 382054
rect 164426 381498 164662 381734
rect 164746 381498 164982 381734
rect 164426 345818 164662 346054
rect 164746 345818 164982 346054
rect 164426 345498 164662 345734
rect 164746 345498 164982 345734
rect 164426 309818 164662 310054
rect 164746 309818 164982 310054
rect 164426 309498 164662 309734
rect 164746 309498 164982 309734
rect 164426 273818 164662 274054
rect 164746 273818 164982 274054
rect 164426 273498 164662 273734
rect 164746 273498 164982 273734
rect 164426 237818 164662 238054
rect 164746 237818 164982 238054
rect 164426 237498 164662 237734
rect 164746 237498 164982 237734
rect 164426 201818 164662 202054
rect 164746 201818 164982 202054
rect 164426 201498 164662 201734
rect 164746 201498 164982 201734
rect 164426 165818 164662 166054
rect 164746 165818 164982 166054
rect 164426 165498 164662 165734
rect 164746 165498 164982 165734
rect 164426 129818 164662 130054
rect 164746 129818 164982 130054
rect 164426 129498 164662 129734
rect 164746 129498 164982 129734
rect 164426 93818 164662 94054
rect 164746 93818 164982 94054
rect 164426 93498 164662 93734
rect 164746 93498 164982 93734
rect 164426 57818 164662 58054
rect 164746 57818 164982 58054
rect 164426 57498 164662 57734
rect 164746 57498 164982 57734
rect 164426 21818 164662 22054
rect 164746 21818 164982 22054
rect 164426 21498 164662 21734
rect 164746 21498 164982 21734
rect 164426 -5382 164662 -5146
rect 164746 -5382 164982 -5146
rect 164426 -5702 164662 -5466
rect 164746 -5702 164982 -5466
rect 171866 569258 172102 569494
rect 172186 569258 172422 569494
rect 171866 568938 172102 569174
rect 172186 568938 172422 569174
rect 168146 529538 168382 529774
rect 168466 529538 168702 529774
rect 168146 529218 168382 529454
rect 168466 529218 168702 529454
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 705562 185782 705798
rect 185866 705562 186102 705798
rect 185546 705242 185782 705478
rect 185866 705242 186102 705478
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 706522 189502 706758
rect 189586 706522 189822 706758
rect 189266 706202 189502 706438
rect 189586 706202 189822 706438
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 192986 707482 193222 707718
rect 193306 707482 193542 707718
rect 192986 707162 193222 707398
rect 193306 707162 193542 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 196706 708442 196942 708678
rect 197026 708442 197262 708678
rect 196706 708122 196942 708358
rect 197026 708122 197262 708358
rect 196706 666098 196942 666334
rect 197026 666098 197262 666334
rect 196706 665778 196942 666014
rect 197026 665778 197262 666014
rect 200426 709402 200662 709638
rect 200746 709402 200982 709638
rect 200426 709082 200662 709318
rect 200746 709082 200982 709318
rect 200426 669818 200662 670054
rect 200746 669818 200982 670054
rect 200426 669498 200662 669734
rect 200746 669498 200982 669734
rect 200426 633818 200662 634054
rect 200746 633818 200982 634054
rect 200426 633498 200662 633734
rect 200746 633498 200982 633734
rect 204146 710362 204382 710598
rect 204466 710362 204702 710598
rect 204146 710042 204382 710278
rect 204466 710042 204702 710278
rect 204146 673538 204382 673774
rect 204466 673538 204702 673774
rect 204146 673218 204382 673454
rect 204466 673218 204702 673454
rect 204146 637538 204382 637774
rect 204466 637538 204702 637774
rect 204146 637218 204382 637454
rect 204466 637218 204702 637454
rect 207866 711322 208102 711558
rect 208186 711322 208422 711558
rect 207866 711002 208102 711238
rect 208186 711002 208422 711238
rect 207866 677258 208102 677494
rect 208186 677258 208422 677494
rect 207866 676938 208102 677174
rect 208186 676938 208422 677174
rect 207866 641258 208102 641494
rect 208186 641258 208422 641494
rect 207866 640938 208102 641174
rect 208186 640938 208422 641174
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 705562 221782 705798
rect 221866 705562 222102 705798
rect 221546 705242 221782 705478
rect 221866 705242 222102 705478
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 706522 225502 706758
rect 225586 706522 225822 706758
rect 225266 706202 225502 706438
rect 225586 706202 225822 706438
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 228986 707482 229222 707718
rect 229306 707482 229542 707718
rect 228986 707162 229222 707398
rect 229306 707162 229542 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 232706 708442 232942 708678
rect 233026 708442 233262 708678
rect 232706 708122 232942 708358
rect 233026 708122 233262 708358
rect 232706 666098 232942 666334
rect 233026 666098 233262 666334
rect 232706 665778 232942 666014
rect 233026 665778 233262 666014
rect 236426 709402 236662 709638
rect 236746 709402 236982 709638
rect 236426 709082 236662 709318
rect 236746 709082 236982 709318
rect 236426 669818 236662 670054
rect 236746 669818 236982 670054
rect 236426 669498 236662 669734
rect 236746 669498 236982 669734
rect 236426 633818 236662 634054
rect 236746 633818 236982 634054
rect 236426 633498 236662 633734
rect 236746 633498 236982 633734
rect 240146 710362 240382 710598
rect 240466 710362 240702 710598
rect 240146 710042 240382 710278
rect 240466 710042 240702 710278
rect 240146 673538 240382 673774
rect 240466 673538 240702 673774
rect 240146 673218 240382 673454
rect 240466 673218 240702 673454
rect 240146 637538 240382 637774
rect 240466 637538 240702 637774
rect 240146 637218 240382 637454
rect 240466 637218 240702 637454
rect 243866 711322 244102 711558
rect 244186 711322 244422 711558
rect 243866 711002 244102 711238
rect 244186 711002 244422 711238
rect 243866 677258 244102 677494
rect 244186 677258 244422 677494
rect 243866 676938 244102 677174
rect 244186 676938 244422 677174
rect 243866 641258 244102 641494
rect 244186 641258 244422 641494
rect 243866 640938 244102 641174
rect 244186 640938 244422 641174
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 705562 257782 705798
rect 257866 705562 258102 705798
rect 257546 705242 257782 705478
rect 257866 705242 258102 705478
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 199610 618938 199846 619174
rect 199610 618618 199846 618854
rect 230330 618938 230566 619174
rect 230330 618618 230566 618854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 184250 615218 184486 615454
rect 184250 614898 184486 615134
rect 214970 615218 215206 615454
rect 214970 614898 215206 615134
rect 245690 615218 245926 615454
rect 245690 614898 245926 615134
rect 171866 533258 172102 533494
rect 172186 533258 172422 533494
rect 171866 532938 172102 533174
rect 172186 532938 172422 533174
rect 199610 582938 199846 583174
rect 199610 582618 199846 582854
rect 230330 582938 230566 583174
rect 230330 582618 230566 582854
rect 184250 579218 184486 579454
rect 184250 578898 184486 579134
rect 214970 579218 215206 579454
rect 214970 578898 215206 579134
rect 245690 579218 245926 579454
rect 245690 578898 245926 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 171770 510938 172006 511174
rect 171770 510618 172006 510854
rect 168146 493538 168382 493774
rect 168466 493538 168702 493774
rect 168146 493218 168382 493454
rect 168466 493218 168702 493454
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 171770 474938 172006 475174
rect 171770 474618 172006 474854
rect 168146 457538 168382 457774
rect 168466 457538 168702 457774
rect 168146 457218 168382 457454
rect 168466 457218 168702 457454
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 171770 438938 172006 439174
rect 171770 438618 172006 438854
rect 168146 421538 168382 421774
rect 168466 421538 168702 421774
rect 168146 421218 168382 421454
rect 168466 421218 168702 421454
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 171770 402938 172006 403174
rect 171770 402618 172006 402854
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 168146 385538 168382 385774
rect 168466 385538 168702 385774
rect 168146 385218 168382 385454
rect 168466 385218 168702 385454
rect 168146 349538 168382 349774
rect 168466 349538 168702 349774
rect 168146 349218 168382 349454
rect 168466 349218 168702 349454
rect 168146 313538 168382 313774
rect 168466 313538 168702 313774
rect 168146 313218 168382 313454
rect 168466 313218 168702 313454
rect 168146 277538 168382 277774
rect 168466 277538 168702 277774
rect 168146 277218 168382 277454
rect 168466 277218 168702 277454
rect 168146 241538 168382 241774
rect 168466 241538 168702 241774
rect 168146 241218 168382 241454
rect 168466 241218 168702 241454
rect 168146 205538 168382 205774
rect 168466 205538 168702 205774
rect 168146 205218 168382 205454
rect 168466 205218 168702 205454
rect 168146 169538 168382 169774
rect 168466 169538 168702 169774
rect 168146 169218 168382 169454
rect 168466 169218 168702 169454
rect 168146 133538 168382 133774
rect 168466 133538 168702 133774
rect 168146 133218 168382 133454
rect 168466 133218 168702 133454
rect 168146 97538 168382 97774
rect 168466 97538 168702 97774
rect 168146 97218 168382 97454
rect 168466 97218 168702 97454
rect 168146 61538 168382 61774
rect 168466 61538 168702 61774
rect 168146 61218 168382 61454
rect 168466 61218 168702 61454
rect 168146 25538 168382 25774
rect 168466 25538 168702 25774
rect 168146 25218 168382 25454
rect 168466 25218 168702 25454
rect 168146 -6342 168382 -6106
rect 168466 -6342 168702 -6106
rect 168146 -6662 168382 -6426
rect 168466 -6662 168702 -6426
rect 171866 389258 172102 389494
rect 172186 389258 172422 389494
rect 171866 388938 172102 389174
rect 172186 388938 172422 389174
rect 171866 353258 172102 353494
rect 172186 353258 172422 353494
rect 171866 352938 172102 353174
rect 172186 352938 172422 353174
rect 171866 317258 172102 317494
rect 172186 317258 172422 317494
rect 171866 316938 172102 317174
rect 172186 316938 172422 317174
rect 171866 281258 172102 281494
rect 172186 281258 172422 281494
rect 171866 280938 172102 281174
rect 172186 280938 172422 281174
rect 171866 245258 172102 245494
rect 172186 245258 172422 245494
rect 171866 244938 172102 245174
rect 172186 244938 172422 245174
rect 171866 209258 172102 209494
rect 172186 209258 172422 209494
rect 171866 208938 172102 209174
rect 172186 208938 172422 209174
rect 171866 173258 172102 173494
rect 172186 173258 172422 173494
rect 171866 172938 172102 173174
rect 172186 172938 172422 173174
rect 171866 137258 172102 137494
rect 172186 137258 172422 137494
rect 171866 136938 172102 137174
rect 172186 136938 172422 137174
rect 171866 101258 172102 101494
rect 172186 101258 172422 101494
rect 171866 100938 172102 101174
rect 172186 100938 172422 101174
rect 171866 65258 172102 65494
rect 172186 65258 172422 65494
rect 171866 64938 172102 65174
rect 172186 64938 172422 65174
rect 171866 29258 172102 29494
rect 172186 29258 172422 29494
rect 171866 28938 172102 29174
rect 172186 28938 172422 29174
rect 171866 -7302 172102 -7066
rect 172186 -7302 172422 -7066
rect 171866 -7622 172102 -7386
rect 172186 -7622 172422 -7386
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 187130 471218 187366 471454
rect 187130 470898 187366 471134
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 187130 435218 187366 435454
rect 187130 434898 187366 435134
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 187130 399218 187366 399454
rect 187130 398898 187366 399134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -1542 185782 -1306
rect 185866 -1542 186102 -1306
rect 185546 -1862 185782 -1626
rect 185866 -1862 186102 -1626
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -2502 189502 -2266
rect 189586 -2502 189822 -2266
rect 189266 -2822 189502 -2586
rect 189586 -2822 189822 -2586
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 192986 -3462 193222 -3226
rect 193306 -3462 193542 -3226
rect 192986 -3782 193222 -3546
rect 193306 -3782 193542 -3546
rect 196706 558098 196942 558334
rect 197026 558098 197262 558334
rect 196706 557778 196942 558014
rect 197026 557778 197262 558014
rect 196706 522098 196942 522334
rect 197026 522098 197262 522334
rect 232706 558098 232942 558334
rect 233026 558098 233262 558334
rect 232706 557778 232942 558014
rect 233026 557778 233262 558014
rect 196706 521778 196942 522014
rect 197026 521778 197262 522014
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 261266 706522 261502 706758
rect 261586 706522 261822 706758
rect 261266 706202 261502 706438
rect 261586 706202 261822 706438
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 264986 707482 265222 707718
rect 265306 707482 265542 707718
rect 264986 707162 265222 707398
rect 265306 707162 265542 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 268706 708442 268942 708678
rect 269026 708442 269262 708678
rect 268706 708122 268942 708358
rect 269026 708122 269262 708358
rect 268706 666098 268942 666334
rect 269026 666098 269262 666334
rect 268706 665778 268942 666014
rect 269026 665778 269262 666014
rect 268706 630098 268942 630334
rect 269026 630098 269262 630334
rect 268706 629778 268942 630014
rect 269026 629778 269262 630014
rect 268706 594098 268942 594334
rect 269026 594098 269262 594334
rect 268706 593778 268942 594014
rect 269026 593778 269262 594014
rect 268706 558098 268942 558334
rect 269026 558098 269262 558334
rect 268706 557778 268942 558014
rect 269026 557778 269262 558014
rect 272426 709402 272662 709638
rect 272746 709402 272982 709638
rect 272426 709082 272662 709318
rect 272746 709082 272982 709318
rect 272426 669818 272662 670054
rect 272746 669818 272982 670054
rect 272426 669498 272662 669734
rect 272746 669498 272982 669734
rect 272426 633818 272662 634054
rect 272746 633818 272982 634054
rect 272426 633498 272662 633734
rect 272746 633498 272982 633734
rect 272426 597818 272662 598054
rect 272746 597818 272982 598054
rect 272426 597498 272662 597734
rect 272746 597498 272982 597734
rect 272426 561818 272662 562054
rect 272746 561818 272982 562054
rect 272426 561498 272662 561734
rect 272746 561498 272982 561734
rect 272426 525818 272662 526054
rect 272746 525818 272982 526054
rect 272426 525498 272662 525734
rect 272746 525498 272982 525734
rect 276146 710362 276382 710598
rect 276466 710362 276702 710598
rect 276146 710042 276382 710278
rect 276466 710042 276702 710278
rect 276146 673538 276382 673774
rect 276466 673538 276702 673774
rect 276146 673218 276382 673454
rect 276466 673218 276702 673454
rect 276146 637538 276382 637774
rect 276466 637538 276702 637774
rect 276146 637218 276382 637454
rect 276466 637218 276702 637454
rect 276146 601538 276382 601774
rect 276466 601538 276702 601774
rect 276146 601218 276382 601454
rect 276466 601218 276702 601454
rect 276146 565538 276382 565774
rect 276466 565538 276702 565774
rect 276146 565218 276382 565454
rect 276466 565218 276702 565454
rect 276146 529538 276382 529774
rect 276466 529538 276702 529774
rect 276146 529218 276382 529454
rect 276466 529218 276702 529454
rect 279866 711322 280102 711558
rect 280186 711322 280422 711558
rect 279866 711002 280102 711238
rect 280186 711002 280422 711238
rect 279866 677258 280102 677494
rect 280186 677258 280422 677494
rect 279866 676938 280102 677174
rect 280186 676938 280422 677174
rect 279866 641258 280102 641494
rect 280186 641258 280422 641494
rect 279866 640938 280102 641174
rect 280186 640938 280422 641174
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 279866 605258 280102 605494
rect 280186 605258 280422 605494
rect 279866 604938 280102 605174
rect 280186 604938 280422 605174
rect 279866 569258 280102 569494
rect 280186 569258 280422 569494
rect 279866 568938 280102 569174
rect 280186 568938 280422 569174
rect 279866 533258 280102 533494
rect 280186 533258 280422 533494
rect 279866 532938 280102 533174
rect 280186 532938 280422 533174
rect 293546 705562 293782 705798
rect 293866 705562 294102 705798
rect 293546 705242 293782 705478
rect 293866 705242 294102 705478
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 297266 706522 297502 706758
rect 297586 706522 297822 706758
rect 297266 706202 297502 706438
rect 297586 706202 297822 706438
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 300986 707482 301222 707718
rect 301306 707482 301542 707718
rect 300986 707162 301222 707398
rect 301306 707162 301542 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 304706 708442 304942 708678
rect 305026 708442 305262 708678
rect 304706 708122 304942 708358
rect 305026 708122 305262 708358
rect 304706 666098 304942 666334
rect 305026 666098 305262 666334
rect 304706 665778 304942 666014
rect 305026 665778 305262 666014
rect 308426 709402 308662 709638
rect 308746 709402 308982 709638
rect 308426 709082 308662 709318
rect 308746 709082 308982 709318
rect 308426 669818 308662 670054
rect 308746 669818 308982 670054
rect 308426 669498 308662 669734
rect 308746 669498 308982 669734
rect 308426 633818 308662 634054
rect 308746 633818 308982 634054
rect 308426 633498 308662 633734
rect 308746 633498 308982 633734
rect 312146 710362 312382 710598
rect 312466 710362 312702 710598
rect 312146 710042 312382 710278
rect 312466 710042 312702 710278
rect 312146 673538 312382 673774
rect 312466 673538 312702 673774
rect 312146 673218 312382 673454
rect 312466 673218 312702 673454
rect 312146 637538 312382 637774
rect 312466 637538 312702 637774
rect 312146 637218 312382 637454
rect 312466 637218 312702 637454
rect 315866 711322 316102 711558
rect 316186 711322 316422 711558
rect 315866 711002 316102 711238
rect 316186 711002 316422 711238
rect 315866 677258 316102 677494
rect 316186 677258 316422 677494
rect 315866 676938 316102 677174
rect 316186 676938 316422 677174
rect 315866 641258 316102 641494
rect 316186 641258 316422 641494
rect 315866 640938 316102 641174
rect 316186 640938 316422 641174
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 705562 329782 705798
rect 329866 705562 330102 705798
rect 329546 705242 329782 705478
rect 329866 705242 330102 705478
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 706522 333502 706758
rect 333586 706522 333822 706758
rect 333266 706202 333502 706438
rect 333586 706202 333822 706438
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 336986 707482 337222 707718
rect 337306 707482 337542 707718
rect 336986 707162 337222 707398
rect 337306 707162 337542 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 340706 708442 340942 708678
rect 341026 708442 341262 708678
rect 340706 708122 340942 708358
rect 341026 708122 341262 708358
rect 340706 666098 340942 666334
rect 341026 666098 341262 666334
rect 340706 665778 340942 666014
rect 341026 665778 341262 666014
rect 344426 709402 344662 709638
rect 344746 709402 344982 709638
rect 344426 709082 344662 709318
rect 344746 709082 344982 709318
rect 344426 669818 344662 670054
rect 344746 669818 344982 670054
rect 344426 669498 344662 669734
rect 344746 669498 344982 669734
rect 344426 633818 344662 634054
rect 344746 633818 344982 634054
rect 344426 633498 344662 633734
rect 344746 633498 344982 633734
rect 348146 710362 348382 710598
rect 348466 710362 348702 710598
rect 348146 710042 348382 710278
rect 348466 710042 348702 710278
rect 348146 673538 348382 673774
rect 348466 673538 348702 673774
rect 348146 673218 348382 673454
rect 348466 673218 348702 673454
rect 348146 637538 348382 637774
rect 348466 637538 348702 637774
rect 348146 637218 348382 637454
rect 348466 637218 348702 637454
rect 351866 711322 352102 711558
rect 352186 711322 352422 711558
rect 351866 711002 352102 711238
rect 352186 711002 352422 711238
rect 351866 677258 352102 677494
rect 352186 677258 352422 677494
rect 351866 676938 352102 677174
rect 352186 676938 352422 677174
rect 351866 641258 352102 641494
rect 352186 641258 352422 641494
rect 351866 640938 352102 641174
rect 352186 640938 352422 641174
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 705562 365782 705798
rect 365866 705562 366102 705798
rect 365546 705242 365782 705478
rect 365866 705242 366102 705478
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 706522 369502 706758
rect 369586 706522 369822 706758
rect 369266 706202 369502 706438
rect 369586 706202 369822 706438
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 372986 707482 373222 707718
rect 373306 707482 373542 707718
rect 372986 707162 373222 707398
rect 373306 707162 373542 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 376706 708442 376942 708678
rect 377026 708442 377262 708678
rect 376706 708122 376942 708358
rect 377026 708122 377262 708358
rect 376706 666098 376942 666334
rect 377026 666098 377262 666334
rect 376706 665778 376942 666014
rect 377026 665778 377262 666014
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 380426 709402 380662 709638
rect 380746 709402 380982 709638
rect 380426 709082 380662 709318
rect 380746 709082 380982 709318
rect 380426 669818 380662 670054
rect 380746 669818 380982 670054
rect 380426 669498 380662 669734
rect 380746 669498 380982 669734
rect 376706 630098 376942 630334
rect 377026 630098 377262 630334
rect 376706 629778 376942 630014
rect 377026 629778 377262 630014
rect 319610 618938 319846 619174
rect 319610 618618 319846 618854
rect 350330 618938 350566 619174
rect 350330 618618 350566 618854
rect 304250 615218 304486 615454
rect 304250 614898 304486 615134
rect 334970 615218 335206 615454
rect 334970 614898 335206 615134
rect 365690 615218 365926 615454
rect 365690 614898 365926 615134
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 380426 633818 380662 634054
rect 380746 633818 380982 634054
rect 380426 633498 380662 633734
rect 380746 633498 380982 633734
rect 376706 594098 376942 594334
rect 377026 594098 377262 594334
rect 376706 593778 376942 594014
rect 377026 593778 377262 594014
rect 319610 582938 319846 583174
rect 319610 582618 319846 582854
rect 350330 582938 350566 583174
rect 350330 582618 350566 582854
rect 304250 579218 304486 579454
rect 304250 578898 304486 579134
rect 334970 579218 335206 579454
rect 334970 578898 335206 579134
rect 365690 579218 365926 579454
rect 365690 578898 365926 579134
rect 304706 558098 304942 558334
rect 305026 558098 305262 558334
rect 304706 557778 304942 558014
rect 305026 557778 305262 558014
rect 340706 558098 340942 558334
rect 341026 558098 341262 558334
rect 340706 557778 340942 558014
rect 341026 557778 341262 558014
rect 380426 597818 380662 598054
rect 380746 597818 380982 598054
rect 380426 597498 380662 597734
rect 380746 597498 380982 597734
rect 376706 558098 376942 558334
rect 377026 558098 377262 558334
rect 376706 557778 376942 558014
rect 377026 557778 377262 558014
rect 384146 710362 384382 710598
rect 384466 710362 384702 710598
rect 384146 710042 384382 710278
rect 384466 710042 384702 710278
rect 384146 673538 384382 673774
rect 384466 673538 384702 673774
rect 384146 673218 384382 673454
rect 384466 673218 384702 673454
rect 384146 637538 384382 637774
rect 384466 637538 384702 637774
rect 384146 637218 384382 637454
rect 384466 637218 384702 637454
rect 384146 601538 384382 601774
rect 384466 601538 384702 601774
rect 384146 601218 384382 601454
rect 384466 601218 384702 601454
rect 380426 561818 380662 562054
rect 380746 561818 380982 562054
rect 380426 561498 380662 561734
rect 380746 561498 380982 561734
rect 384146 565538 384382 565774
rect 384466 565538 384702 565774
rect 384146 565218 384382 565454
rect 384466 565218 384702 565454
rect 380426 525818 380662 526054
rect 380746 525818 380982 526054
rect 380426 525498 380662 525734
rect 380746 525498 380982 525734
rect 384146 529538 384382 529774
rect 384466 529538 384702 529774
rect 384146 529218 384382 529454
rect 384466 529218 384702 529454
rect 387866 711322 388102 711558
rect 388186 711322 388422 711558
rect 387866 711002 388102 711238
rect 388186 711002 388422 711238
rect 387866 677258 388102 677494
rect 388186 677258 388422 677494
rect 387866 676938 388102 677174
rect 388186 676938 388422 677174
rect 387866 641258 388102 641494
rect 388186 641258 388422 641494
rect 387866 640938 388102 641174
rect 388186 640938 388422 641174
rect 387866 605258 388102 605494
rect 388186 605258 388422 605494
rect 387866 604938 388102 605174
rect 388186 604938 388422 605174
rect 387866 569258 388102 569494
rect 388186 569258 388422 569494
rect 387866 568938 388102 569174
rect 388186 568938 388422 569174
rect 387866 533258 388102 533494
rect 388186 533258 388422 533494
rect 387866 532938 388102 533174
rect 388186 532938 388422 533174
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 401546 705562 401782 705798
rect 401866 705562 402102 705798
rect 401546 705242 401782 705478
rect 401866 705242 402102 705478
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 405266 706522 405502 706758
rect 405586 706522 405822 706758
rect 405266 706202 405502 706438
rect 405586 706202 405822 706438
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 408986 707482 409222 707718
rect 409306 707482 409542 707718
rect 408986 707162 409222 707398
rect 409306 707162 409542 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 412706 708442 412942 708678
rect 413026 708442 413262 708678
rect 412706 708122 412942 708358
rect 413026 708122 413262 708358
rect 412706 666098 412942 666334
rect 413026 666098 413262 666334
rect 412706 665778 412942 666014
rect 413026 665778 413262 666014
rect 412706 630098 412942 630334
rect 413026 630098 413262 630334
rect 412706 629778 412942 630014
rect 413026 629778 413262 630014
rect 412706 594098 412942 594334
rect 413026 594098 413262 594334
rect 412706 593778 412942 594014
rect 413026 593778 413262 594014
rect 412706 558098 412942 558334
rect 413026 558098 413262 558334
rect 412706 557778 412942 558014
rect 413026 557778 413262 558014
rect 416426 709402 416662 709638
rect 416746 709402 416982 709638
rect 416426 709082 416662 709318
rect 416746 709082 416982 709318
rect 416426 669818 416662 670054
rect 416746 669818 416982 670054
rect 416426 669498 416662 669734
rect 416746 669498 416982 669734
rect 416426 633818 416662 634054
rect 416746 633818 416982 634054
rect 416426 633498 416662 633734
rect 416746 633498 416982 633734
rect 416426 597818 416662 598054
rect 416746 597818 416982 598054
rect 416426 597498 416662 597734
rect 416746 597498 416982 597734
rect 416426 561818 416662 562054
rect 416746 561818 416982 562054
rect 416426 561498 416662 561734
rect 416746 561498 416982 561734
rect 416426 525818 416662 526054
rect 416746 525818 416982 526054
rect 416426 525498 416662 525734
rect 416746 525498 416982 525734
rect 420146 710362 420382 710598
rect 420466 710362 420702 710598
rect 420146 710042 420382 710278
rect 420466 710042 420702 710278
rect 420146 673538 420382 673774
rect 420466 673538 420702 673774
rect 420146 673218 420382 673454
rect 420466 673218 420702 673454
rect 420146 637538 420382 637774
rect 420466 637538 420702 637774
rect 420146 637218 420382 637454
rect 420466 637218 420702 637454
rect 420146 601538 420382 601774
rect 420466 601538 420702 601774
rect 420146 601218 420382 601454
rect 420466 601218 420702 601454
rect 420146 565538 420382 565774
rect 420466 565538 420702 565774
rect 420146 565218 420382 565454
rect 420466 565218 420702 565454
rect 420146 529538 420382 529774
rect 420466 529538 420702 529774
rect 420146 529218 420382 529454
rect 420466 529218 420702 529454
rect 423866 711322 424102 711558
rect 424186 711322 424422 711558
rect 423866 711002 424102 711238
rect 424186 711002 424422 711238
rect 423866 677258 424102 677494
rect 424186 677258 424422 677494
rect 423866 676938 424102 677174
rect 424186 676938 424422 677174
rect 423866 641258 424102 641494
rect 424186 641258 424422 641494
rect 423866 640938 424102 641174
rect 424186 640938 424422 641174
rect 423866 605258 424102 605494
rect 424186 605258 424422 605494
rect 423866 604938 424102 605174
rect 424186 604938 424422 605174
rect 423866 569258 424102 569494
rect 424186 569258 424422 569494
rect 423866 568938 424102 569174
rect 424186 568938 424422 569174
rect 423866 533258 424102 533494
rect 424186 533258 424422 533494
rect 423866 532938 424102 533174
rect 424186 532938 424422 533174
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 437546 705562 437782 705798
rect 437866 705562 438102 705798
rect 437546 705242 437782 705478
rect 437866 705242 438102 705478
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 441266 706522 441502 706758
rect 441586 706522 441822 706758
rect 441266 706202 441502 706438
rect 441586 706202 441822 706438
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 444986 707482 445222 707718
rect 445306 707482 445542 707718
rect 444986 707162 445222 707398
rect 445306 707162 445542 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 448706 708442 448942 708678
rect 449026 708442 449262 708678
rect 448706 708122 448942 708358
rect 449026 708122 449262 708358
rect 448706 666098 448942 666334
rect 449026 666098 449262 666334
rect 448706 665778 448942 666014
rect 449026 665778 449262 666014
rect 452426 709402 452662 709638
rect 452746 709402 452982 709638
rect 452426 709082 452662 709318
rect 452746 709082 452982 709318
rect 452426 669818 452662 670054
rect 452746 669818 452982 670054
rect 452426 669498 452662 669734
rect 452746 669498 452982 669734
rect 448706 630098 448942 630334
rect 449026 630098 449262 630334
rect 448706 629778 448942 630014
rect 449026 629778 449262 630014
rect 448706 594098 448942 594334
rect 449026 594098 449262 594334
rect 448706 593778 448942 594014
rect 449026 593778 449262 594014
rect 448706 558098 448942 558334
rect 449026 558098 449262 558334
rect 448706 557778 448942 558014
rect 449026 557778 449262 558014
rect 452426 633818 452662 634054
rect 452746 633818 452982 634054
rect 452426 633498 452662 633734
rect 452746 633498 452982 633734
rect 452426 597818 452662 598054
rect 452746 597818 452982 598054
rect 452426 597498 452662 597734
rect 452746 597498 452982 597734
rect 452426 561818 452662 562054
rect 452746 561818 452982 562054
rect 452426 561498 452662 561734
rect 452746 561498 452982 561734
rect 452426 525818 452662 526054
rect 452746 525818 452982 526054
rect 452426 525498 452662 525734
rect 452746 525498 452982 525734
rect 456146 710362 456382 710598
rect 456466 710362 456702 710598
rect 456146 710042 456382 710278
rect 456466 710042 456702 710278
rect 456146 673538 456382 673774
rect 456466 673538 456702 673774
rect 456146 673218 456382 673454
rect 456466 673218 456702 673454
rect 456146 637538 456382 637774
rect 456466 637538 456702 637774
rect 456146 637218 456382 637454
rect 456466 637218 456702 637454
rect 456146 601538 456382 601774
rect 456466 601538 456702 601774
rect 456146 601218 456382 601454
rect 456466 601218 456702 601454
rect 456146 565538 456382 565774
rect 456466 565538 456702 565774
rect 456146 565218 456382 565454
rect 456466 565218 456702 565454
rect 456146 529538 456382 529774
rect 456466 529538 456702 529774
rect 456146 529218 456382 529454
rect 456466 529218 456702 529454
rect 459866 711322 460102 711558
rect 460186 711322 460422 711558
rect 459866 711002 460102 711238
rect 460186 711002 460422 711238
rect 459866 677258 460102 677494
rect 460186 677258 460422 677494
rect 459866 676938 460102 677174
rect 460186 676938 460422 677174
rect 459866 641258 460102 641494
rect 460186 641258 460422 641494
rect 459866 640938 460102 641174
rect 460186 640938 460422 641174
rect 459866 605258 460102 605494
rect 460186 605258 460422 605494
rect 459866 604938 460102 605174
rect 460186 604938 460422 605174
rect 459866 569258 460102 569494
rect 460186 569258 460422 569494
rect 459866 568938 460102 569174
rect 460186 568938 460422 569174
rect 459866 533258 460102 533494
rect 460186 533258 460422 533494
rect 459866 532938 460102 533174
rect 460186 532938 460422 533174
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 473546 705562 473782 705798
rect 473866 705562 474102 705798
rect 473546 705242 473782 705478
rect 473866 705242 474102 705478
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 706522 477502 706758
rect 477586 706522 477822 706758
rect 477266 706202 477502 706438
rect 477586 706202 477822 706438
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 480986 707482 481222 707718
rect 481306 707482 481542 707718
rect 480986 707162 481222 707398
rect 481306 707162 481542 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 484706 708442 484942 708678
rect 485026 708442 485262 708678
rect 484706 708122 484942 708358
rect 485026 708122 485262 708358
rect 484706 666098 484942 666334
rect 485026 666098 485262 666334
rect 484706 665778 484942 666014
rect 485026 665778 485262 666014
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 484706 630098 484942 630334
rect 485026 630098 485262 630334
rect 484706 629778 484942 630014
rect 485026 629778 485262 630014
rect 484706 594098 484942 594334
rect 485026 594098 485262 594334
rect 484706 593778 484942 594014
rect 485026 593778 485262 594014
rect 484706 558098 484942 558334
rect 485026 558098 485262 558334
rect 484706 557778 484942 558014
rect 485026 557778 485262 558014
rect 488426 709402 488662 709638
rect 488746 709402 488982 709638
rect 488426 709082 488662 709318
rect 488746 709082 488982 709318
rect 488426 669818 488662 670054
rect 488746 669818 488982 670054
rect 488426 669498 488662 669734
rect 488746 669498 488982 669734
rect 488426 633818 488662 634054
rect 488746 633818 488982 634054
rect 488426 633498 488662 633734
rect 488746 633498 488982 633734
rect 488426 597818 488662 598054
rect 488746 597818 488982 598054
rect 488426 597498 488662 597734
rect 488746 597498 488982 597734
rect 488426 561818 488662 562054
rect 488746 561818 488982 562054
rect 488426 561498 488662 561734
rect 488746 561498 488982 561734
rect 488426 525818 488662 526054
rect 488746 525818 488982 526054
rect 488426 525498 488662 525734
rect 488746 525498 488982 525734
rect 492146 710362 492382 710598
rect 492466 710362 492702 710598
rect 492146 710042 492382 710278
rect 492466 710042 492702 710278
rect 492146 673538 492382 673774
rect 492466 673538 492702 673774
rect 492146 673218 492382 673454
rect 492466 673218 492702 673454
rect 495866 711322 496102 711558
rect 496186 711322 496422 711558
rect 495866 711002 496102 711238
rect 496186 711002 496422 711238
rect 495866 677258 496102 677494
rect 496186 677258 496422 677494
rect 495866 676938 496102 677174
rect 496186 676938 496422 677174
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 509546 705562 509782 705798
rect 509866 705562 510102 705798
rect 509546 705242 509782 705478
rect 509866 705242 510102 705478
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 513266 706522 513502 706758
rect 513586 706522 513822 706758
rect 513266 706202 513502 706438
rect 513586 706202 513822 706438
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 516986 707482 517222 707718
rect 517306 707482 517542 707718
rect 516986 707162 517222 707398
rect 517306 707162 517542 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 520706 708442 520942 708678
rect 521026 708442 521262 708678
rect 520706 708122 520942 708358
rect 521026 708122 521262 708358
rect 520706 666098 520942 666334
rect 521026 666098 521262 666334
rect 520706 665778 520942 666014
rect 521026 665778 521262 666014
rect 524426 709402 524662 709638
rect 524746 709402 524982 709638
rect 524426 709082 524662 709318
rect 524746 709082 524982 709318
rect 524426 669818 524662 670054
rect 524746 669818 524982 670054
rect 524426 669498 524662 669734
rect 524746 669498 524982 669734
rect 528146 710362 528382 710598
rect 528466 710362 528702 710598
rect 528146 710042 528382 710278
rect 528466 710042 528702 710278
rect 528146 673538 528382 673774
rect 528466 673538 528702 673774
rect 528146 673218 528382 673454
rect 528466 673218 528702 673454
rect 531866 711322 532102 711558
rect 532186 711322 532422 711558
rect 531866 711002 532102 711238
rect 532186 711002 532422 711238
rect 531866 677258 532102 677494
rect 532186 677258 532422 677494
rect 531866 676938 532102 677174
rect 532186 676938 532422 677174
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 494250 651218 494486 651454
rect 494250 650898 494486 651134
rect 524970 651218 525206 651454
rect 524970 650898 525206 651134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 492146 637538 492382 637774
rect 492466 637538 492702 637774
rect 492146 637218 492382 637454
rect 492466 637218 492702 637454
rect 509610 618938 509846 619174
rect 509610 618618 509846 618854
rect 494250 615218 494486 615454
rect 494250 614898 494486 615134
rect 524970 615218 525206 615454
rect 524970 614898 525206 615134
rect 545546 705562 545782 705798
rect 545866 705562 546102 705798
rect 545546 705242 545782 705478
rect 545866 705242 546102 705478
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 492146 601538 492382 601774
rect 492466 601538 492702 601774
rect 492146 601218 492382 601454
rect 492466 601218 492702 601454
rect 492146 565538 492382 565774
rect 492466 565538 492702 565774
rect 492146 565218 492382 565454
rect 492466 565218 492702 565454
rect 492146 529538 492382 529774
rect 492466 529538 492702 529774
rect 492146 529218 492382 529454
rect 492466 529218 492702 529454
rect 495866 569258 496102 569494
rect 496186 569258 496422 569494
rect 495866 568938 496102 569174
rect 496186 568938 496422 569174
rect 495866 533258 496102 533494
rect 496186 533258 496422 533494
rect 495866 532938 496102 533174
rect 496186 532938 496422 533174
rect 202490 510938 202726 511174
rect 202490 510618 202726 510854
rect 233210 510938 233446 511174
rect 233210 510618 233446 510854
rect 263930 510938 264166 511174
rect 263930 510618 264166 510854
rect 294650 510938 294886 511174
rect 294650 510618 294886 510854
rect 325370 510938 325606 511174
rect 325370 510618 325606 510854
rect 356090 510938 356326 511174
rect 356090 510618 356326 510854
rect 386810 510938 387046 511174
rect 386810 510618 387046 510854
rect 417530 510938 417766 511174
rect 417530 510618 417766 510854
rect 448250 510938 448486 511174
rect 448250 510618 448486 510854
rect 478970 510938 479206 511174
rect 478970 510618 479206 510854
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 310010 507218 310246 507454
rect 310010 506898 310246 507134
rect 340730 507218 340966 507454
rect 340730 506898 340966 507134
rect 371450 507218 371686 507454
rect 371450 506898 371686 507134
rect 402170 507218 402406 507454
rect 402170 506898 402406 507134
rect 432890 507218 433126 507454
rect 432890 506898 433126 507134
rect 463610 507218 463846 507454
rect 463610 506898 463846 507134
rect 494330 507218 494566 507454
rect 494330 506898 494566 507134
rect 196706 486098 196942 486334
rect 197026 486098 197262 486334
rect 196706 485778 196942 486014
rect 197026 485778 197262 486014
rect 202490 474938 202726 475174
rect 202490 474618 202726 474854
rect 233210 474938 233446 475174
rect 233210 474618 233446 474854
rect 263930 474938 264166 475174
rect 263930 474618 264166 474854
rect 294650 474938 294886 475174
rect 294650 474618 294886 474854
rect 325370 474938 325606 475174
rect 325370 474618 325606 474854
rect 356090 474938 356326 475174
rect 356090 474618 356326 474854
rect 386810 474938 387046 475174
rect 386810 474618 387046 474854
rect 417530 474938 417766 475174
rect 417530 474618 417766 474854
rect 448250 474938 448486 475174
rect 448250 474618 448486 474854
rect 478970 474938 479206 475174
rect 478970 474618 479206 474854
rect 217850 471218 218086 471454
rect 217850 470898 218086 471134
rect 248570 471218 248806 471454
rect 248570 470898 248806 471134
rect 279290 471218 279526 471454
rect 279290 470898 279526 471134
rect 310010 471218 310246 471454
rect 310010 470898 310246 471134
rect 340730 471218 340966 471454
rect 340730 470898 340966 471134
rect 371450 471218 371686 471454
rect 371450 470898 371686 471134
rect 402170 471218 402406 471454
rect 402170 470898 402406 471134
rect 432890 471218 433126 471454
rect 432890 470898 433126 471134
rect 463610 471218 463846 471454
rect 463610 470898 463846 471134
rect 494330 471218 494566 471454
rect 494330 470898 494566 471134
rect 196706 450098 196942 450334
rect 197026 450098 197262 450334
rect 196706 449778 196942 450014
rect 197026 449778 197262 450014
rect 202490 438938 202726 439174
rect 202490 438618 202726 438854
rect 233210 438938 233446 439174
rect 233210 438618 233446 438854
rect 263930 438938 264166 439174
rect 263930 438618 264166 438854
rect 294650 438938 294886 439174
rect 294650 438618 294886 438854
rect 325370 438938 325606 439174
rect 325370 438618 325606 438854
rect 356090 438938 356326 439174
rect 356090 438618 356326 438854
rect 386810 438938 387046 439174
rect 386810 438618 387046 438854
rect 417530 438938 417766 439174
rect 417530 438618 417766 438854
rect 448250 438938 448486 439174
rect 448250 438618 448486 438854
rect 478970 438938 479206 439174
rect 478970 438618 479206 438854
rect 217850 435218 218086 435454
rect 217850 434898 218086 435134
rect 248570 435218 248806 435454
rect 248570 434898 248806 435134
rect 279290 435218 279526 435454
rect 279290 434898 279526 435134
rect 310010 435218 310246 435454
rect 310010 434898 310246 435134
rect 340730 435218 340966 435454
rect 340730 434898 340966 435134
rect 371450 435218 371686 435454
rect 371450 434898 371686 435134
rect 402170 435218 402406 435454
rect 402170 434898 402406 435134
rect 432890 435218 433126 435454
rect 432890 434898 433126 435134
rect 463610 435218 463846 435454
rect 463610 434898 463846 435134
rect 494330 435218 494566 435454
rect 494330 434898 494566 435134
rect 196706 414098 196942 414334
rect 197026 414098 197262 414334
rect 196706 413778 196942 414014
rect 197026 413778 197262 414014
rect 202490 402938 202726 403174
rect 202490 402618 202726 402854
rect 233210 402938 233446 403174
rect 233210 402618 233446 402854
rect 263930 402938 264166 403174
rect 263930 402618 264166 402854
rect 294650 402938 294886 403174
rect 294650 402618 294886 402854
rect 325370 402938 325606 403174
rect 325370 402618 325606 402854
rect 356090 402938 356326 403174
rect 356090 402618 356326 402854
rect 386810 402938 387046 403174
rect 386810 402618 387046 402854
rect 417530 402938 417766 403174
rect 417530 402618 417766 402854
rect 448250 402938 448486 403174
rect 448250 402618 448486 402854
rect 478970 402938 479206 403174
rect 478970 402618 479206 402854
rect 217850 399218 218086 399454
rect 217850 398898 218086 399134
rect 248570 399218 248806 399454
rect 248570 398898 248806 399134
rect 279290 399218 279526 399454
rect 279290 398898 279526 399134
rect 310010 399218 310246 399454
rect 310010 398898 310246 399134
rect 340730 399218 340966 399454
rect 340730 398898 340966 399134
rect 371450 399218 371686 399454
rect 371450 398898 371686 399134
rect 402170 399218 402406 399454
rect 402170 398898 402406 399134
rect 432890 399218 433126 399454
rect 432890 398898 433126 399134
rect 463610 399218 463846 399454
rect 463610 398898 463846 399134
rect 494330 399218 494566 399454
rect 494330 398898 494566 399134
rect 196706 378098 196942 378334
rect 197026 378098 197262 378334
rect 196706 377778 196942 378014
rect 197026 377778 197262 378014
rect 196706 342098 196942 342334
rect 197026 342098 197262 342334
rect 196706 341778 196942 342014
rect 197026 341778 197262 342014
rect 196706 306098 196942 306334
rect 197026 306098 197262 306334
rect 196706 305778 196942 306014
rect 197026 305778 197262 306014
rect 196706 270098 196942 270334
rect 197026 270098 197262 270334
rect 196706 269778 196942 270014
rect 197026 269778 197262 270014
rect 200426 381818 200662 382054
rect 200746 381818 200982 382054
rect 200426 381498 200662 381734
rect 200746 381498 200982 381734
rect 200426 345818 200662 346054
rect 200746 345818 200982 346054
rect 200426 345498 200662 345734
rect 200746 345498 200982 345734
rect 200426 309818 200662 310054
rect 200746 309818 200982 310054
rect 200426 309498 200662 309734
rect 200746 309498 200982 309734
rect 200426 273818 200662 274054
rect 200746 273818 200982 274054
rect 200426 273498 200662 273734
rect 200746 273498 200982 273734
rect 196706 234098 196942 234334
rect 197026 234098 197262 234334
rect 196706 233778 196942 234014
rect 197026 233778 197262 234014
rect 196706 198098 196942 198334
rect 197026 198098 197262 198334
rect 196706 197778 196942 198014
rect 197026 197778 197262 198014
rect 200426 237818 200662 238054
rect 200746 237818 200982 238054
rect 200426 237498 200662 237734
rect 200746 237498 200982 237734
rect 200426 201818 200662 202054
rect 200746 201818 200982 202054
rect 200426 201498 200662 201734
rect 200746 201498 200982 201734
rect 196706 162098 196942 162334
rect 197026 162098 197262 162334
rect 196706 161778 196942 162014
rect 197026 161778 197262 162014
rect 196706 126098 196942 126334
rect 197026 126098 197262 126334
rect 196706 125778 196942 126014
rect 197026 125778 197262 126014
rect 196706 90098 196942 90334
rect 197026 90098 197262 90334
rect 196706 89778 196942 90014
rect 197026 89778 197262 90014
rect 196706 54098 196942 54334
rect 197026 54098 197262 54334
rect 196706 53778 196942 54014
rect 197026 53778 197262 54014
rect 196706 18098 196942 18334
rect 197026 18098 197262 18334
rect 196706 17778 196942 18014
rect 197026 17778 197262 18014
rect 196706 -4422 196942 -4186
rect 197026 -4422 197262 -4186
rect 196706 -4742 196942 -4506
rect 197026 -4742 197262 -4506
rect 200426 165818 200662 166054
rect 200746 165818 200982 166054
rect 200426 165498 200662 165734
rect 200746 165498 200982 165734
rect 200426 129818 200662 130054
rect 200746 129818 200982 130054
rect 200426 129498 200662 129734
rect 200746 129498 200982 129734
rect 200426 93818 200662 94054
rect 200746 93818 200982 94054
rect 200426 93498 200662 93734
rect 200746 93498 200982 93734
rect 200426 57818 200662 58054
rect 200746 57818 200982 58054
rect 200426 57498 200662 57734
rect 200746 57498 200982 57734
rect 200426 21818 200662 22054
rect 200746 21818 200982 22054
rect 200426 21498 200662 21734
rect 200746 21498 200982 21734
rect 200426 -5382 200662 -5146
rect 200746 -5382 200982 -5146
rect 200426 -5702 200662 -5466
rect 200746 -5702 200982 -5466
rect 204146 385538 204382 385774
rect 204466 385538 204702 385774
rect 204146 385218 204382 385454
rect 204466 385218 204702 385454
rect 204146 349538 204382 349774
rect 204466 349538 204702 349774
rect 204146 349218 204382 349454
rect 204466 349218 204702 349454
rect 204146 313538 204382 313774
rect 204466 313538 204702 313774
rect 204146 313218 204382 313454
rect 204466 313218 204702 313454
rect 204146 277538 204382 277774
rect 204466 277538 204702 277774
rect 204146 277218 204382 277454
rect 204466 277218 204702 277454
rect 204146 241538 204382 241774
rect 204466 241538 204702 241774
rect 204146 241218 204382 241454
rect 204466 241218 204702 241454
rect 204146 205538 204382 205774
rect 204466 205538 204702 205774
rect 204146 205218 204382 205454
rect 204466 205218 204702 205454
rect 204146 169538 204382 169774
rect 204466 169538 204702 169774
rect 204146 169218 204382 169454
rect 204466 169218 204702 169454
rect 204146 133538 204382 133774
rect 204466 133538 204702 133774
rect 204146 133218 204382 133454
rect 204466 133218 204702 133454
rect 204146 97538 204382 97774
rect 204466 97538 204702 97774
rect 204146 97218 204382 97454
rect 204466 97218 204702 97454
rect 204146 61538 204382 61774
rect 204466 61538 204702 61774
rect 204146 61218 204382 61454
rect 204466 61218 204702 61454
rect 204146 25538 204382 25774
rect 204466 25538 204702 25774
rect 204146 25218 204382 25454
rect 204466 25218 204702 25454
rect 204146 -6342 204382 -6106
rect 204466 -6342 204702 -6106
rect 204146 -6662 204382 -6426
rect 204466 -6662 204702 -6426
rect 207866 353258 208102 353494
rect 208186 353258 208422 353494
rect 207866 352938 208102 353174
rect 208186 352938 208422 353174
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 207866 317258 208102 317494
rect 208186 317258 208422 317494
rect 207866 316938 208102 317174
rect 208186 316938 208422 317174
rect 207866 281258 208102 281494
rect 208186 281258 208422 281494
rect 207866 280938 208102 281174
rect 208186 280938 208422 281174
rect 207866 245258 208102 245494
rect 208186 245258 208422 245494
rect 207866 244938 208102 245174
rect 208186 244938 208422 245174
rect 207866 209258 208102 209494
rect 208186 209258 208422 209494
rect 207866 208938 208102 209174
rect 208186 208938 208422 209174
rect 207866 173258 208102 173494
rect 208186 173258 208422 173494
rect 207866 172938 208102 173174
rect 208186 172938 208422 173174
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 207866 137258 208102 137494
rect 208186 137258 208422 137494
rect 207866 136938 208102 137174
rect 208186 136938 208422 137174
rect 207866 101258 208102 101494
rect 208186 101258 208422 101494
rect 207866 100938 208102 101174
rect 208186 100938 208422 101174
rect 207866 65258 208102 65494
rect 208186 65258 208422 65494
rect 207866 64938 208102 65174
rect 208186 64938 208422 65174
rect 207866 29258 208102 29494
rect 208186 29258 208422 29494
rect 207866 28938 208102 29174
rect 208186 28938 208422 29174
rect 207866 -7302 208102 -7066
rect 208186 -7302 208422 -7066
rect 207866 -7622 208102 -7386
rect 208186 -7622 208422 -7386
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 217826 111218 218062 111454
rect 218146 111218 218382 111454
rect 217826 110898 218062 111134
rect 218146 110898 218382 111134
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 221546 114938 221782 115174
rect 221866 114938 222102 115174
rect 221546 114618 221782 114854
rect 221866 114618 222102 114854
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -1542 221782 -1306
rect 221866 -1542 222102 -1306
rect 221546 -1862 221782 -1626
rect 221866 -1862 222102 -1626
rect 232706 378098 232942 378334
rect 233026 378098 233262 378334
rect 232706 377778 232942 378014
rect 233026 377778 233262 378014
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 225266 118658 225502 118894
rect 225586 118658 225822 118894
rect 225266 118338 225502 118574
rect 225586 118338 225822 118574
rect 236426 381818 236662 382054
rect 236746 381818 236982 382054
rect 236426 381498 236662 381734
rect 236746 381498 236982 381734
rect 232706 342098 232942 342334
rect 233026 342098 233262 342334
rect 232706 341778 232942 342014
rect 233026 341778 233262 342014
rect 232706 306098 232942 306334
rect 233026 306098 233262 306334
rect 232706 305778 232942 306014
rect 233026 305778 233262 306014
rect 232706 270098 232942 270334
rect 233026 270098 233262 270334
rect 232706 269778 232942 270014
rect 233026 269778 233262 270014
rect 232706 234098 232942 234334
rect 233026 234098 233262 234334
rect 232706 233778 232942 234014
rect 233026 233778 233262 234014
rect 232706 198098 232942 198334
rect 233026 198098 233262 198334
rect 232706 197778 232942 198014
rect 233026 197778 233262 198014
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -2502 225502 -2266
rect 225586 -2502 225822 -2266
rect 225266 -2822 225502 -2586
rect 225586 -2822 225822 -2586
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 232706 162098 232942 162334
rect 233026 162098 233262 162334
rect 232706 161778 232942 162014
rect 233026 161778 233262 162014
rect 240146 385538 240382 385774
rect 240466 385538 240702 385774
rect 240146 385218 240382 385454
rect 240466 385218 240702 385454
rect 236426 345818 236662 346054
rect 236746 345818 236982 346054
rect 236426 345498 236662 345734
rect 236746 345498 236982 345734
rect 236426 309818 236662 310054
rect 236746 309818 236982 310054
rect 236426 309498 236662 309734
rect 236746 309498 236982 309734
rect 236426 273818 236662 274054
rect 236746 273818 236982 274054
rect 236426 273498 236662 273734
rect 236746 273498 236982 273734
rect 236426 237818 236662 238054
rect 236746 237818 236982 238054
rect 236426 237498 236662 237734
rect 236746 237498 236982 237734
rect 236426 201818 236662 202054
rect 236746 201818 236982 202054
rect 236426 201498 236662 201734
rect 236746 201498 236982 201734
rect 236426 165818 236662 166054
rect 236746 165818 236982 166054
rect 236426 165498 236662 165734
rect 236746 165498 236982 165734
rect 232706 126098 232942 126334
rect 233026 126098 233262 126334
rect 232706 125778 232942 126014
rect 233026 125778 233262 126014
rect 232706 90098 232942 90334
rect 233026 90098 233262 90334
rect 232706 89778 232942 90014
rect 233026 89778 233262 90014
rect 232706 54098 232942 54334
rect 233026 54098 233262 54334
rect 232706 53778 232942 54014
rect 233026 53778 233262 54014
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 228986 -3462 229222 -3226
rect 229306 -3462 229542 -3226
rect 228986 -3782 229222 -3546
rect 229306 -3782 229542 -3546
rect 232706 18098 232942 18334
rect 233026 18098 233262 18334
rect 232706 17778 232942 18014
rect 233026 17778 233262 18014
rect 236426 129818 236662 130054
rect 236746 129818 236982 130054
rect 236426 129498 236662 129734
rect 236746 129498 236982 129734
rect 240146 349538 240382 349774
rect 240466 349538 240702 349774
rect 240146 349218 240382 349454
rect 240466 349218 240702 349454
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 268706 378098 268942 378334
rect 269026 378098 269262 378334
rect 268706 377778 268942 378014
rect 269026 377778 269262 378014
rect 268706 342098 268942 342334
rect 269026 342098 269262 342334
rect 268706 341778 268942 342014
rect 269026 341778 269262 342014
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 272426 381818 272662 382054
rect 272746 381818 272982 382054
rect 272426 381498 272662 381734
rect 272746 381498 272982 381734
rect 272426 345818 272662 346054
rect 272746 345818 272982 346054
rect 272426 345498 272662 345734
rect 272746 345498 272982 345734
rect 276146 385538 276382 385774
rect 276466 385538 276702 385774
rect 276146 385218 276382 385454
rect 276466 385218 276702 385454
rect 276146 349538 276382 349774
rect 276466 349538 276702 349774
rect 276146 349218 276382 349454
rect 276466 349218 276702 349454
rect 259610 330938 259846 331174
rect 259610 330618 259846 330854
rect 244250 327218 244486 327454
rect 244250 326898 244486 327134
rect 274970 327218 275206 327454
rect 274970 326898 275206 327134
rect 259610 294938 259846 295174
rect 259610 294618 259846 294854
rect 244250 291218 244486 291454
rect 244250 290898 244486 291134
rect 274970 291218 275206 291454
rect 274970 290898 275206 291134
rect 259610 258938 259846 259174
rect 259610 258618 259846 258854
rect 244250 255218 244486 255454
rect 244250 254898 244486 255134
rect 274970 255218 275206 255454
rect 274970 254898 275206 255134
rect 259610 222938 259846 223174
rect 259610 222618 259846 222854
rect 244250 219218 244486 219454
rect 244250 218898 244486 219134
rect 274970 219218 275206 219454
rect 274970 218898 275206 219134
rect 259610 186938 259846 187174
rect 259610 186618 259846 186854
rect 244250 183218 244486 183454
rect 244250 182898 244486 183134
rect 274970 183218 275206 183454
rect 274970 182898 275206 183134
rect 259610 150938 259846 151174
rect 259610 150618 259846 150854
rect 244250 147218 244486 147454
rect 244250 146898 244486 147134
rect 274970 147218 275206 147454
rect 274970 146898 275206 147134
rect 236426 93818 236662 94054
rect 236746 93818 236982 94054
rect 236426 93498 236662 93734
rect 236746 93498 236982 93734
rect 236426 57818 236662 58054
rect 236746 57818 236982 58054
rect 236426 57498 236662 57734
rect 236746 57498 236982 57734
rect 240146 97538 240382 97774
rect 240466 97538 240702 97774
rect 240146 97218 240382 97454
rect 240466 97218 240702 97454
rect 240146 61538 240382 61774
rect 240466 61538 240702 61774
rect 240146 61218 240382 61454
rect 240466 61218 240702 61454
rect 236426 21818 236662 22054
rect 236746 21818 236982 22054
rect 236426 21498 236662 21734
rect 236746 21498 236982 21734
rect 232706 -4422 232942 -4186
rect 233026 -4422 233262 -4186
rect 232706 -4742 232942 -4506
rect 233026 -4742 233262 -4506
rect 236426 -5382 236662 -5146
rect 236746 -5382 236982 -5146
rect 236426 -5702 236662 -5466
rect 236746 -5702 236982 -5466
rect 240146 25538 240382 25774
rect 240466 25538 240702 25774
rect 240146 25218 240382 25454
rect 240466 25218 240702 25454
rect 240146 -6342 240382 -6106
rect 240466 -6342 240702 -6106
rect 240146 -6662 240382 -6426
rect 240466 -6662 240702 -6426
rect 243866 101258 244102 101494
rect 244186 101258 244422 101494
rect 243866 100938 244102 101174
rect 244186 100938 244422 101174
rect 243866 65258 244102 65494
rect 244186 65258 244422 65494
rect 243866 64938 244102 65174
rect 244186 64938 244422 65174
rect 243866 29258 244102 29494
rect 244186 29258 244422 29494
rect 243866 28938 244102 29174
rect 244186 28938 244422 29174
rect 243866 -7302 244102 -7066
rect 244186 -7302 244422 -7066
rect 243866 -7622 244102 -7386
rect 244186 -7622 244422 -7386
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -1542 257782 -1306
rect 257866 -1542 258102 -1306
rect 257546 -1862 257782 -1626
rect 257866 -1862 258102 -1626
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -2502 261502 -2266
rect 261586 -2502 261822 -2266
rect 261266 -2822 261502 -2586
rect 261586 -2822 261822 -2586
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 264986 -3462 265222 -3226
rect 265306 -3462 265542 -3226
rect 264986 -3782 265222 -3546
rect 265306 -3782 265542 -3546
rect 268706 126098 268942 126334
rect 269026 126098 269262 126334
rect 268706 125778 268942 126014
rect 269026 125778 269262 126014
rect 268706 90098 268942 90334
rect 269026 90098 269262 90334
rect 268706 89778 268942 90014
rect 269026 89778 269262 90014
rect 268706 54098 268942 54334
rect 269026 54098 269262 54334
rect 268706 53778 268942 54014
rect 269026 53778 269262 54014
rect 268706 18098 268942 18334
rect 269026 18098 269262 18334
rect 268706 17778 268942 18014
rect 269026 17778 269262 18014
rect 268706 -4422 268942 -4186
rect 269026 -4422 269262 -4186
rect 268706 -4742 268942 -4506
rect 269026 -4742 269262 -4506
rect 272426 129818 272662 130054
rect 272746 129818 272982 130054
rect 272426 129498 272662 129734
rect 272746 129498 272982 129734
rect 272426 93818 272662 94054
rect 272746 93818 272982 94054
rect 272426 93498 272662 93734
rect 272746 93498 272982 93734
rect 272426 57818 272662 58054
rect 272746 57818 272982 58054
rect 272426 57498 272662 57734
rect 272746 57498 272982 57734
rect 272426 21818 272662 22054
rect 272746 21818 272982 22054
rect 272426 21498 272662 21734
rect 272746 21498 272982 21734
rect 272426 -5382 272662 -5146
rect 272746 -5382 272982 -5146
rect 272426 -5702 272662 -5466
rect 272746 -5702 272982 -5466
rect 276146 97538 276382 97774
rect 276466 97538 276702 97774
rect 276146 97218 276382 97454
rect 276466 97218 276702 97454
rect 279866 101258 280102 101494
rect 280186 101258 280422 101494
rect 279866 100938 280102 101174
rect 280186 100938 280422 101174
rect 276146 61538 276382 61774
rect 276466 61538 276702 61774
rect 276146 61218 276382 61454
rect 276466 61218 276702 61454
rect 276146 25538 276382 25774
rect 276466 25538 276702 25774
rect 276146 25218 276382 25454
rect 276466 25218 276702 25454
rect 276146 -6342 276382 -6106
rect 276466 -6342 276702 -6106
rect 276146 -6662 276382 -6426
rect 276466 -6662 276702 -6426
rect 279866 65258 280102 65494
rect 280186 65258 280422 65494
rect 279866 64938 280102 65174
rect 280186 64938 280422 65174
rect 279866 29258 280102 29494
rect 280186 29258 280422 29494
rect 279866 28938 280102 29174
rect 280186 28938 280422 29174
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 279866 -7302 280102 -7066
rect 280186 -7302 280422 -7066
rect 279866 -7622 280102 -7386
rect 280186 -7622 280422 -7386
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 304706 378098 304942 378334
rect 305026 378098 305262 378334
rect 304706 377778 304942 378014
rect 305026 377778 305262 378014
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 308426 381818 308662 382054
rect 308746 381818 308982 382054
rect 308426 381498 308662 381734
rect 308746 381498 308982 381734
rect 308426 345818 308662 346054
rect 308746 345818 308982 346054
rect 308426 345498 308662 345734
rect 308746 345498 308982 345734
rect 304706 342098 304942 342334
rect 305026 342098 305262 342334
rect 304706 341778 304942 342014
rect 305026 341778 305262 342014
rect 304706 306098 304942 306334
rect 305026 306098 305262 306334
rect 304706 305778 304942 306014
rect 305026 305778 305262 306014
rect 304706 270098 304942 270334
rect 305026 270098 305262 270334
rect 304706 269778 304942 270014
rect 305026 269778 305262 270014
rect 304706 234098 304942 234334
rect 305026 234098 305262 234334
rect 304706 233778 304942 234014
rect 305026 233778 305262 234014
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -1542 293782 -1306
rect 293866 -1542 294102 -1306
rect 293546 -1862 293782 -1626
rect 293866 -1862 294102 -1626
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 308426 309818 308662 310054
rect 308746 309818 308982 310054
rect 308426 309498 308662 309734
rect 308746 309498 308982 309734
rect 308426 273818 308662 274054
rect 308746 273818 308982 274054
rect 308426 273498 308662 273734
rect 308746 273498 308982 273734
rect 308426 237818 308662 238054
rect 308746 237818 308982 238054
rect 308426 237498 308662 237734
rect 308746 237498 308982 237734
rect 304706 198098 304942 198334
rect 305026 198098 305262 198334
rect 304706 197778 304942 198014
rect 305026 197778 305262 198014
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 308426 201818 308662 202054
rect 308746 201818 308982 202054
rect 308426 201498 308662 201734
rect 308746 201498 308982 201734
rect 304706 162098 304942 162334
rect 305026 162098 305262 162334
rect 304706 161778 304942 162014
rect 305026 161778 305262 162014
rect 304706 126098 304942 126334
rect 305026 126098 305262 126334
rect 304706 125778 304942 126014
rect 305026 125778 305262 126014
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -2502 297502 -2266
rect 297586 -2502 297822 -2266
rect 297266 -2822 297502 -2586
rect 297586 -2822 297822 -2586
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 300986 -3462 301222 -3226
rect 301306 -3462 301542 -3226
rect 300986 -3782 301222 -3546
rect 301306 -3782 301542 -3546
rect 304706 90098 304942 90334
rect 305026 90098 305262 90334
rect 304706 89778 304942 90014
rect 305026 89778 305262 90014
rect 312146 385538 312382 385774
rect 312466 385538 312702 385774
rect 312146 385218 312382 385454
rect 312466 385218 312702 385454
rect 312146 349538 312382 349774
rect 312466 349538 312702 349774
rect 312146 349218 312382 349454
rect 312466 349218 312702 349454
rect 312146 313538 312382 313774
rect 312466 313538 312702 313774
rect 312146 313218 312382 313454
rect 312466 313218 312702 313454
rect 312146 277538 312382 277774
rect 312466 277538 312702 277774
rect 312146 277218 312382 277454
rect 312466 277218 312702 277454
rect 312146 241538 312382 241774
rect 312466 241538 312702 241774
rect 312146 241218 312382 241454
rect 312466 241218 312702 241454
rect 312146 205538 312382 205774
rect 312466 205538 312702 205774
rect 312146 205218 312382 205454
rect 312466 205218 312702 205454
rect 308426 165818 308662 166054
rect 308746 165818 308982 166054
rect 308426 165498 308662 165734
rect 308746 165498 308982 165734
rect 308426 129818 308662 130054
rect 308746 129818 308982 130054
rect 308426 129498 308662 129734
rect 308746 129498 308982 129734
rect 315866 353258 316102 353494
rect 316186 353258 316422 353494
rect 315866 352938 316102 353174
rect 316186 352938 316422 353174
rect 315866 317258 316102 317494
rect 316186 317258 316422 317494
rect 315866 316938 316102 317174
rect 316186 316938 316422 317174
rect 315866 281258 316102 281494
rect 316186 281258 316422 281494
rect 315866 280938 316102 281174
rect 316186 280938 316422 281174
rect 315866 245258 316102 245494
rect 316186 245258 316422 245494
rect 315866 244938 316102 245174
rect 316186 244938 316422 245174
rect 315866 209258 316102 209494
rect 316186 209258 316422 209494
rect 315866 208938 316102 209174
rect 316186 208938 316422 209174
rect 312146 169538 312382 169774
rect 312466 169538 312702 169774
rect 312146 169218 312382 169454
rect 312466 169218 312702 169454
rect 312146 133538 312382 133774
rect 312466 133538 312702 133774
rect 312146 133218 312382 133454
rect 312466 133218 312702 133454
rect 308426 93818 308662 94054
rect 308746 93818 308982 94054
rect 308426 93498 308662 93734
rect 308746 93498 308982 93734
rect 304706 54098 304942 54334
rect 305026 54098 305262 54334
rect 304706 53778 304942 54014
rect 305026 53778 305262 54014
rect 304706 18098 304942 18334
rect 305026 18098 305262 18334
rect 304706 17778 304942 18014
rect 305026 17778 305262 18014
rect 304706 -4422 304942 -4186
rect 305026 -4422 305262 -4186
rect 304706 -4742 304942 -4506
rect 305026 -4742 305262 -4506
rect 308426 57818 308662 58054
rect 308746 57818 308982 58054
rect 308426 57498 308662 57734
rect 308746 57498 308982 57734
rect 308426 21818 308662 22054
rect 308746 21818 308982 22054
rect 308426 21498 308662 21734
rect 308746 21498 308982 21734
rect 308426 -5382 308662 -5146
rect 308746 -5382 308982 -5146
rect 308426 -5702 308662 -5466
rect 308746 -5702 308982 -5466
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 315866 173258 316102 173494
rect 316186 173258 316422 173494
rect 315866 172938 316102 173174
rect 316186 172938 316422 173174
rect 315866 137258 316102 137494
rect 316186 137258 316422 137494
rect 315866 136938 316102 137174
rect 316186 136938 316422 137174
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 315866 101258 316102 101494
rect 316186 101258 316422 101494
rect 315866 100938 316102 101174
rect 316186 100938 316422 101174
rect 312146 97538 312382 97774
rect 312466 97538 312702 97774
rect 312146 97218 312382 97454
rect 312466 97218 312702 97454
rect 312146 61538 312382 61774
rect 312466 61538 312702 61774
rect 312146 61218 312382 61454
rect 312466 61218 312702 61454
rect 312146 25538 312382 25774
rect 312466 25538 312702 25774
rect 312146 25218 312382 25454
rect 312466 25218 312702 25454
rect 312146 -6342 312382 -6106
rect 312466 -6342 312702 -6106
rect 312146 -6662 312382 -6426
rect 312466 -6662 312702 -6426
rect 315866 65258 316102 65494
rect 316186 65258 316422 65494
rect 315866 64938 316102 65174
rect 316186 64938 316422 65174
rect 315866 29258 316102 29494
rect 316186 29258 316422 29494
rect 315866 28938 316102 29174
rect 316186 28938 316422 29174
rect 315866 -7302 316102 -7066
rect 316186 -7302 316422 -7066
rect 315866 -7622 316102 -7386
rect 316186 -7622 316422 -7386
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -1542 329782 -1306
rect 329866 -1542 330102 -1306
rect 329546 -1862 329782 -1626
rect 329866 -1862 330102 -1626
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 340706 378098 340942 378334
rect 341026 378098 341262 378334
rect 340706 377778 340942 378014
rect 341026 377778 341262 378014
rect 340706 342098 340942 342334
rect 341026 342098 341262 342334
rect 340706 341778 340942 342014
rect 341026 341778 341262 342014
rect 340706 306098 340942 306334
rect 341026 306098 341262 306334
rect 340706 305778 340942 306014
rect 341026 305778 341262 306014
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 340706 270098 340942 270334
rect 341026 270098 341262 270334
rect 340706 269778 340942 270014
rect 341026 269778 341262 270014
rect 340706 234098 340942 234334
rect 341026 234098 341262 234334
rect 340706 233778 340942 234014
rect 341026 233778 341262 234014
rect 340706 198098 340942 198334
rect 341026 198098 341262 198334
rect 340706 197778 340942 198014
rect 341026 197778 341262 198014
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -2502 333502 -2266
rect 333586 -2502 333822 -2266
rect 333266 -2822 333502 -2586
rect 333586 -2822 333822 -2586
rect 344426 381818 344662 382054
rect 344746 381818 344982 382054
rect 344426 381498 344662 381734
rect 344746 381498 344982 381734
rect 344426 345818 344662 346054
rect 344746 345818 344982 346054
rect 344426 345498 344662 345734
rect 344746 345498 344982 345734
rect 344426 309818 344662 310054
rect 344746 309818 344982 310054
rect 344426 309498 344662 309734
rect 344746 309498 344982 309734
rect 344426 273818 344662 274054
rect 344746 273818 344982 274054
rect 344426 273498 344662 273734
rect 344746 273498 344982 273734
rect 348146 385538 348382 385774
rect 348466 385538 348702 385774
rect 348146 385218 348382 385454
rect 348466 385218 348702 385454
rect 348146 349538 348382 349774
rect 348466 349538 348702 349774
rect 348146 349218 348382 349454
rect 348466 349218 348702 349454
rect 348146 313538 348382 313774
rect 348466 313538 348702 313774
rect 348146 313218 348382 313454
rect 348466 313218 348702 313454
rect 348146 277538 348382 277774
rect 348466 277538 348702 277774
rect 348146 277218 348382 277454
rect 348466 277218 348702 277454
rect 344426 237818 344662 238054
rect 344746 237818 344982 238054
rect 344426 237498 344662 237734
rect 344746 237498 344982 237734
rect 344426 201818 344662 202054
rect 344746 201818 344982 202054
rect 344426 201498 344662 201734
rect 344746 201498 344982 201734
rect 340706 162098 340942 162334
rect 341026 162098 341262 162334
rect 340706 161778 340942 162014
rect 341026 161778 341262 162014
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 336986 -3462 337222 -3226
rect 337306 -3462 337542 -3226
rect 336986 -3782 337222 -3546
rect 337306 -3782 337542 -3546
rect 351866 353258 352102 353494
rect 352186 353258 352422 353494
rect 351866 352938 352102 353174
rect 352186 352938 352422 353174
rect 351866 317258 352102 317494
rect 352186 317258 352422 317494
rect 351866 316938 352102 317174
rect 352186 316938 352422 317174
rect 351866 281258 352102 281494
rect 352186 281258 352422 281494
rect 351866 280938 352102 281174
rect 352186 280938 352422 281174
rect 348146 241538 348382 241774
rect 348466 241538 348702 241774
rect 348146 241218 348382 241454
rect 348466 241218 348702 241454
rect 348146 205538 348382 205774
rect 348466 205538 348702 205774
rect 348146 205218 348382 205454
rect 348466 205218 348702 205454
rect 344426 165818 344662 166054
rect 344746 165818 344982 166054
rect 344426 165498 344662 165734
rect 344746 165498 344982 165734
rect 351866 245258 352102 245494
rect 352186 245258 352422 245494
rect 351866 244938 352102 245174
rect 352186 244938 352422 245174
rect 351866 209258 352102 209494
rect 352186 209258 352422 209494
rect 351866 208938 352102 209174
rect 352186 208938 352422 209174
rect 348146 169538 348382 169774
rect 348466 169538 348702 169774
rect 348146 169218 348382 169454
rect 348466 169218 348702 169454
rect 344426 129818 344662 130054
rect 344746 129818 344982 130054
rect 344426 129498 344662 129734
rect 344746 129498 344982 129734
rect 340706 126098 340942 126334
rect 341026 126098 341262 126334
rect 340706 125778 340942 126014
rect 341026 125778 341262 126014
rect 340706 90098 340942 90334
rect 341026 90098 341262 90334
rect 340706 89778 340942 90014
rect 341026 89778 341262 90014
rect 340706 54098 340942 54334
rect 341026 54098 341262 54334
rect 340706 53778 340942 54014
rect 341026 53778 341262 54014
rect 340706 18098 340942 18334
rect 341026 18098 341262 18334
rect 340706 17778 340942 18014
rect 341026 17778 341262 18014
rect 340706 -4422 340942 -4186
rect 341026 -4422 341262 -4186
rect 340706 -4742 340942 -4506
rect 341026 -4742 341262 -4506
rect 344426 93818 344662 94054
rect 344746 93818 344982 94054
rect 344426 93498 344662 93734
rect 344746 93498 344982 93734
rect 344426 57818 344662 58054
rect 344746 57818 344982 58054
rect 344426 57498 344662 57734
rect 344746 57498 344982 57734
rect 344426 21818 344662 22054
rect 344746 21818 344982 22054
rect 344426 21498 344662 21734
rect 344746 21498 344982 21734
rect 344426 -5382 344662 -5146
rect 344746 -5382 344982 -5146
rect 344426 -5702 344662 -5466
rect 344746 -5702 344982 -5466
rect 348146 133538 348382 133774
rect 348466 133538 348702 133774
rect 348146 133218 348382 133454
rect 348466 133218 348702 133454
rect 351866 173258 352102 173494
rect 352186 173258 352422 173494
rect 351866 172938 352102 173174
rect 352186 172938 352422 173174
rect 351866 137258 352102 137494
rect 352186 137258 352422 137494
rect 351866 136938 352102 137174
rect 352186 136938 352422 137174
rect 348146 97538 348382 97774
rect 348466 97538 348702 97774
rect 348146 97218 348382 97454
rect 348466 97218 348702 97454
rect 348146 61538 348382 61774
rect 348466 61538 348702 61774
rect 348146 61218 348382 61454
rect 348466 61218 348702 61454
rect 348146 25538 348382 25774
rect 348466 25538 348702 25774
rect 348146 25218 348382 25454
rect 348466 25218 348702 25454
rect 348146 -6342 348382 -6106
rect 348466 -6342 348702 -6106
rect 348146 -6662 348382 -6426
rect 348466 -6662 348702 -6426
rect 384146 385538 384382 385774
rect 384466 385538 384702 385774
rect 384146 385218 384382 385454
rect 384466 385218 384702 385454
rect 384146 349538 384382 349774
rect 384466 349538 384702 349774
rect 384146 349218 384382 349454
rect 384466 349218 384702 349454
rect 420146 385538 420382 385774
rect 420466 385538 420702 385774
rect 420146 385218 420382 385454
rect 420466 385218 420702 385454
rect 420146 349538 420382 349774
rect 420466 349538 420702 349774
rect 456146 385538 456382 385774
rect 456466 385538 456702 385774
rect 456146 385218 456382 385454
rect 456466 385218 456702 385454
rect 492146 385538 492382 385774
rect 492466 385538 492702 385774
rect 492146 385218 492382 385454
rect 492466 385218 492702 385454
rect 420146 349218 420382 349454
rect 420466 349218 420702 349454
rect 492146 349538 492382 349774
rect 492466 349538 492702 349774
rect 492146 349218 492382 349454
rect 492466 349218 492702 349454
rect 379610 330938 379846 331174
rect 379610 330618 379846 330854
rect 410330 330938 410566 331174
rect 410330 330618 410566 330854
rect 441050 330938 441286 331174
rect 441050 330618 441286 330854
rect 471770 330938 472006 331174
rect 471770 330618 472006 330854
rect 364250 327218 364486 327454
rect 364250 326898 364486 327134
rect 394970 327218 395206 327454
rect 394970 326898 395206 327134
rect 425690 327218 425926 327454
rect 425690 326898 425926 327134
rect 456410 327218 456646 327454
rect 456410 326898 456646 327134
rect 487130 327218 487366 327454
rect 487130 326898 487366 327134
rect 379610 294938 379846 295174
rect 379610 294618 379846 294854
rect 410330 294938 410566 295174
rect 410330 294618 410566 294854
rect 441050 294938 441286 295174
rect 441050 294618 441286 294854
rect 471770 294938 472006 295174
rect 471770 294618 472006 294854
rect 364250 291218 364486 291454
rect 364250 290898 364486 291134
rect 394970 291218 395206 291454
rect 394970 290898 395206 291134
rect 425690 291218 425926 291454
rect 425690 290898 425926 291134
rect 456410 291218 456646 291454
rect 456410 290898 456646 291134
rect 487130 291218 487366 291454
rect 487130 290898 487366 291134
rect 379610 258938 379846 259174
rect 379610 258618 379846 258854
rect 410330 258938 410566 259174
rect 410330 258618 410566 258854
rect 441050 258938 441286 259174
rect 441050 258618 441286 258854
rect 471770 258938 472006 259174
rect 471770 258618 472006 258854
rect 364250 255218 364486 255454
rect 364250 254898 364486 255134
rect 394970 255218 395206 255454
rect 394970 254898 395206 255134
rect 425690 255218 425926 255454
rect 425690 254898 425926 255134
rect 456410 255218 456646 255454
rect 456410 254898 456646 255134
rect 487130 255218 487366 255454
rect 487130 254898 487366 255134
rect 379610 222938 379846 223174
rect 379610 222618 379846 222854
rect 410330 222938 410566 223174
rect 410330 222618 410566 222854
rect 441050 222938 441286 223174
rect 441050 222618 441286 222854
rect 471770 222938 472006 223174
rect 471770 222618 472006 222854
rect 364250 219218 364486 219454
rect 364250 218898 364486 219134
rect 394970 219218 395206 219454
rect 394970 218898 395206 219134
rect 425690 219218 425926 219454
rect 425690 218898 425926 219134
rect 456410 219218 456646 219454
rect 456410 218898 456646 219134
rect 487130 219218 487366 219454
rect 487130 218898 487366 219134
rect 379610 186938 379846 187174
rect 379610 186618 379846 186854
rect 410330 186938 410566 187174
rect 410330 186618 410566 186854
rect 441050 186938 441286 187174
rect 441050 186618 441286 186854
rect 471770 186938 472006 187174
rect 471770 186618 472006 186854
rect 364250 183218 364486 183454
rect 364250 182898 364486 183134
rect 394970 183218 395206 183454
rect 394970 182898 395206 183134
rect 425690 183218 425926 183454
rect 425690 182898 425926 183134
rect 456410 183218 456646 183454
rect 456410 182898 456646 183134
rect 487130 183218 487366 183454
rect 487130 182898 487366 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 379610 114938 379846 115174
rect 379610 114618 379846 114854
rect 364250 111218 364486 111454
rect 364250 110898 364486 111134
rect 394970 111218 395206 111454
rect 394970 110898 395206 111134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 351866 101258 352102 101494
rect 352186 101258 352422 101494
rect 351866 100938 352102 101174
rect 352186 100938 352422 101174
rect 351866 65258 352102 65494
rect 352186 65258 352422 65494
rect 351866 64938 352102 65174
rect 352186 64938 352422 65174
rect 351866 29258 352102 29494
rect 352186 29258 352422 29494
rect 351866 28938 352102 29174
rect 352186 28938 352422 29174
rect 351866 -7302 352102 -7066
rect 352186 -7302 352422 -7066
rect 351866 -7622 352102 -7386
rect 352186 -7622 352422 -7386
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -1542 365782 -1306
rect 365866 -1542 366102 -1306
rect 365546 -1862 365782 -1626
rect 365866 -1862 366102 -1626
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -2502 369502 -2266
rect 369586 -2502 369822 -2266
rect 369266 -2822 369502 -2586
rect 369586 -2822 369822 -2586
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 372986 -3462 373222 -3226
rect 373306 -3462 373542 -3226
rect 372986 -3782 373222 -3546
rect 373306 -3782 373542 -3546
rect 376706 90098 376942 90334
rect 377026 90098 377262 90334
rect 376706 89778 376942 90014
rect 377026 89778 377262 90014
rect 376706 54098 376942 54334
rect 377026 54098 377262 54334
rect 376706 53778 376942 54014
rect 377026 53778 377262 54014
rect 376706 18098 376942 18334
rect 377026 18098 377262 18334
rect 376706 17778 376942 18014
rect 377026 17778 377262 18014
rect 376706 -4422 376942 -4186
rect 377026 -4422 377262 -4186
rect 376706 -4742 376942 -4506
rect 377026 -4742 377262 -4506
rect 380426 93818 380662 94054
rect 380746 93818 380982 94054
rect 380426 93498 380662 93734
rect 380746 93498 380982 93734
rect 380426 57818 380662 58054
rect 380746 57818 380982 58054
rect 380426 57498 380662 57734
rect 380746 57498 380982 57734
rect 380426 21818 380662 22054
rect 380746 21818 380982 22054
rect 380426 21498 380662 21734
rect 380746 21498 380982 21734
rect 380426 -5382 380662 -5146
rect 380746 -5382 380982 -5146
rect 380426 -5702 380662 -5466
rect 380746 -5702 380982 -5466
rect 384146 97538 384382 97774
rect 384466 97538 384702 97774
rect 384146 97218 384382 97454
rect 384466 97218 384702 97454
rect 384146 61538 384382 61774
rect 384466 61538 384702 61774
rect 384146 61218 384382 61454
rect 384466 61218 384702 61454
rect 384146 25538 384382 25774
rect 384466 25538 384702 25774
rect 384146 25218 384382 25454
rect 384466 25218 384702 25454
rect 384146 -6342 384382 -6106
rect 384466 -6342 384702 -6106
rect 384146 -6662 384382 -6426
rect 384466 -6662 384702 -6426
rect 387866 65258 388102 65494
rect 388186 65258 388422 65494
rect 387866 64938 388102 65174
rect 388186 64938 388422 65174
rect 387866 29258 388102 29494
rect 388186 29258 388422 29494
rect 387866 28938 388102 29174
rect 388186 28938 388422 29174
rect 387866 -7302 388102 -7066
rect 388186 -7302 388422 -7066
rect 387866 -7622 388102 -7386
rect 388186 -7622 388422 -7386
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -1542 401782 -1306
rect 401866 -1542 402102 -1306
rect 401546 -1862 401782 -1626
rect 401866 -1862 402102 -1626
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -2502 405502 -2266
rect 405586 -2502 405822 -2266
rect 405266 -2822 405502 -2586
rect 405586 -2822 405822 -2586
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 408986 -3462 409222 -3226
rect 409306 -3462 409542 -3226
rect 408986 -3782 409222 -3546
rect 409306 -3782 409542 -3546
rect 412706 162098 412942 162334
rect 413026 162098 413262 162334
rect 412706 161778 412942 162014
rect 413026 161778 413262 162014
rect 412706 126098 412942 126334
rect 413026 126098 413262 126334
rect 412706 125778 412942 126014
rect 413026 125778 413262 126014
rect 412706 90098 412942 90334
rect 413026 90098 413262 90334
rect 412706 89778 412942 90014
rect 413026 89778 413262 90014
rect 412706 54098 412942 54334
rect 413026 54098 413262 54334
rect 412706 53778 412942 54014
rect 413026 53778 413262 54014
rect 412706 18098 412942 18334
rect 413026 18098 413262 18334
rect 412706 17778 412942 18014
rect 413026 17778 413262 18014
rect 412706 -4422 412942 -4186
rect 413026 -4422 413262 -4186
rect 412706 -4742 412942 -4506
rect 413026 -4742 413262 -4506
rect 416426 165818 416662 166054
rect 416746 165818 416982 166054
rect 416426 165498 416662 165734
rect 416746 165498 416982 165734
rect 416426 129818 416662 130054
rect 416746 129818 416982 130054
rect 416426 129498 416662 129734
rect 416746 129498 416982 129734
rect 416426 93818 416662 94054
rect 416746 93818 416982 94054
rect 416426 93498 416662 93734
rect 416746 93498 416982 93734
rect 416426 57818 416662 58054
rect 416746 57818 416982 58054
rect 416426 57498 416662 57734
rect 416746 57498 416982 57734
rect 416426 21818 416662 22054
rect 416746 21818 416982 22054
rect 416426 21498 416662 21734
rect 416746 21498 416982 21734
rect 416426 -5382 416662 -5146
rect 416746 -5382 416982 -5146
rect 416426 -5702 416662 -5466
rect 416746 -5702 416982 -5466
rect 420146 169538 420382 169774
rect 420466 169538 420702 169774
rect 420146 169218 420382 169454
rect 420466 169218 420702 169454
rect 420146 133538 420382 133774
rect 420466 133538 420702 133774
rect 420146 133218 420382 133454
rect 420466 133218 420702 133454
rect 420146 97538 420382 97774
rect 420466 97538 420702 97774
rect 420146 97218 420382 97454
rect 420466 97218 420702 97454
rect 420146 61538 420382 61774
rect 420466 61538 420702 61774
rect 420146 61218 420382 61454
rect 420466 61218 420702 61454
rect 420146 25538 420382 25774
rect 420466 25538 420702 25774
rect 420146 25218 420382 25454
rect 420466 25218 420702 25454
rect 420146 -6342 420382 -6106
rect 420466 -6342 420702 -6106
rect 420146 -6662 420382 -6426
rect 420466 -6662 420702 -6426
rect 423866 173258 424102 173494
rect 424186 173258 424422 173494
rect 423866 172938 424102 173174
rect 424186 172938 424422 173174
rect 423866 137258 424102 137494
rect 424186 137258 424422 137494
rect 423866 136938 424102 137174
rect 424186 136938 424422 137174
rect 423866 101258 424102 101494
rect 424186 101258 424422 101494
rect 423866 100938 424102 101174
rect 424186 100938 424422 101174
rect 423866 65258 424102 65494
rect 424186 65258 424422 65494
rect 423866 64938 424102 65174
rect 424186 64938 424422 65174
rect 423866 29258 424102 29494
rect 424186 29258 424422 29494
rect 423866 28938 424102 29174
rect 424186 28938 424422 29174
rect 423866 -7302 424102 -7066
rect 424186 -7302 424422 -7066
rect 423866 -7622 424102 -7386
rect 424186 -7622 424422 -7386
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -1542 437782 -1306
rect 437866 -1542 438102 -1306
rect 437546 -1862 437782 -1626
rect 437866 -1862 438102 -1626
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -2502 441502 -2266
rect 441586 -2502 441822 -2266
rect 441266 -2822 441502 -2586
rect 441586 -2822 441822 -2586
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 444986 -3462 445222 -3226
rect 445306 -3462 445542 -3226
rect 444986 -3782 445222 -3546
rect 445306 -3782 445542 -3546
rect 448706 162098 448942 162334
rect 449026 162098 449262 162334
rect 448706 161778 448942 162014
rect 449026 161778 449262 162014
rect 448706 126098 448942 126334
rect 449026 126098 449262 126334
rect 448706 125778 448942 126014
rect 449026 125778 449262 126014
rect 448706 90098 448942 90334
rect 449026 90098 449262 90334
rect 448706 89778 448942 90014
rect 449026 89778 449262 90014
rect 448706 54098 448942 54334
rect 449026 54098 449262 54334
rect 448706 53778 448942 54014
rect 449026 53778 449262 54014
rect 448706 18098 448942 18334
rect 449026 18098 449262 18334
rect 448706 17778 448942 18014
rect 449026 17778 449262 18014
rect 448706 -4422 448942 -4186
rect 449026 -4422 449262 -4186
rect 448706 -4742 448942 -4506
rect 449026 -4742 449262 -4506
rect 452426 165818 452662 166054
rect 452746 165818 452982 166054
rect 452426 165498 452662 165734
rect 452746 165498 452982 165734
rect 452426 129818 452662 130054
rect 452746 129818 452982 130054
rect 452426 129498 452662 129734
rect 452746 129498 452982 129734
rect 452426 93818 452662 94054
rect 452746 93818 452982 94054
rect 452426 93498 452662 93734
rect 452746 93498 452982 93734
rect 452426 57818 452662 58054
rect 452746 57818 452982 58054
rect 452426 57498 452662 57734
rect 452746 57498 452982 57734
rect 452426 21818 452662 22054
rect 452746 21818 452982 22054
rect 452426 21498 452662 21734
rect 452746 21498 452982 21734
rect 452426 -5382 452662 -5146
rect 452746 -5382 452982 -5146
rect 452426 -5702 452662 -5466
rect 452746 -5702 452982 -5466
rect 456146 169538 456382 169774
rect 456466 169538 456702 169774
rect 456146 169218 456382 169454
rect 456466 169218 456702 169454
rect 456146 133538 456382 133774
rect 456466 133538 456702 133774
rect 456146 133218 456382 133454
rect 456466 133218 456702 133454
rect 456146 97538 456382 97774
rect 456466 97538 456702 97774
rect 456146 97218 456382 97454
rect 456466 97218 456702 97454
rect 456146 61538 456382 61774
rect 456466 61538 456702 61774
rect 456146 61218 456382 61454
rect 456466 61218 456702 61454
rect 456146 25538 456382 25774
rect 456466 25538 456702 25774
rect 456146 25218 456382 25454
rect 456466 25218 456702 25454
rect 456146 -6342 456382 -6106
rect 456466 -6342 456702 -6106
rect 456146 -6662 456382 -6426
rect 456466 -6662 456702 -6426
rect 459866 173258 460102 173494
rect 460186 173258 460422 173494
rect 459866 172938 460102 173174
rect 460186 172938 460422 173174
rect 459866 137258 460102 137494
rect 460186 137258 460422 137494
rect 459866 136938 460102 137174
rect 460186 136938 460422 137174
rect 459866 101258 460102 101494
rect 460186 101258 460422 101494
rect 459866 100938 460102 101174
rect 460186 100938 460422 101174
rect 459866 65258 460102 65494
rect 460186 65258 460422 65494
rect 459866 64938 460102 65174
rect 460186 64938 460422 65174
rect 459866 29258 460102 29494
rect 460186 29258 460422 29494
rect 459866 28938 460102 29174
rect 460186 28938 460422 29174
rect 459866 -7302 460102 -7066
rect 460186 -7302 460422 -7066
rect 459866 -7622 460102 -7386
rect 460186 -7622 460422 -7386
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -1542 473782 -1306
rect 473866 -1542 474102 -1306
rect 473546 -1862 473782 -1626
rect 473866 -1862 474102 -1626
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -2502 477502 -2266
rect 477586 -2502 477822 -2266
rect 477266 -2822 477502 -2586
rect 477586 -2822 477822 -2586
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 480986 -3462 481222 -3226
rect 481306 -3462 481542 -3226
rect 480986 -3782 481222 -3546
rect 481306 -3782 481542 -3546
rect 484706 162098 484942 162334
rect 485026 162098 485262 162334
rect 484706 161778 484942 162014
rect 485026 161778 485262 162014
rect 484706 126098 484942 126334
rect 485026 126098 485262 126334
rect 484706 125778 484942 126014
rect 485026 125778 485262 126014
rect 484706 90098 484942 90334
rect 485026 90098 485262 90334
rect 484706 89778 484942 90014
rect 485026 89778 485262 90014
rect 484706 54098 484942 54334
rect 485026 54098 485262 54334
rect 484706 53778 484942 54014
rect 485026 53778 485262 54014
rect 484706 18098 484942 18334
rect 485026 18098 485262 18334
rect 484706 17778 484942 18014
rect 485026 17778 485262 18014
rect 484706 -4422 484942 -4186
rect 485026 -4422 485262 -4186
rect 484706 -4742 484942 -4506
rect 485026 -4742 485262 -4506
rect 488426 165818 488662 166054
rect 488746 165818 488982 166054
rect 488426 165498 488662 165734
rect 488746 165498 488982 165734
rect 488426 129818 488662 130054
rect 488746 129818 488982 130054
rect 488426 129498 488662 129734
rect 488746 129498 488982 129734
rect 488426 93818 488662 94054
rect 488746 93818 488982 94054
rect 488426 93498 488662 93734
rect 488746 93498 488982 93734
rect 488426 57818 488662 58054
rect 488746 57818 488982 58054
rect 488426 57498 488662 57734
rect 488746 57498 488982 57734
rect 488426 21818 488662 22054
rect 488746 21818 488982 22054
rect 488426 21498 488662 21734
rect 488746 21498 488982 21734
rect 488426 -5382 488662 -5146
rect 488746 -5382 488982 -5146
rect 488426 -5702 488662 -5466
rect 488746 -5702 488982 -5466
rect 492146 169538 492382 169774
rect 492466 169538 492702 169774
rect 492146 169218 492382 169454
rect 492466 169218 492702 169454
rect 492146 133538 492382 133774
rect 492466 133538 492702 133774
rect 492146 133218 492382 133454
rect 492466 133218 492702 133454
rect 492146 97538 492382 97774
rect 492466 97538 492702 97774
rect 492146 97218 492382 97454
rect 492466 97218 492702 97454
rect 492146 61538 492382 61774
rect 492466 61538 492702 61774
rect 492146 61218 492382 61454
rect 492466 61218 492702 61454
rect 492146 25538 492382 25774
rect 492466 25538 492702 25774
rect 492146 25218 492382 25454
rect 492466 25218 492702 25454
rect 492146 -6342 492382 -6106
rect 492466 -6342 492702 -6106
rect 492146 -6662 492382 -6426
rect 492466 -6662 492702 -6426
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 495866 173258 496102 173494
rect 496186 173258 496422 173494
rect 495866 172938 496102 173174
rect 496186 172938 496422 173174
rect 495866 137258 496102 137494
rect 496186 137258 496422 137494
rect 495866 136938 496102 137174
rect 496186 136938 496422 137174
rect 495866 101258 496102 101494
rect 496186 101258 496422 101494
rect 495866 100938 496102 101174
rect 496186 100938 496422 101174
rect 495866 65258 496102 65494
rect 496186 65258 496422 65494
rect 495866 64938 496102 65174
rect 496186 64938 496422 65174
rect 495866 29258 496102 29494
rect 496186 29258 496422 29494
rect 495866 28938 496102 29174
rect 496186 28938 496422 29174
rect 495866 -7302 496102 -7066
rect 496186 -7302 496422 -7066
rect 495866 -7622 496102 -7386
rect 496186 -7622 496422 -7386
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -1542 509782 -1306
rect 509866 -1542 510102 -1306
rect 509546 -1862 509782 -1626
rect 509866 -1862 510102 -1626
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 520706 594098 520942 594334
rect 521026 594098 521262 594334
rect 520706 593778 520942 594014
rect 521026 593778 521262 594014
rect 524426 597818 524662 598054
rect 524746 597818 524982 598054
rect 524426 597498 524662 597734
rect 524746 597498 524982 597734
rect 524426 561818 524662 562054
rect 524746 561818 524982 562054
rect 524426 561498 524662 561734
rect 524746 561498 524982 561734
rect 520706 558098 520942 558334
rect 521026 558098 521262 558334
rect 520706 557778 520942 558014
rect 521026 557778 521262 558014
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -2502 513502 -2266
rect 513586 -2502 513822 -2266
rect 513266 -2822 513502 -2586
rect 513586 -2822 513822 -2586
rect 520706 522098 520942 522334
rect 521026 522098 521262 522334
rect 520706 521778 520942 522014
rect 521026 521778 521262 522014
rect 520706 486098 520942 486334
rect 521026 486098 521262 486334
rect 520706 485778 520942 486014
rect 521026 485778 521262 486014
rect 520706 450098 520942 450334
rect 521026 450098 521262 450334
rect 520706 449778 520942 450014
rect 521026 449778 521262 450014
rect 520706 414098 520942 414334
rect 521026 414098 521262 414334
rect 520706 413778 520942 414014
rect 521026 413778 521262 414014
rect 520706 378098 520942 378334
rect 521026 378098 521262 378334
rect 520706 377778 520942 378014
rect 521026 377778 521262 378014
rect 520706 342098 520942 342334
rect 521026 342098 521262 342334
rect 520706 341778 520942 342014
rect 521026 341778 521262 342014
rect 520706 306098 520942 306334
rect 521026 306098 521262 306334
rect 520706 305778 520942 306014
rect 521026 305778 521262 306014
rect 520706 270098 520942 270334
rect 521026 270098 521262 270334
rect 520706 269778 520942 270014
rect 521026 269778 521262 270014
rect 520706 234098 520942 234334
rect 521026 234098 521262 234334
rect 520706 233778 520942 234014
rect 521026 233778 521262 234014
rect 520706 198098 520942 198334
rect 521026 198098 521262 198334
rect 520706 197778 520942 198014
rect 521026 197778 521262 198014
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 516986 -3462 517222 -3226
rect 517306 -3462 517542 -3226
rect 516986 -3782 517222 -3546
rect 517306 -3782 517542 -3546
rect 528146 565538 528382 565774
rect 528466 565538 528702 565774
rect 528146 565218 528382 565454
rect 528466 565218 528702 565454
rect 524426 525818 524662 526054
rect 524746 525818 524982 526054
rect 524426 525498 524662 525734
rect 524746 525498 524982 525734
rect 524426 489818 524662 490054
rect 524746 489818 524982 490054
rect 524426 489498 524662 489734
rect 524746 489498 524982 489734
rect 524426 453818 524662 454054
rect 524746 453818 524982 454054
rect 524426 453498 524662 453734
rect 524746 453498 524982 453734
rect 524426 417818 524662 418054
rect 524746 417818 524982 418054
rect 524426 417498 524662 417734
rect 524746 417498 524982 417734
rect 524426 381818 524662 382054
rect 524746 381818 524982 382054
rect 524426 381498 524662 381734
rect 524746 381498 524982 381734
rect 524426 345818 524662 346054
rect 524746 345818 524982 346054
rect 524426 345498 524662 345734
rect 524746 345498 524982 345734
rect 524426 309818 524662 310054
rect 524746 309818 524982 310054
rect 524426 309498 524662 309734
rect 524746 309498 524982 309734
rect 524426 273818 524662 274054
rect 524746 273818 524982 274054
rect 524426 273498 524662 273734
rect 524746 273498 524982 273734
rect 524426 237818 524662 238054
rect 524746 237818 524982 238054
rect 524426 237498 524662 237734
rect 524746 237498 524982 237734
rect 524426 201818 524662 202054
rect 524746 201818 524982 202054
rect 524426 201498 524662 201734
rect 524746 201498 524982 201734
rect 520706 162098 520942 162334
rect 521026 162098 521262 162334
rect 520706 161778 520942 162014
rect 521026 161778 521262 162014
rect 520706 126098 520942 126334
rect 521026 126098 521262 126334
rect 520706 125778 520942 126014
rect 521026 125778 521262 126014
rect 520706 90098 520942 90334
rect 521026 90098 521262 90334
rect 520706 89778 520942 90014
rect 521026 89778 521262 90014
rect 520706 54098 520942 54334
rect 521026 54098 521262 54334
rect 520706 53778 520942 54014
rect 521026 53778 521262 54014
rect 520706 18098 520942 18334
rect 521026 18098 521262 18334
rect 520706 17778 520942 18014
rect 521026 17778 521262 18014
rect 520706 -4422 520942 -4186
rect 521026 -4422 521262 -4186
rect 520706 -4742 520942 -4506
rect 521026 -4742 521262 -4506
rect 531866 569258 532102 569494
rect 532186 569258 532422 569494
rect 531866 568938 532102 569174
rect 532186 568938 532422 569174
rect 528146 529538 528382 529774
rect 528466 529538 528702 529774
rect 528146 529218 528382 529454
rect 528466 529218 528702 529454
rect 528146 493538 528382 493774
rect 528466 493538 528702 493774
rect 528146 493218 528382 493454
rect 528466 493218 528702 493454
rect 531866 533258 532102 533494
rect 532186 533258 532422 533494
rect 531866 532938 532102 533174
rect 532186 532938 532422 533174
rect 528146 457538 528382 457774
rect 528466 457538 528702 457774
rect 528146 457218 528382 457454
rect 528466 457218 528702 457454
rect 528146 421538 528382 421774
rect 528466 421538 528702 421774
rect 528146 421218 528382 421454
rect 528466 421218 528702 421454
rect 528146 385538 528382 385774
rect 528466 385538 528702 385774
rect 528146 385218 528382 385454
rect 528466 385218 528702 385454
rect 528146 349538 528382 349774
rect 528466 349538 528702 349774
rect 528146 349218 528382 349454
rect 528466 349218 528702 349454
rect 528146 313538 528382 313774
rect 528466 313538 528702 313774
rect 528146 313218 528382 313454
rect 528466 313218 528702 313454
rect 528146 277538 528382 277774
rect 528466 277538 528702 277774
rect 528146 277218 528382 277454
rect 528466 277218 528702 277454
rect 528146 241538 528382 241774
rect 528466 241538 528702 241774
rect 528146 241218 528382 241454
rect 528466 241218 528702 241454
rect 528146 205538 528382 205774
rect 528466 205538 528702 205774
rect 528146 205218 528382 205454
rect 528466 205218 528702 205454
rect 524426 165818 524662 166054
rect 524746 165818 524982 166054
rect 524426 165498 524662 165734
rect 524746 165498 524982 165734
rect 524426 129818 524662 130054
rect 524746 129818 524982 130054
rect 524426 129498 524662 129734
rect 524746 129498 524982 129734
rect 524426 93818 524662 94054
rect 524746 93818 524982 94054
rect 524426 93498 524662 93734
rect 524746 93498 524982 93734
rect 524426 57818 524662 58054
rect 524746 57818 524982 58054
rect 524426 57498 524662 57734
rect 524746 57498 524982 57734
rect 524426 21818 524662 22054
rect 524746 21818 524982 22054
rect 524426 21498 524662 21734
rect 524746 21498 524982 21734
rect 524426 -5382 524662 -5146
rect 524746 -5382 524982 -5146
rect 524426 -5702 524662 -5466
rect 524746 -5702 524982 -5466
rect 531866 497258 532102 497494
rect 532186 497258 532422 497494
rect 531866 496938 532102 497174
rect 532186 496938 532422 497174
rect 531866 461258 532102 461494
rect 532186 461258 532422 461494
rect 531866 460938 532102 461174
rect 532186 460938 532422 461174
rect 531866 425258 532102 425494
rect 532186 425258 532422 425494
rect 531866 424938 532102 425174
rect 532186 424938 532422 425174
rect 531866 389258 532102 389494
rect 532186 389258 532422 389494
rect 531866 388938 532102 389174
rect 532186 388938 532422 389174
rect 531866 353258 532102 353494
rect 532186 353258 532422 353494
rect 531866 352938 532102 353174
rect 532186 352938 532422 353174
rect 531866 317258 532102 317494
rect 532186 317258 532422 317494
rect 531866 316938 532102 317174
rect 532186 316938 532422 317174
rect 531866 281258 532102 281494
rect 532186 281258 532422 281494
rect 531866 280938 532102 281174
rect 532186 280938 532422 281174
rect 531866 245258 532102 245494
rect 532186 245258 532422 245494
rect 531866 244938 532102 245174
rect 532186 244938 532422 245174
rect 531866 209258 532102 209494
rect 532186 209258 532422 209494
rect 531866 208938 532102 209174
rect 532186 208938 532422 209174
rect 528146 169538 528382 169774
rect 528466 169538 528702 169774
rect 528146 169218 528382 169454
rect 528466 169218 528702 169454
rect 528146 133538 528382 133774
rect 528466 133538 528702 133774
rect 528146 133218 528382 133454
rect 528466 133218 528702 133454
rect 528146 97538 528382 97774
rect 528466 97538 528702 97774
rect 528146 97218 528382 97454
rect 528466 97218 528702 97454
rect 528146 61538 528382 61774
rect 528466 61538 528702 61774
rect 528146 61218 528382 61454
rect 528466 61218 528702 61454
rect 528146 25538 528382 25774
rect 528466 25538 528702 25774
rect 528146 25218 528382 25454
rect 528466 25218 528702 25454
rect 528146 -6342 528382 -6106
rect 528466 -6342 528702 -6106
rect 528146 -6662 528382 -6426
rect 528466 -6662 528702 -6426
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 549266 706522 549502 706758
rect 549586 706522 549822 706758
rect 549266 706202 549502 706438
rect 549586 706202 549822 706438
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 531866 173258 532102 173494
rect 532186 173258 532422 173494
rect 531866 172938 532102 173174
rect 532186 172938 532422 173174
rect 531866 137258 532102 137494
rect 532186 137258 532422 137494
rect 531866 136938 532102 137174
rect 532186 136938 532422 137174
rect 531866 101258 532102 101494
rect 532186 101258 532422 101494
rect 531866 100938 532102 101174
rect 532186 100938 532422 101174
rect 531866 65258 532102 65494
rect 532186 65258 532422 65494
rect 531866 64938 532102 65174
rect 532186 64938 532422 65174
rect 531866 29258 532102 29494
rect 532186 29258 532422 29494
rect 531866 28938 532102 29174
rect 532186 28938 532422 29174
rect 531866 -7302 532102 -7066
rect 532186 -7302 532422 -7066
rect 531866 -7622 532102 -7386
rect 532186 -7622 532422 -7386
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 552986 707482 553222 707718
rect 553306 707482 553542 707718
rect 552986 707162 553222 707398
rect 553306 707162 553542 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 556706 708442 556942 708678
rect 557026 708442 557262 708678
rect 556706 708122 556942 708358
rect 557026 708122 557262 708358
rect 560426 709402 560662 709638
rect 560746 709402 560982 709638
rect 560426 709082 560662 709318
rect 560746 709082 560982 709318
rect 556706 666098 556942 666334
rect 557026 666098 557262 666334
rect 556706 665778 556942 666014
rect 557026 665778 557262 666014
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -1542 545782 -1306
rect 545866 -1542 546102 -1306
rect 545546 -1862 545782 -1626
rect 545866 -1862 546102 -1626
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -2502 549502 -2266
rect 549586 -2502 549822 -2266
rect 549266 -2822 549502 -2586
rect 549586 -2822 549822 -2586
rect 556706 630098 556942 630334
rect 557026 630098 557262 630334
rect 556706 629778 556942 630014
rect 557026 629778 557262 630014
rect 556706 594098 556942 594334
rect 557026 594098 557262 594334
rect 556706 593778 556942 594014
rect 557026 593778 557262 594014
rect 556706 558098 556942 558334
rect 557026 558098 557262 558334
rect 556706 557778 556942 558014
rect 557026 557778 557262 558014
rect 556706 522098 556942 522334
rect 557026 522098 557262 522334
rect 556706 521778 556942 522014
rect 557026 521778 557262 522014
rect 556706 486098 556942 486334
rect 557026 486098 557262 486334
rect 556706 485778 556942 486014
rect 557026 485778 557262 486014
rect 556706 450098 556942 450334
rect 557026 450098 557262 450334
rect 556706 449778 556942 450014
rect 557026 449778 557262 450014
rect 556706 414098 556942 414334
rect 557026 414098 557262 414334
rect 556706 413778 556942 414014
rect 557026 413778 557262 414014
rect 556706 378098 556942 378334
rect 557026 378098 557262 378334
rect 556706 377778 556942 378014
rect 557026 377778 557262 378014
rect 556706 342098 556942 342334
rect 557026 342098 557262 342334
rect 556706 341778 556942 342014
rect 557026 341778 557262 342014
rect 556706 306098 556942 306334
rect 557026 306098 557262 306334
rect 556706 305778 556942 306014
rect 557026 305778 557262 306014
rect 556706 270098 556942 270334
rect 557026 270098 557262 270334
rect 556706 269778 556942 270014
rect 557026 269778 557262 270014
rect 556706 234098 556942 234334
rect 557026 234098 557262 234334
rect 556706 233778 556942 234014
rect 557026 233778 557262 234014
rect 556706 198098 556942 198334
rect 557026 198098 557262 198334
rect 556706 197778 556942 198014
rect 557026 197778 557262 198014
rect 556706 162098 556942 162334
rect 557026 162098 557262 162334
rect 556706 161778 556942 162014
rect 557026 161778 557262 162014
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 552986 -3462 553222 -3226
rect 553306 -3462 553542 -3226
rect 552986 -3782 553222 -3546
rect 553306 -3782 553542 -3546
rect 560426 669818 560662 670054
rect 560746 669818 560982 670054
rect 560426 669498 560662 669734
rect 560746 669498 560982 669734
rect 560426 633818 560662 634054
rect 560746 633818 560982 634054
rect 560426 633498 560662 633734
rect 560746 633498 560982 633734
rect 560426 597818 560662 598054
rect 560746 597818 560982 598054
rect 560426 597498 560662 597734
rect 560746 597498 560982 597734
rect 560426 561818 560662 562054
rect 560746 561818 560982 562054
rect 560426 561498 560662 561734
rect 560746 561498 560982 561734
rect 560426 525818 560662 526054
rect 560746 525818 560982 526054
rect 560426 525498 560662 525734
rect 560746 525498 560982 525734
rect 560426 489818 560662 490054
rect 560746 489818 560982 490054
rect 560426 489498 560662 489734
rect 560746 489498 560982 489734
rect 560426 453818 560662 454054
rect 560746 453818 560982 454054
rect 560426 453498 560662 453734
rect 560746 453498 560982 453734
rect 560426 417818 560662 418054
rect 560746 417818 560982 418054
rect 560426 417498 560662 417734
rect 560746 417498 560982 417734
rect 560426 381818 560662 382054
rect 560746 381818 560982 382054
rect 560426 381498 560662 381734
rect 560746 381498 560982 381734
rect 560426 345818 560662 346054
rect 560746 345818 560982 346054
rect 560426 345498 560662 345734
rect 560746 345498 560982 345734
rect 560426 309818 560662 310054
rect 560746 309818 560982 310054
rect 560426 309498 560662 309734
rect 560746 309498 560982 309734
rect 560426 273818 560662 274054
rect 560746 273818 560982 274054
rect 560426 273498 560662 273734
rect 560746 273498 560982 273734
rect 560426 237818 560662 238054
rect 560746 237818 560982 238054
rect 560426 237498 560662 237734
rect 560746 237498 560982 237734
rect 560426 201818 560662 202054
rect 560746 201818 560982 202054
rect 560426 201498 560662 201734
rect 560746 201498 560982 201734
rect 560426 165818 560662 166054
rect 560746 165818 560982 166054
rect 560426 165498 560662 165734
rect 560746 165498 560982 165734
rect 556706 126098 556942 126334
rect 557026 126098 557262 126334
rect 556706 125778 556942 126014
rect 557026 125778 557262 126014
rect 556706 90098 556942 90334
rect 557026 90098 557262 90334
rect 556706 89778 556942 90014
rect 557026 89778 557262 90014
rect 556706 54098 556942 54334
rect 557026 54098 557262 54334
rect 556706 53778 556942 54014
rect 557026 53778 557262 54014
rect 556706 18098 556942 18334
rect 557026 18098 557262 18334
rect 556706 17778 556942 18014
rect 557026 17778 557262 18014
rect 556706 -4422 556942 -4186
rect 557026 -4422 557262 -4186
rect 556706 -4742 556942 -4506
rect 557026 -4742 557262 -4506
rect 560426 129818 560662 130054
rect 560746 129818 560982 130054
rect 560426 129498 560662 129734
rect 560746 129498 560982 129734
rect 560426 93818 560662 94054
rect 560746 93818 560982 94054
rect 560426 93498 560662 93734
rect 560746 93498 560982 93734
rect 560426 57818 560662 58054
rect 560746 57818 560982 58054
rect 560426 57498 560662 57734
rect 560746 57498 560982 57734
rect 560426 21818 560662 22054
rect 560746 21818 560982 22054
rect 560426 21498 560662 21734
rect 560746 21498 560982 21734
rect 560426 -5382 560662 -5146
rect 560746 -5382 560982 -5146
rect 560426 -5702 560662 -5466
rect 560746 -5702 560982 -5466
rect 564146 710362 564382 710598
rect 564466 710362 564702 710598
rect 564146 710042 564382 710278
rect 564466 710042 564702 710278
rect 564146 673538 564382 673774
rect 564466 673538 564702 673774
rect 564146 673218 564382 673454
rect 564466 673218 564702 673454
rect 564146 637538 564382 637774
rect 564466 637538 564702 637774
rect 564146 637218 564382 637454
rect 564466 637218 564702 637454
rect 564146 601538 564382 601774
rect 564466 601538 564702 601774
rect 564146 601218 564382 601454
rect 564466 601218 564702 601454
rect 564146 565538 564382 565774
rect 564466 565538 564702 565774
rect 564146 565218 564382 565454
rect 564466 565218 564702 565454
rect 564146 529538 564382 529774
rect 564466 529538 564702 529774
rect 564146 529218 564382 529454
rect 564466 529218 564702 529454
rect 564146 493538 564382 493774
rect 564466 493538 564702 493774
rect 564146 493218 564382 493454
rect 564466 493218 564702 493454
rect 564146 457538 564382 457774
rect 564466 457538 564702 457774
rect 564146 457218 564382 457454
rect 564466 457218 564702 457454
rect 564146 421538 564382 421774
rect 564466 421538 564702 421774
rect 564146 421218 564382 421454
rect 564466 421218 564702 421454
rect 564146 385538 564382 385774
rect 564466 385538 564702 385774
rect 564146 385218 564382 385454
rect 564466 385218 564702 385454
rect 564146 349538 564382 349774
rect 564466 349538 564702 349774
rect 564146 349218 564382 349454
rect 564466 349218 564702 349454
rect 564146 313538 564382 313774
rect 564466 313538 564702 313774
rect 564146 313218 564382 313454
rect 564466 313218 564702 313454
rect 564146 277538 564382 277774
rect 564466 277538 564702 277774
rect 564146 277218 564382 277454
rect 564466 277218 564702 277454
rect 564146 241538 564382 241774
rect 564466 241538 564702 241774
rect 564146 241218 564382 241454
rect 564466 241218 564702 241454
rect 564146 205538 564382 205774
rect 564466 205538 564702 205774
rect 564146 205218 564382 205454
rect 564466 205218 564702 205454
rect 564146 169538 564382 169774
rect 564466 169538 564702 169774
rect 564146 169218 564382 169454
rect 564466 169218 564702 169454
rect 564146 133538 564382 133774
rect 564466 133538 564702 133774
rect 564146 133218 564382 133454
rect 564466 133218 564702 133454
rect 564146 97538 564382 97774
rect 564466 97538 564702 97774
rect 564146 97218 564382 97454
rect 564466 97218 564702 97454
rect 564146 61538 564382 61774
rect 564466 61538 564702 61774
rect 564146 61218 564382 61454
rect 564466 61218 564702 61454
rect 564146 25538 564382 25774
rect 564466 25538 564702 25774
rect 564146 25218 564382 25454
rect 564466 25218 564702 25454
rect 564146 -6342 564382 -6106
rect 564466 -6342 564702 -6106
rect 564146 -6662 564382 -6426
rect 564466 -6662 564702 -6426
rect 567866 711322 568102 711558
rect 568186 711322 568422 711558
rect 567866 711002 568102 711238
rect 568186 711002 568422 711238
rect 567866 677258 568102 677494
rect 568186 677258 568422 677494
rect 567866 676938 568102 677174
rect 568186 676938 568422 677174
rect 567866 641258 568102 641494
rect 568186 641258 568422 641494
rect 567866 640938 568102 641174
rect 568186 640938 568422 641174
rect 567866 605258 568102 605494
rect 568186 605258 568422 605494
rect 567866 604938 568102 605174
rect 568186 604938 568422 605174
rect 567866 569258 568102 569494
rect 568186 569258 568422 569494
rect 567866 568938 568102 569174
rect 568186 568938 568422 569174
rect 567866 533258 568102 533494
rect 568186 533258 568422 533494
rect 567866 532938 568102 533174
rect 568186 532938 568422 533174
rect 567866 497258 568102 497494
rect 568186 497258 568422 497494
rect 567866 496938 568102 497174
rect 568186 496938 568422 497174
rect 567866 461258 568102 461494
rect 568186 461258 568422 461494
rect 567866 460938 568102 461174
rect 568186 460938 568422 461174
rect 567866 425258 568102 425494
rect 568186 425258 568422 425494
rect 567866 424938 568102 425174
rect 568186 424938 568422 425174
rect 567866 389258 568102 389494
rect 568186 389258 568422 389494
rect 567866 388938 568102 389174
rect 568186 388938 568422 389174
rect 567866 353258 568102 353494
rect 568186 353258 568422 353494
rect 567866 352938 568102 353174
rect 568186 352938 568422 353174
rect 567866 317258 568102 317494
rect 568186 317258 568422 317494
rect 567866 316938 568102 317174
rect 568186 316938 568422 317174
rect 567866 281258 568102 281494
rect 568186 281258 568422 281494
rect 567866 280938 568102 281174
rect 568186 280938 568422 281174
rect 567866 245258 568102 245494
rect 568186 245258 568422 245494
rect 567866 244938 568102 245174
rect 568186 244938 568422 245174
rect 567866 209258 568102 209494
rect 568186 209258 568422 209494
rect 567866 208938 568102 209174
rect 568186 208938 568422 209174
rect 567866 173258 568102 173494
rect 568186 173258 568422 173494
rect 567866 172938 568102 173174
rect 568186 172938 568422 173174
rect 567866 137258 568102 137494
rect 568186 137258 568422 137494
rect 567866 136938 568102 137174
rect 568186 136938 568422 137174
rect 567866 101258 568102 101494
rect 568186 101258 568422 101494
rect 567866 100938 568102 101174
rect 568186 100938 568422 101174
rect 567866 65258 568102 65494
rect 568186 65258 568422 65494
rect 567866 64938 568102 65174
rect 568186 64938 568422 65174
rect 567866 29258 568102 29494
rect 568186 29258 568422 29494
rect 567866 28938 568102 29174
rect 568186 28938 568422 29174
rect 567866 -7302 568102 -7066
rect 568186 -7302 568422 -7066
rect 567866 -7622 568102 -7386
rect 568186 -7622 568422 -7386
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 581546 705562 581782 705798
rect 581866 705562 582102 705798
rect 581546 705242 581782 705478
rect 581866 705242 582102 705478
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 690938 586538 691174
rect 586622 690938 586858 691174
rect 586302 690618 586538 690854
rect 586622 690618 586858 690854
rect 586302 654938 586538 655174
rect 586622 654938 586858 655174
rect 586302 654618 586538 654854
rect 586622 654618 586858 654854
rect 586302 618938 586538 619174
rect 586622 618938 586858 619174
rect 586302 618618 586538 618854
rect 586622 618618 586858 618854
rect 586302 582938 586538 583174
rect 586622 582938 586858 583174
rect 586302 582618 586538 582854
rect 586622 582618 586858 582854
rect 586302 546938 586538 547174
rect 586622 546938 586858 547174
rect 586302 546618 586538 546854
rect 586622 546618 586858 546854
rect 586302 510938 586538 511174
rect 586622 510938 586858 511174
rect 586302 510618 586538 510854
rect 586622 510618 586858 510854
rect 586302 474938 586538 475174
rect 586622 474938 586858 475174
rect 586302 474618 586538 474854
rect 586622 474618 586858 474854
rect 586302 438938 586538 439174
rect 586622 438938 586858 439174
rect 586302 438618 586538 438854
rect 586622 438618 586858 438854
rect 586302 402938 586538 403174
rect 586622 402938 586858 403174
rect 586302 402618 586538 402854
rect 586622 402618 586858 402854
rect 586302 366938 586538 367174
rect 586622 366938 586858 367174
rect 586302 366618 586538 366854
rect 586622 366618 586858 366854
rect 586302 330938 586538 331174
rect 586622 330938 586858 331174
rect 586302 330618 586538 330854
rect 586622 330618 586858 330854
rect 586302 294938 586538 295174
rect 586622 294938 586858 295174
rect 586302 294618 586538 294854
rect 586622 294618 586858 294854
rect 586302 258938 586538 259174
rect 586622 258938 586858 259174
rect 586302 258618 586538 258854
rect 586622 258618 586858 258854
rect 586302 222938 586538 223174
rect 586622 222938 586858 223174
rect 586302 222618 586538 222854
rect 586622 222618 586858 222854
rect 586302 186938 586538 187174
rect 586622 186938 586858 187174
rect 586302 186618 586538 186854
rect 586622 186618 586858 186854
rect 586302 150938 586538 151174
rect 586622 150938 586858 151174
rect 586302 150618 586538 150854
rect 586622 150618 586858 150854
rect 586302 114938 586538 115174
rect 586622 114938 586858 115174
rect 586302 114618 586538 114854
rect 586622 114618 586858 114854
rect 586302 78938 586538 79174
rect 586622 78938 586858 79174
rect 586302 78618 586538 78854
rect 586622 78618 586858 78854
rect 586302 42938 586538 43174
rect 586622 42938 586858 43174
rect 586302 42618 586538 42854
rect 586622 42618 586858 42854
rect 586302 6938 586538 7174
rect 586622 6938 586858 7174
rect 586302 6618 586538 6854
rect 586622 6618 586858 6854
rect 581546 -1542 581782 -1306
rect 581866 -1542 582102 -1306
rect 581546 -1862 581782 -1626
rect 581866 -1862 582102 -1626
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 694658 587498 694894
rect 587582 694658 587818 694894
rect 587262 694338 587498 694574
rect 587582 694338 587818 694574
rect 587262 658658 587498 658894
rect 587582 658658 587818 658894
rect 587262 658338 587498 658574
rect 587582 658338 587818 658574
rect 587262 622658 587498 622894
rect 587582 622658 587818 622894
rect 587262 622338 587498 622574
rect 587582 622338 587818 622574
rect 587262 586658 587498 586894
rect 587582 586658 587818 586894
rect 587262 586338 587498 586574
rect 587582 586338 587818 586574
rect 587262 550658 587498 550894
rect 587582 550658 587818 550894
rect 587262 550338 587498 550574
rect 587582 550338 587818 550574
rect 587262 514658 587498 514894
rect 587582 514658 587818 514894
rect 587262 514338 587498 514574
rect 587582 514338 587818 514574
rect 587262 478658 587498 478894
rect 587582 478658 587818 478894
rect 587262 478338 587498 478574
rect 587582 478338 587818 478574
rect 587262 442658 587498 442894
rect 587582 442658 587818 442894
rect 587262 442338 587498 442574
rect 587582 442338 587818 442574
rect 587262 406658 587498 406894
rect 587582 406658 587818 406894
rect 587262 406338 587498 406574
rect 587582 406338 587818 406574
rect 587262 370658 587498 370894
rect 587582 370658 587818 370894
rect 587262 370338 587498 370574
rect 587582 370338 587818 370574
rect 587262 334658 587498 334894
rect 587582 334658 587818 334894
rect 587262 334338 587498 334574
rect 587582 334338 587818 334574
rect 587262 298658 587498 298894
rect 587582 298658 587818 298894
rect 587262 298338 587498 298574
rect 587582 298338 587818 298574
rect 587262 262658 587498 262894
rect 587582 262658 587818 262894
rect 587262 262338 587498 262574
rect 587582 262338 587818 262574
rect 587262 226658 587498 226894
rect 587582 226658 587818 226894
rect 587262 226338 587498 226574
rect 587582 226338 587818 226574
rect 587262 190658 587498 190894
rect 587582 190658 587818 190894
rect 587262 190338 587498 190574
rect 587582 190338 587818 190574
rect 587262 154658 587498 154894
rect 587582 154658 587818 154894
rect 587262 154338 587498 154574
rect 587582 154338 587818 154574
rect 587262 118658 587498 118894
rect 587582 118658 587818 118894
rect 587262 118338 587498 118574
rect 587582 118338 587818 118574
rect 587262 82658 587498 82894
rect 587582 82658 587818 82894
rect 587262 82338 587498 82574
rect 587582 82338 587818 82574
rect 587262 46658 587498 46894
rect 587582 46658 587818 46894
rect 587262 46338 587498 46574
rect 587582 46338 587818 46574
rect 587262 10658 587498 10894
rect 587582 10658 587818 10894
rect 587262 10338 587498 10574
rect 587582 10338 587818 10574
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 698378 588458 698614
rect 588542 698378 588778 698614
rect 588222 698058 588458 698294
rect 588542 698058 588778 698294
rect 588222 662378 588458 662614
rect 588542 662378 588778 662614
rect 588222 662058 588458 662294
rect 588542 662058 588778 662294
rect 588222 626378 588458 626614
rect 588542 626378 588778 626614
rect 588222 626058 588458 626294
rect 588542 626058 588778 626294
rect 588222 590378 588458 590614
rect 588542 590378 588778 590614
rect 588222 590058 588458 590294
rect 588542 590058 588778 590294
rect 588222 554378 588458 554614
rect 588542 554378 588778 554614
rect 588222 554058 588458 554294
rect 588542 554058 588778 554294
rect 588222 518378 588458 518614
rect 588542 518378 588778 518614
rect 588222 518058 588458 518294
rect 588542 518058 588778 518294
rect 588222 482378 588458 482614
rect 588542 482378 588778 482614
rect 588222 482058 588458 482294
rect 588542 482058 588778 482294
rect 588222 446378 588458 446614
rect 588542 446378 588778 446614
rect 588222 446058 588458 446294
rect 588542 446058 588778 446294
rect 588222 410378 588458 410614
rect 588542 410378 588778 410614
rect 588222 410058 588458 410294
rect 588542 410058 588778 410294
rect 588222 374378 588458 374614
rect 588542 374378 588778 374614
rect 588222 374058 588458 374294
rect 588542 374058 588778 374294
rect 588222 338378 588458 338614
rect 588542 338378 588778 338614
rect 588222 338058 588458 338294
rect 588542 338058 588778 338294
rect 588222 302378 588458 302614
rect 588542 302378 588778 302614
rect 588222 302058 588458 302294
rect 588542 302058 588778 302294
rect 588222 266378 588458 266614
rect 588542 266378 588778 266614
rect 588222 266058 588458 266294
rect 588542 266058 588778 266294
rect 588222 230378 588458 230614
rect 588542 230378 588778 230614
rect 588222 230058 588458 230294
rect 588542 230058 588778 230294
rect 588222 194378 588458 194614
rect 588542 194378 588778 194614
rect 588222 194058 588458 194294
rect 588542 194058 588778 194294
rect 588222 158378 588458 158614
rect 588542 158378 588778 158614
rect 588222 158058 588458 158294
rect 588542 158058 588778 158294
rect 588222 122378 588458 122614
rect 588542 122378 588778 122614
rect 588222 122058 588458 122294
rect 588542 122058 588778 122294
rect 588222 86378 588458 86614
rect 588542 86378 588778 86614
rect 588222 86058 588458 86294
rect 588542 86058 588778 86294
rect 588222 50378 588458 50614
rect 588542 50378 588778 50614
rect 588222 50058 588458 50294
rect 588542 50058 588778 50294
rect 588222 14378 588458 14614
rect 588542 14378 588778 14614
rect 588222 14058 588458 14294
rect 588542 14058 588778 14294
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 666098 589418 666334
rect 589502 666098 589738 666334
rect 589182 665778 589418 666014
rect 589502 665778 589738 666014
rect 589182 630098 589418 630334
rect 589502 630098 589738 630334
rect 589182 629778 589418 630014
rect 589502 629778 589738 630014
rect 589182 594098 589418 594334
rect 589502 594098 589738 594334
rect 589182 593778 589418 594014
rect 589502 593778 589738 594014
rect 589182 558098 589418 558334
rect 589502 558098 589738 558334
rect 589182 557778 589418 558014
rect 589502 557778 589738 558014
rect 589182 522098 589418 522334
rect 589502 522098 589738 522334
rect 589182 521778 589418 522014
rect 589502 521778 589738 522014
rect 589182 486098 589418 486334
rect 589502 486098 589738 486334
rect 589182 485778 589418 486014
rect 589502 485778 589738 486014
rect 589182 450098 589418 450334
rect 589502 450098 589738 450334
rect 589182 449778 589418 450014
rect 589502 449778 589738 450014
rect 589182 414098 589418 414334
rect 589502 414098 589738 414334
rect 589182 413778 589418 414014
rect 589502 413778 589738 414014
rect 589182 378098 589418 378334
rect 589502 378098 589738 378334
rect 589182 377778 589418 378014
rect 589502 377778 589738 378014
rect 589182 342098 589418 342334
rect 589502 342098 589738 342334
rect 589182 341778 589418 342014
rect 589502 341778 589738 342014
rect 589182 306098 589418 306334
rect 589502 306098 589738 306334
rect 589182 305778 589418 306014
rect 589502 305778 589738 306014
rect 589182 270098 589418 270334
rect 589502 270098 589738 270334
rect 589182 269778 589418 270014
rect 589502 269778 589738 270014
rect 589182 234098 589418 234334
rect 589502 234098 589738 234334
rect 589182 233778 589418 234014
rect 589502 233778 589738 234014
rect 589182 198098 589418 198334
rect 589502 198098 589738 198334
rect 589182 197778 589418 198014
rect 589502 197778 589738 198014
rect 589182 162098 589418 162334
rect 589502 162098 589738 162334
rect 589182 161778 589418 162014
rect 589502 161778 589738 162014
rect 589182 126098 589418 126334
rect 589502 126098 589738 126334
rect 589182 125778 589418 126014
rect 589502 125778 589738 126014
rect 589182 90098 589418 90334
rect 589502 90098 589738 90334
rect 589182 89778 589418 90014
rect 589502 89778 589738 90014
rect 589182 54098 589418 54334
rect 589502 54098 589738 54334
rect 589182 53778 589418 54014
rect 589502 53778 589738 54014
rect 589182 18098 589418 18334
rect 589502 18098 589738 18334
rect 589182 17778 589418 18014
rect 589502 17778 589738 18014
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 669818 590378 670054
rect 590462 669818 590698 670054
rect 590142 669498 590378 669734
rect 590462 669498 590698 669734
rect 590142 633818 590378 634054
rect 590462 633818 590698 634054
rect 590142 633498 590378 633734
rect 590462 633498 590698 633734
rect 590142 597818 590378 598054
rect 590462 597818 590698 598054
rect 590142 597498 590378 597734
rect 590462 597498 590698 597734
rect 590142 561818 590378 562054
rect 590462 561818 590698 562054
rect 590142 561498 590378 561734
rect 590462 561498 590698 561734
rect 590142 525818 590378 526054
rect 590462 525818 590698 526054
rect 590142 525498 590378 525734
rect 590462 525498 590698 525734
rect 590142 489818 590378 490054
rect 590462 489818 590698 490054
rect 590142 489498 590378 489734
rect 590462 489498 590698 489734
rect 590142 453818 590378 454054
rect 590462 453818 590698 454054
rect 590142 453498 590378 453734
rect 590462 453498 590698 453734
rect 590142 417818 590378 418054
rect 590462 417818 590698 418054
rect 590142 417498 590378 417734
rect 590462 417498 590698 417734
rect 590142 381818 590378 382054
rect 590462 381818 590698 382054
rect 590142 381498 590378 381734
rect 590462 381498 590698 381734
rect 590142 345818 590378 346054
rect 590462 345818 590698 346054
rect 590142 345498 590378 345734
rect 590462 345498 590698 345734
rect 590142 309818 590378 310054
rect 590462 309818 590698 310054
rect 590142 309498 590378 309734
rect 590462 309498 590698 309734
rect 590142 273818 590378 274054
rect 590462 273818 590698 274054
rect 590142 273498 590378 273734
rect 590462 273498 590698 273734
rect 590142 237818 590378 238054
rect 590462 237818 590698 238054
rect 590142 237498 590378 237734
rect 590462 237498 590698 237734
rect 590142 201818 590378 202054
rect 590462 201818 590698 202054
rect 590142 201498 590378 201734
rect 590462 201498 590698 201734
rect 590142 165818 590378 166054
rect 590462 165818 590698 166054
rect 590142 165498 590378 165734
rect 590462 165498 590698 165734
rect 590142 129818 590378 130054
rect 590462 129818 590698 130054
rect 590142 129498 590378 129734
rect 590462 129498 590698 129734
rect 590142 93818 590378 94054
rect 590462 93818 590698 94054
rect 590142 93498 590378 93734
rect 590462 93498 590698 93734
rect 590142 57818 590378 58054
rect 590462 57818 590698 58054
rect 590142 57498 590378 57734
rect 590462 57498 590698 57734
rect 590142 21818 590378 22054
rect 590462 21818 590698 22054
rect 590142 21498 590378 21734
rect 590462 21498 590698 21734
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 673538 591338 673774
rect 591422 673538 591658 673774
rect 591102 673218 591338 673454
rect 591422 673218 591658 673454
rect 591102 637538 591338 637774
rect 591422 637538 591658 637774
rect 591102 637218 591338 637454
rect 591422 637218 591658 637454
rect 591102 601538 591338 601774
rect 591422 601538 591658 601774
rect 591102 601218 591338 601454
rect 591422 601218 591658 601454
rect 591102 565538 591338 565774
rect 591422 565538 591658 565774
rect 591102 565218 591338 565454
rect 591422 565218 591658 565454
rect 591102 529538 591338 529774
rect 591422 529538 591658 529774
rect 591102 529218 591338 529454
rect 591422 529218 591658 529454
rect 591102 493538 591338 493774
rect 591422 493538 591658 493774
rect 591102 493218 591338 493454
rect 591422 493218 591658 493454
rect 591102 457538 591338 457774
rect 591422 457538 591658 457774
rect 591102 457218 591338 457454
rect 591422 457218 591658 457454
rect 591102 421538 591338 421774
rect 591422 421538 591658 421774
rect 591102 421218 591338 421454
rect 591422 421218 591658 421454
rect 591102 385538 591338 385774
rect 591422 385538 591658 385774
rect 591102 385218 591338 385454
rect 591422 385218 591658 385454
rect 591102 349538 591338 349774
rect 591422 349538 591658 349774
rect 591102 349218 591338 349454
rect 591422 349218 591658 349454
rect 591102 313538 591338 313774
rect 591422 313538 591658 313774
rect 591102 313218 591338 313454
rect 591422 313218 591658 313454
rect 591102 277538 591338 277774
rect 591422 277538 591658 277774
rect 591102 277218 591338 277454
rect 591422 277218 591658 277454
rect 591102 241538 591338 241774
rect 591422 241538 591658 241774
rect 591102 241218 591338 241454
rect 591422 241218 591658 241454
rect 591102 205538 591338 205774
rect 591422 205538 591658 205774
rect 591102 205218 591338 205454
rect 591422 205218 591658 205454
rect 591102 169538 591338 169774
rect 591422 169538 591658 169774
rect 591102 169218 591338 169454
rect 591422 169218 591658 169454
rect 591102 133538 591338 133774
rect 591422 133538 591658 133774
rect 591102 133218 591338 133454
rect 591422 133218 591658 133454
rect 591102 97538 591338 97774
rect 591422 97538 591658 97774
rect 591102 97218 591338 97454
rect 591422 97218 591658 97454
rect 591102 61538 591338 61774
rect 591422 61538 591658 61774
rect 591102 61218 591338 61454
rect 591422 61218 591658 61454
rect 591102 25538 591338 25774
rect 591422 25538 591658 25774
rect 591102 25218 591338 25454
rect 591422 25218 591658 25454
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 677258 592298 677494
rect 592382 677258 592618 677494
rect 592062 676938 592298 677174
rect 592382 676938 592618 677174
rect 592062 641258 592298 641494
rect 592382 641258 592618 641494
rect 592062 640938 592298 641174
rect 592382 640938 592618 641174
rect 592062 605258 592298 605494
rect 592382 605258 592618 605494
rect 592062 604938 592298 605174
rect 592382 604938 592618 605174
rect 592062 569258 592298 569494
rect 592382 569258 592618 569494
rect 592062 568938 592298 569174
rect 592382 568938 592618 569174
rect 592062 533258 592298 533494
rect 592382 533258 592618 533494
rect 592062 532938 592298 533174
rect 592382 532938 592618 533174
rect 592062 497258 592298 497494
rect 592382 497258 592618 497494
rect 592062 496938 592298 497174
rect 592382 496938 592618 497174
rect 592062 461258 592298 461494
rect 592382 461258 592618 461494
rect 592062 460938 592298 461174
rect 592382 460938 592618 461174
rect 592062 425258 592298 425494
rect 592382 425258 592618 425494
rect 592062 424938 592298 425174
rect 592382 424938 592618 425174
rect 592062 389258 592298 389494
rect 592382 389258 592618 389494
rect 592062 388938 592298 389174
rect 592382 388938 592618 389174
rect 592062 353258 592298 353494
rect 592382 353258 592618 353494
rect 592062 352938 592298 353174
rect 592382 352938 592618 353174
rect 592062 317258 592298 317494
rect 592382 317258 592618 317494
rect 592062 316938 592298 317174
rect 592382 316938 592618 317174
rect 592062 281258 592298 281494
rect 592382 281258 592618 281494
rect 592062 280938 592298 281174
rect 592382 280938 592618 281174
rect 592062 245258 592298 245494
rect 592382 245258 592618 245494
rect 592062 244938 592298 245174
rect 592382 244938 592618 245174
rect 592062 209258 592298 209494
rect 592382 209258 592618 209494
rect 592062 208938 592298 209174
rect 592382 208938 592618 209174
rect 592062 173258 592298 173494
rect 592382 173258 592618 173494
rect 592062 172938 592298 173174
rect 592382 172938 592618 173174
rect 592062 137258 592298 137494
rect 592382 137258 592618 137494
rect 592062 136938 592298 137174
rect 592382 136938 592618 137174
rect 592062 101258 592298 101494
rect 592382 101258 592618 101494
rect 592062 100938 592298 101174
rect 592382 100938 592618 101174
rect 592062 65258 592298 65494
rect 592382 65258 592618 65494
rect 592062 64938 592298 65174
rect 592382 64938 592618 65174
rect 592062 29258 592298 29494
rect 592382 29258 592618 29494
rect 592062 28938 592298 29174
rect 592382 28938 592618 29174
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 27866 711558
rect 28102 711322 28186 711558
rect 28422 711322 63866 711558
rect 64102 711322 64186 711558
rect 64422 711322 99866 711558
rect 100102 711322 100186 711558
rect 100422 711322 135866 711558
rect 136102 711322 136186 711558
rect 136422 711322 171866 711558
rect 172102 711322 172186 711558
rect 172422 711322 207866 711558
rect 208102 711322 208186 711558
rect 208422 711322 243866 711558
rect 244102 711322 244186 711558
rect 244422 711322 279866 711558
rect 280102 711322 280186 711558
rect 280422 711322 315866 711558
rect 316102 711322 316186 711558
rect 316422 711322 351866 711558
rect 352102 711322 352186 711558
rect 352422 711322 387866 711558
rect 388102 711322 388186 711558
rect 388422 711322 423866 711558
rect 424102 711322 424186 711558
rect 424422 711322 459866 711558
rect 460102 711322 460186 711558
rect 460422 711322 495866 711558
rect 496102 711322 496186 711558
rect 496422 711322 531866 711558
rect 532102 711322 532186 711558
rect 532422 711322 567866 711558
rect 568102 711322 568186 711558
rect 568422 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 27866 711238
rect 28102 711002 28186 711238
rect 28422 711002 63866 711238
rect 64102 711002 64186 711238
rect 64422 711002 99866 711238
rect 100102 711002 100186 711238
rect 100422 711002 135866 711238
rect 136102 711002 136186 711238
rect 136422 711002 171866 711238
rect 172102 711002 172186 711238
rect 172422 711002 207866 711238
rect 208102 711002 208186 711238
rect 208422 711002 243866 711238
rect 244102 711002 244186 711238
rect 244422 711002 279866 711238
rect 280102 711002 280186 711238
rect 280422 711002 315866 711238
rect 316102 711002 316186 711238
rect 316422 711002 351866 711238
rect 352102 711002 352186 711238
rect 352422 711002 387866 711238
rect 388102 711002 388186 711238
rect 388422 711002 423866 711238
rect 424102 711002 424186 711238
rect 424422 711002 459866 711238
rect 460102 711002 460186 711238
rect 460422 711002 495866 711238
rect 496102 711002 496186 711238
rect 496422 711002 531866 711238
rect 532102 711002 532186 711238
rect 532422 711002 567866 711238
rect 568102 711002 568186 711238
rect 568422 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 24146 710598
rect 24382 710362 24466 710598
rect 24702 710362 60146 710598
rect 60382 710362 60466 710598
rect 60702 710362 96146 710598
rect 96382 710362 96466 710598
rect 96702 710362 132146 710598
rect 132382 710362 132466 710598
rect 132702 710362 168146 710598
rect 168382 710362 168466 710598
rect 168702 710362 204146 710598
rect 204382 710362 204466 710598
rect 204702 710362 240146 710598
rect 240382 710362 240466 710598
rect 240702 710362 276146 710598
rect 276382 710362 276466 710598
rect 276702 710362 312146 710598
rect 312382 710362 312466 710598
rect 312702 710362 348146 710598
rect 348382 710362 348466 710598
rect 348702 710362 384146 710598
rect 384382 710362 384466 710598
rect 384702 710362 420146 710598
rect 420382 710362 420466 710598
rect 420702 710362 456146 710598
rect 456382 710362 456466 710598
rect 456702 710362 492146 710598
rect 492382 710362 492466 710598
rect 492702 710362 528146 710598
rect 528382 710362 528466 710598
rect 528702 710362 564146 710598
rect 564382 710362 564466 710598
rect 564702 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 24146 710278
rect 24382 710042 24466 710278
rect 24702 710042 60146 710278
rect 60382 710042 60466 710278
rect 60702 710042 96146 710278
rect 96382 710042 96466 710278
rect 96702 710042 132146 710278
rect 132382 710042 132466 710278
rect 132702 710042 168146 710278
rect 168382 710042 168466 710278
rect 168702 710042 204146 710278
rect 204382 710042 204466 710278
rect 204702 710042 240146 710278
rect 240382 710042 240466 710278
rect 240702 710042 276146 710278
rect 276382 710042 276466 710278
rect 276702 710042 312146 710278
rect 312382 710042 312466 710278
rect 312702 710042 348146 710278
rect 348382 710042 348466 710278
rect 348702 710042 384146 710278
rect 384382 710042 384466 710278
rect 384702 710042 420146 710278
rect 420382 710042 420466 710278
rect 420702 710042 456146 710278
rect 456382 710042 456466 710278
rect 456702 710042 492146 710278
rect 492382 710042 492466 710278
rect 492702 710042 528146 710278
rect 528382 710042 528466 710278
rect 528702 710042 564146 710278
rect 564382 710042 564466 710278
rect 564702 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 20426 709638
rect 20662 709402 20746 709638
rect 20982 709402 56426 709638
rect 56662 709402 56746 709638
rect 56982 709402 92426 709638
rect 92662 709402 92746 709638
rect 92982 709402 128426 709638
rect 128662 709402 128746 709638
rect 128982 709402 164426 709638
rect 164662 709402 164746 709638
rect 164982 709402 200426 709638
rect 200662 709402 200746 709638
rect 200982 709402 236426 709638
rect 236662 709402 236746 709638
rect 236982 709402 272426 709638
rect 272662 709402 272746 709638
rect 272982 709402 308426 709638
rect 308662 709402 308746 709638
rect 308982 709402 344426 709638
rect 344662 709402 344746 709638
rect 344982 709402 380426 709638
rect 380662 709402 380746 709638
rect 380982 709402 416426 709638
rect 416662 709402 416746 709638
rect 416982 709402 452426 709638
rect 452662 709402 452746 709638
rect 452982 709402 488426 709638
rect 488662 709402 488746 709638
rect 488982 709402 524426 709638
rect 524662 709402 524746 709638
rect 524982 709402 560426 709638
rect 560662 709402 560746 709638
rect 560982 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 20426 709318
rect 20662 709082 20746 709318
rect 20982 709082 56426 709318
rect 56662 709082 56746 709318
rect 56982 709082 92426 709318
rect 92662 709082 92746 709318
rect 92982 709082 128426 709318
rect 128662 709082 128746 709318
rect 128982 709082 164426 709318
rect 164662 709082 164746 709318
rect 164982 709082 200426 709318
rect 200662 709082 200746 709318
rect 200982 709082 236426 709318
rect 236662 709082 236746 709318
rect 236982 709082 272426 709318
rect 272662 709082 272746 709318
rect 272982 709082 308426 709318
rect 308662 709082 308746 709318
rect 308982 709082 344426 709318
rect 344662 709082 344746 709318
rect 344982 709082 380426 709318
rect 380662 709082 380746 709318
rect 380982 709082 416426 709318
rect 416662 709082 416746 709318
rect 416982 709082 452426 709318
rect 452662 709082 452746 709318
rect 452982 709082 488426 709318
rect 488662 709082 488746 709318
rect 488982 709082 524426 709318
rect 524662 709082 524746 709318
rect 524982 709082 560426 709318
rect 560662 709082 560746 709318
rect 560982 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 16706 708678
rect 16942 708442 17026 708678
rect 17262 708442 52706 708678
rect 52942 708442 53026 708678
rect 53262 708442 88706 708678
rect 88942 708442 89026 708678
rect 89262 708442 124706 708678
rect 124942 708442 125026 708678
rect 125262 708442 160706 708678
rect 160942 708442 161026 708678
rect 161262 708442 196706 708678
rect 196942 708442 197026 708678
rect 197262 708442 232706 708678
rect 232942 708442 233026 708678
rect 233262 708442 268706 708678
rect 268942 708442 269026 708678
rect 269262 708442 304706 708678
rect 304942 708442 305026 708678
rect 305262 708442 340706 708678
rect 340942 708442 341026 708678
rect 341262 708442 376706 708678
rect 376942 708442 377026 708678
rect 377262 708442 412706 708678
rect 412942 708442 413026 708678
rect 413262 708442 448706 708678
rect 448942 708442 449026 708678
rect 449262 708442 484706 708678
rect 484942 708442 485026 708678
rect 485262 708442 520706 708678
rect 520942 708442 521026 708678
rect 521262 708442 556706 708678
rect 556942 708442 557026 708678
rect 557262 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 16706 708358
rect 16942 708122 17026 708358
rect 17262 708122 52706 708358
rect 52942 708122 53026 708358
rect 53262 708122 88706 708358
rect 88942 708122 89026 708358
rect 89262 708122 124706 708358
rect 124942 708122 125026 708358
rect 125262 708122 160706 708358
rect 160942 708122 161026 708358
rect 161262 708122 196706 708358
rect 196942 708122 197026 708358
rect 197262 708122 232706 708358
rect 232942 708122 233026 708358
rect 233262 708122 268706 708358
rect 268942 708122 269026 708358
rect 269262 708122 304706 708358
rect 304942 708122 305026 708358
rect 305262 708122 340706 708358
rect 340942 708122 341026 708358
rect 341262 708122 376706 708358
rect 376942 708122 377026 708358
rect 377262 708122 412706 708358
rect 412942 708122 413026 708358
rect 413262 708122 448706 708358
rect 448942 708122 449026 708358
rect 449262 708122 484706 708358
rect 484942 708122 485026 708358
rect 485262 708122 520706 708358
rect 520942 708122 521026 708358
rect 521262 708122 556706 708358
rect 556942 708122 557026 708358
rect 557262 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 12986 707718
rect 13222 707482 13306 707718
rect 13542 707482 48986 707718
rect 49222 707482 49306 707718
rect 49542 707482 84986 707718
rect 85222 707482 85306 707718
rect 85542 707482 120986 707718
rect 121222 707482 121306 707718
rect 121542 707482 156986 707718
rect 157222 707482 157306 707718
rect 157542 707482 192986 707718
rect 193222 707482 193306 707718
rect 193542 707482 228986 707718
rect 229222 707482 229306 707718
rect 229542 707482 264986 707718
rect 265222 707482 265306 707718
rect 265542 707482 300986 707718
rect 301222 707482 301306 707718
rect 301542 707482 336986 707718
rect 337222 707482 337306 707718
rect 337542 707482 372986 707718
rect 373222 707482 373306 707718
rect 373542 707482 408986 707718
rect 409222 707482 409306 707718
rect 409542 707482 444986 707718
rect 445222 707482 445306 707718
rect 445542 707482 480986 707718
rect 481222 707482 481306 707718
rect 481542 707482 516986 707718
rect 517222 707482 517306 707718
rect 517542 707482 552986 707718
rect 553222 707482 553306 707718
rect 553542 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 12986 707398
rect 13222 707162 13306 707398
rect 13542 707162 48986 707398
rect 49222 707162 49306 707398
rect 49542 707162 84986 707398
rect 85222 707162 85306 707398
rect 85542 707162 120986 707398
rect 121222 707162 121306 707398
rect 121542 707162 156986 707398
rect 157222 707162 157306 707398
rect 157542 707162 192986 707398
rect 193222 707162 193306 707398
rect 193542 707162 228986 707398
rect 229222 707162 229306 707398
rect 229542 707162 264986 707398
rect 265222 707162 265306 707398
rect 265542 707162 300986 707398
rect 301222 707162 301306 707398
rect 301542 707162 336986 707398
rect 337222 707162 337306 707398
rect 337542 707162 372986 707398
rect 373222 707162 373306 707398
rect 373542 707162 408986 707398
rect 409222 707162 409306 707398
rect 409542 707162 444986 707398
rect 445222 707162 445306 707398
rect 445542 707162 480986 707398
rect 481222 707162 481306 707398
rect 481542 707162 516986 707398
rect 517222 707162 517306 707398
rect 517542 707162 552986 707398
rect 553222 707162 553306 707398
rect 553542 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 9266 706758
rect 9502 706522 9586 706758
rect 9822 706522 45266 706758
rect 45502 706522 45586 706758
rect 45822 706522 81266 706758
rect 81502 706522 81586 706758
rect 81822 706522 117266 706758
rect 117502 706522 117586 706758
rect 117822 706522 153266 706758
rect 153502 706522 153586 706758
rect 153822 706522 189266 706758
rect 189502 706522 189586 706758
rect 189822 706522 225266 706758
rect 225502 706522 225586 706758
rect 225822 706522 261266 706758
rect 261502 706522 261586 706758
rect 261822 706522 297266 706758
rect 297502 706522 297586 706758
rect 297822 706522 333266 706758
rect 333502 706522 333586 706758
rect 333822 706522 369266 706758
rect 369502 706522 369586 706758
rect 369822 706522 405266 706758
rect 405502 706522 405586 706758
rect 405822 706522 441266 706758
rect 441502 706522 441586 706758
rect 441822 706522 477266 706758
rect 477502 706522 477586 706758
rect 477822 706522 513266 706758
rect 513502 706522 513586 706758
rect 513822 706522 549266 706758
rect 549502 706522 549586 706758
rect 549822 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 9266 706438
rect 9502 706202 9586 706438
rect 9822 706202 45266 706438
rect 45502 706202 45586 706438
rect 45822 706202 81266 706438
rect 81502 706202 81586 706438
rect 81822 706202 117266 706438
rect 117502 706202 117586 706438
rect 117822 706202 153266 706438
rect 153502 706202 153586 706438
rect 153822 706202 189266 706438
rect 189502 706202 189586 706438
rect 189822 706202 225266 706438
rect 225502 706202 225586 706438
rect 225822 706202 261266 706438
rect 261502 706202 261586 706438
rect 261822 706202 297266 706438
rect 297502 706202 297586 706438
rect 297822 706202 333266 706438
rect 333502 706202 333586 706438
rect 333822 706202 369266 706438
rect 369502 706202 369586 706438
rect 369822 706202 405266 706438
rect 405502 706202 405586 706438
rect 405822 706202 441266 706438
rect 441502 706202 441586 706438
rect 441822 706202 477266 706438
rect 477502 706202 477586 706438
rect 477822 706202 513266 706438
rect 513502 706202 513586 706438
rect 513822 706202 549266 706438
rect 549502 706202 549586 706438
rect 549822 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 5546 705798
rect 5782 705562 5866 705798
rect 6102 705562 41546 705798
rect 41782 705562 41866 705798
rect 42102 705562 77546 705798
rect 77782 705562 77866 705798
rect 78102 705562 113546 705798
rect 113782 705562 113866 705798
rect 114102 705562 149546 705798
rect 149782 705562 149866 705798
rect 150102 705562 185546 705798
rect 185782 705562 185866 705798
rect 186102 705562 221546 705798
rect 221782 705562 221866 705798
rect 222102 705562 257546 705798
rect 257782 705562 257866 705798
rect 258102 705562 293546 705798
rect 293782 705562 293866 705798
rect 294102 705562 329546 705798
rect 329782 705562 329866 705798
rect 330102 705562 365546 705798
rect 365782 705562 365866 705798
rect 366102 705562 401546 705798
rect 401782 705562 401866 705798
rect 402102 705562 437546 705798
rect 437782 705562 437866 705798
rect 438102 705562 473546 705798
rect 473782 705562 473866 705798
rect 474102 705562 509546 705798
rect 509782 705562 509866 705798
rect 510102 705562 545546 705798
rect 545782 705562 545866 705798
rect 546102 705562 581546 705798
rect 581782 705562 581866 705798
rect 582102 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 5546 705478
rect 5782 705242 5866 705478
rect 6102 705242 41546 705478
rect 41782 705242 41866 705478
rect 42102 705242 77546 705478
rect 77782 705242 77866 705478
rect 78102 705242 113546 705478
rect 113782 705242 113866 705478
rect 114102 705242 149546 705478
rect 149782 705242 149866 705478
rect 150102 705242 185546 705478
rect 185782 705242 185866 705478
rect 186102 705242 221546 705478
rect 221782 705242 221866 705478
rect 222102 705242 257546 705478
rect 257782 705242 257866 705478
rect 258102 705242 293546 705478
rect 293782 705242 293866 705478
rect 294102 705242 329546 705478
rect 329782 705242 329866 705478
rect 330102 705242 365546 705478
rect 365782 705242 365866 705478
rect 366102 705242 401546 705478
rect 401782 705242 401866 705478
rect 402102 705242 437546 705478
rect 437782 705242 437866 705478
rect 438102 705242 473546 705478
rect 473782 705242 473866 705478
rect 474102 705242 509546 705478
rect 509782 705242 509866 705478
rect 510102 705242 545546 705478
rect 545782 705242 545866 705478
rect 546102 705242 581546 705478
rect 581782 705242 581866 705478
rect 582102 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -4854 698614
rect -4618 698378 -4534 698614
rect -4298 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 588222 698614
rect 588458 698378 588542 698614
rect 588778 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -4854 698294
rect -4618 698058 -4534 698294
rect -4298 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 588222 698294
rect 588458 698058 588542 698294
rect 588778 698058 592650 698294
rect -8726 698026 592650 698058
rect -8726 694894 592650 694926
rect -8726 694658 -3894 694894
rect -3658 694658 -3574 694894
rect -3338 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 587262 694894
rect 587498 694658 587582 694894
rect 587818 694658 592650 694894
rect -8726 694574 592650 694658
rect -8726 694338 -3894 694574
rect -3658 694338 -3574 694574
rect -3338 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 587262 694574
rect 587498 694338 587582 694574
rect 587818 694338 592650 694574
rect -8726 694306 592650 694338
rect -8726 691174 592650 691206
rect -8726 690938 -2934 691174
rect -2698 690938 -2614 691174
rect -2378 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 586302 691174
rect 586538 690938 586622 691174
rect 586858 690938 592650 691174
rect -8726 690854 592650 690938
rect -8726 690618 -2934 690854
rect -2698 690618 -2614 690854
rect -2378 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 586302 690854
rect 586538 690618 586622 690854
rect 586858 690618 592650 690854
rect -8726 690586 592650 690618
rect -8726 687454 592650 687486
rect -8726 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 592650 687454
rect -8726 687134 592650 687218
rect -8726 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 592650 687134
rect -8726 686866 592650 686898
rect -8726 677494 592650 677526
rect -8726 677258 -8694 677494
rect -8458 677258 -8374 677494
rect -8138 677258 27866 677494
rect 28102 677258 28186 677494
rect 28422 677258 63866 677494
rect 64102 677258 64186 677494
rect 64422 677258 99866 677494
rect 100102 677258 100186 677494
rect 100422 677258 135866 677494
rect 136102 677258 136186 677494
rect 136422 677258 171866 677494
rect 172102 677258 172186 677494
rect 172422 677258 207866 677494
rect 208102 677258 208186 677494
rect 208422 677258 243866 677494
rect 244102 677258 244186 677494
rect 244422 677258 279866 677494
rect 280102 677258 280186 677494
rect 280422 677258 315866 677494
rect 316102 677258 316186 677494
rect 316422 677258 351866 677494
rect 352102 677258 352186 677494
rect 352422 677258 387866 677494
rect 388102 677258 388186 677494
rect 388422 677258 423866 677494
rect 424102 677258 424186 677494
rect 424422 677258 459866 677494
rect 460102 677258 460186 677494
rect 460422 677258 495866 677494
rect 496102 677258 496186 677494
rect 496422 677258 531866 677494
rect 532102 677258 532186 677494
rect 532422 677258 567866 677494
rect 568102 677258 568186 677494
rect 568422 677258 592062 677494
rect 592298 677258 592382 677494
rect 592618 677258 592650 677494
rect -8726 677174 592650 677258
rect -8726 676938 -8694 677174
rect -8458 676938 -8374 677174
rect -8138 676938 27866 677174
rect 28102 676938 28186 677174
rect 28422 676938 63866 677174
rect 64102 676938 64186 677174
rect 64422 676938 99866 677174
rect 100102 676938 100186 677174
rect 100422 676938 135866 677174
rect 136102 676938 136186 677174
rect 136422 676938 171866 677174
rect 172102 676938 172186 677174
rect 172422 676938 207866 677174
rect 208102 676938 208186 677174
rect 208422 676938 243866 677174
rect 244102 676938 244186 677174
rect 244422 676938 279866 677174
rect 280102 676938 280186 677174
rect 280422 676938 315866 677174
rect 316102 676938 316186 677174
rect 316422 676938 351866 677174
rect 352102 676938 352186 677174
rect 352422 676938 387866 677174
rect 388102 676938 388186 677174
rect 388422 676938 423866 677174
rect 424102 676938 424186 677174
rect 424422 676938 459866 677174
rect 460102 676938 460186 677174
rect 460422 676938 495866 677174
rect 496102 676938 496186 677174
rect 496422 676938 531866 677174
rect 532102 676938 532186 677174
rect 532422 676938 567866 677174
rect 568102 676938 568186 677174
rect 568422 676938 592062 677174
rect 592298 676938 592382 677174
rect 592618 676938 592650 677174
rect -8726 676906 592650 676938
rect -8726 673774 592650 673806
rect -8726 673538 -7734 673774
rect -7498 673538 -7414 673774
rect -7178 673538 24146 673774
rect 24382 673538 24466 673774
rect 24702 673538 60146 673774
rect 60382 673538 60466 673774
rect 60702 673538 96146 673774
rect 96382 673538 96466 673774
rect 96702 673538 132146 673774
rect 132382 673538 132466 673774
rect 132702 673538 168146 673774
rect 168382 673538 168466 673774
rect 168702 673538 204146 673774
rect 204382 673538 204466 673774
rect 204702 673538 240146 673774
rect 240382 673538 240466 673774
rect 240702 673538 276146 673774
rect 276382 673538 276466 673774
rect 276702 673538 312146 673774
rect 312382 673538 312466 673774
rect 312702 673538 348146 673774
rect 348382 673538 348466 673774
rect 348702 673538 384146 673774
rect 384382 673538 384466 673774
rect 384702 673538 420146 673774
rect 420382 673538 420466 673774
rect 420702 673538 456146 673774
rect 456382 673538 456466 673774
rect 456702 673538 492146 673774
rect 492382 673538 492466 673774
rect 492702 673538 528146 673774
rect 528382 673538 528466 673774
rect 528702 673538 564146 673774
rect 564382 673538 564466 673774
rect 564702 673538 591102 673774
rect 591338 673538 591422 673774
rect 591658 673538 592650 673774
rect -8726 673454 592650 673538
rect -8726 673218 -7734 673454
rect -7498 673218 -7414 673454
rect -7178 673218 24146 673454
rect 24382 673218 24466 673454
rect 24702 673218 60146 673454
rect 60382 673218 60466 673454
rect 60702 673218 96146 673454
rect 96382 673218 96466 673454
rect 96702 673218 132146 673454
rect 132382 673218 132466 673454
rect 132702 673218 168146 673454
rect 168382 673218 168466 673454
rect 168702 673218 204146 673454
rect 204382 673218 204466 673454
rect 204702 673218 240146 673454
rect 240382 673218 240466 673454
rect 240702 673218 276146 673454
rect 276382 673218 276466 673454
rect 276702 673218 312146 673454
rect 312382 673218 312466 673454
rect 312702 673218 348146 673454
rect 348382 673218 348466 673454
rect 348702 673218 384146 673454
rect 384382 673218 384466 673454
rect 384702 673218 420146 673454
rect 420382 673218 420466 673454
rect 420702 673218 456146 673454
rect 456382 673218 456466 673454
rect 456702 673218 492146 673454
rect 492382 673218 492466 673454
rect 492702 673218 528146 673454
rect 528382 673218 528466 673454
rect 528702 673218 564146 673454
rect 564382 673218 564466 673454
rect 564702 673218 591102 673454
rect 591338 673218 591422 673454
rect 591658 673218 592650 673454
rect -8726 673186 592650 673218
rect -8726 670054 592650 670086
rect -8726 669818 -6774 670054
rect -6538 669818 -6454 670054
rect -6218 669818 20426 670054
rect 20662 669818 20746 670054
rect 20982 669818 56426 670054
rect 56662 669818 56746 670054
rect 56982 669818 92426 670054
rect 92662 669818 92746 670054
rect 92982 669818 128426 670054
rect 128662 669818 128746 670054
rect 128982 669818 164426 670054
rect 164662 669818 164746 670054
rect 164982 669818 200426 670054
rect 200662 669818 200746 670054
rect 200982 669818 236426 670054
rect 236662 669818 236746 670054
rect 236982 669818 272426 670054
rect 272662 669818 272746 670054
rect 272982 669818 308426 670054
rect 308662 669818 308746 670054
rect 308982 669818 344426 670054
rect 344662 669818 344746 670054
rect 344982 669818 380426 670054
rect 380662 669818 380746 670054
rect 380982 669818 416426 670054
rect 416662 669818 416746 670054
rect 416982 669818 452426 670054
rect 452662 669818 452746 670054
rect 452982 669818 488426 670054
rect 488662 669818 488746 670054
rect 488982 669818 524426 670054
rect 524662 669818 524746 670054
rect 524982 669818 560426 670054
rect 560662 669818 560746 670054
rect 560982 669818 590142 670054
rect 590378 669818 590462 670054
rect 590698 669818 592650 670054
rect -8726 669734 592650 669818
rect -8726 669498 -6774 669734
rect -6538 669498 -6454 669734
rect -6218 669498 20426 669734
rect 20662 669498 20746 669734
rect 20982 669498 56426 669734
rect 56662 669498 56746 669734
rect 56982 669498 92426 669734
rect 92662 669498 92746 669734
rect 92982 669498 128426 669734
rect 128662 669498 128746 669734
rect 128982 669498 164426 669734
rect 164662 669498 164746 669734
rect 164982 669498 200426 669734
rect 200662 669498 200746 669734
rect 200982 669498 236426 669734
rect 236662 669498 236746 669734
rect 236982 669498 272426 669734
rect 272662 669498 272746 669734
rect 272982 669498 308426 669734
rect 308662 669498 308746 669734
rect 308982 669498 344426 669734
rect 344662 669498 344746 669734
rect 344982 669498 380426 669734
rect 380662 669498 380746 669734
rect 380982 669498 416426 669734
rect 416662 669498 416746 669734
rect 416982 669498 452426 669734
rect 452662 669498 452746 669734
rect 452982 669498 488426 669734
rect 488662 669498 488746 669734
rect 488982 669498 524426 669734
rect 524662 669498 524746 669734
rect 524982 669498 560426 669734
rect 560662 669498 560746 669734
rect 560982 669498 590142 669734
rect 590378 669498 590462 669734
rect 590698 669498 592650 669734
rect -8726 669466 592650 669498
rect -8726 666334 592650 666366
rect -8726 666098 -5814 666334
rect -5578 666098 -5494 666334
rect -5258 666098 16706 666334
rect 16942 666098 17026 666334
rect 17262 666098 52706 666334
rect 52942 666098 53026 666334
rect 53262 666098 88706 666334
rect 88942 666098 89026 666334
rect 89262 666098 124706 666334
rect 124942 666098 125026 666334
rect 125262 666098 160706 666334
rect 160942 666098 161026 666334
rect 161262 666098 196706 666334
rect 196942 666098 197026 666334
rect 197262 666098 232706 666334
rect 232942 666098 233026 666334
rect 233262 666098 268706 666334
rect 268942 666098 269026 666334
rect 269262 666098 304706 666334
rect 304942 666098 305026 666334
rect 305262 666098 340706 666334
rect 340942 666098 341026 666334
rect 341262 666098 376706 666334
rect 376942 666098 377026 666334
rect 377262 666098 412706 666334
rect 412942 666098 413026 666334
rect 413262 666098 448706 666334
rect 448942 666098 449026 666334
rect 449262 666098 484706 666334
rect 484942 666098 485026 666334
rect 485262 666098 520706 666334
rect 520942 666098 521026 666334
rect 521262 666098 556706 666334
rect 556942 666098 557026 666334
rect 557262 666098 589182 666334
rect 589418 666098 589502 666334
rect 589738 666098 592650 666334
rect -8726 666014 592650 666098
rect -8726 665778 -5814 666014
rect -5578 665778 -5494 666014
rect -5258 665778 16706 666014
rect 16942 665778 17026 666014
rect 17262 665778 52706 666014
rect 52942 665778 53026 666014
rect 53262 665778 88706 666014
rect 88942 665778 89026 666014
rect 89262 665778 124706 666014
rect 124942 665778 125026 666014
rect 125262 665778 160706 666014
rect 160942 665778 161026 666014
rect 161262 665778 196706 666014
rect 196942 665778 197026 666014
rect 197262 665778 232706 666014
rect 232942 665778 233026 666014
rect 233262 665778 268706 666014
rect 268942 665778 269026 666014
rect 269262 665778 304706 666014
rect 304942 665778 305026 666014
rect 305262 665778 340706 666014
rect 340942 665778 341026 666014
rect 341262 665778 376706 666014
rect 376942 665778 377026 666014
rect 377262 665778 412706 666014
rect 412942 665778 413026 666014
rect 413262 665778 448706 666014
rect 448942 665778 449026 666014
rect 449262 665778 484706 666014
rect 484942 665778 485026 666014
rect 485262 665778 520706 666014
rect 520942 665778 521026 666014
rect 521262 665778 556706 666014
rect 556942 665778 557026 666014
rect 557262 665778 589182 666014
rect 589418 665778 589502 666014
rect 589738 665778 592650 666014
rect -8726 665746 592650 665778
rect -8726 662614 592650 662646
rect -8726 662378 -4854 662614
rect -4618 662378 -4534 662614
rect -4298 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 588222 662614
rect 588458 662378 588542 662614
rect 588778 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -4854 662294
rect -4618 662058 -4534 662294
rect -4298 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 588222 662294
rect 588458 662058 588542 662294
rect 588778 662058 592650 662294
rect -8726 662026 592650 662058
rect -8726 658894 592650 658926
rect -8726 658658 -3894 658894
rect -3658 658658 -3574 658894
rect -3338 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 587262 658894
rect 587498 658658 587582 658894
rect 587818 658658 592650 658894
rect -8726 658574 592650 658658
rect -8726 658338 -3894 658574
rect -3658 658338 -3574 658574
rect -3338 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 587262 658574
rect 587498 658338 587582 658574
rect 587818 658338 592650 658574
rect -8726 658306 592650 658338
rect -8726 655174 592650 655206
rect -8726 654938 -2934 655174
rect -2698 654938 -2614 655174
rect -2378 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 586302 655174
rect 586538 654938 586622 655174
rect 586858 654938 592650 655174
rect -8726 654854 592650 654938
rect -8726 654618 -2934 654854
rect -2698 654618 -2614 654854
rect -2378 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 586302 654854
rect 586538 654618 586622 654854
rect 586858 654618 592650 654854
rect -8726 654586 592650 654618
rect -8726 651454 592650 651486
rect -8726 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 494250 651454
rect 494486 651218 524970 651454
rect 525206 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 592650 651454
rect -8726 651134 592650 651218
rect -8726 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 494250 651134
rect 494486 650898 524970 651134
rect 525206 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 592650 651134
rect -8726 650866 592650 650898
rect -8726 641494 592650 641526
rect -8726 641258 -8694 641494
rect -8458 641258 -8374 641494
rect -8138 641258 27866 641494
rect 28102 641258 28186 641494
rect 28422 641258 63866 641494
rect 64102 641258 64186 641494
rect 64422 641258 99866 641494
rect 100102 641258 100186 641494
rect 100422 641258 135866 641494
rect 136102 641258 136186 641494
rect 136422 641258 171866 641494
rect 172102 641258 172186 641494
rect 172422 641258 207866 641494
rect 208102 641258 208186 641494
rect 208422 641258 243866 641494
rect 244102 641258 244186 641494
rect 244422 641258 279866 641494
rect 280102 641258 280186 641494
rect 280422 641258 315866 641494
rect 316102 641258 316186 641494
rect 316422 641258 351866 641494
rect 352102 641258 352186 641494
rect 352422 641258 387866 641494
rect 388102 641258 388186 641494
rect 388422 641258 423866 641494
rect 424102 641258 424186 641494
rect 424422 641258 459866 641494
rect 460102 641258 460186 641494
rect 460422 641258 567866 641494
rect 568102 641258 568186 641494
rect 568422 641258 592062 641494
rect 592298 641258 592382 641494
rect 592618 641258 592650 641494
rect -8726 641174 592650 641258
rect -8726 640938 -8694 641174
rect -8458 640938 -8374 641174
rect -8138 640938 27866 641174
rect 28102 640938 28186 641174
rect 28422 640938 63866 641174
rect 64102 640938 64186 641174
rect 64422 640938 99866 641174
rect 100102 640938 100186 641174
rect 100422 640938 135866 641174
rect 136102 640938 136186 641174
rect 136422 640938 171866 641174
rect 172102 640938 172186 641174
rect 172422 640938 207866 641174
rect 208102 640938 208186 641174
rect 208422 640938 243866 641174
rect 244102 640938 244186 641174
rect 244422 640938 279866 641174
rect 280102 640938 280186 641174
rect 280422 640938 315866 641174
rect 316102 640938 316186 641174
rect 316422 640938 351866 641174
rect 352102 640938 352186 641174
rect 352422 640938 387866 641174
rect 388102 640938 388186 641174
rect 388422 640938 423866 641174
rect 424102 640938 424186 641174
rect 424422 640938 459866 641174
rect 460102 640938 460186 641174
rect 460422 640938 567866 641174
rect 568102 640938 568186 641174
rect 568422 640938 592062 641174
rect 592298 640938 592382 641174
rect 592618 640938 592650 641174
rect -8726 640906 592650 640938
rect -8726 637774 592650 637806
rect -8726 637538 -7734 637774
rect -7498 637538 -7414 637774
rect -7178 637538 24146 637774
rect 24382 637538 24466 637774
rect 24702 637538 60146 637774
rect 60382 637538 60466 637774
rect 60702 637538 96146 637774
rect 96382 637538 96466 637774
rect 96702 637538 132146 637774
rect 132382 637538 132466 637774
rect 132702 637538 168146 637774
rect 168382 637538 168466 637774
rect 168702 637538 204146 637774
rect 204382 637538 204466 637774
rect 204702 637538 240146 637774
rect 240382 637538 240466 637774
rect 240702 637538 276146 637774
rect 276382 637538 276466 637774
rect 276702 637538 312146 637774
rect 312382 637538 312466 637774
rect 312702 637538 348146 637774
rect 348382 637538 348466 637774
rect 348702 637538 384146 637774
rect 384382 637538 384466 637774
rect 384702 637538 420146 637774
rect 420382 637538 420466 637774
rect 420702 637538 456146 637774
rect 456382 637538 456466 637774
rect 456702 637538 492146 637774
rect 492382 637538 492466 637774
rect 492702 637538 564146 637774
rect 564382 637538 564466 637774
rect 564702 637538 591102 637774
rect 591338 637538 591422 637774
rect 591658 637538 592650 637774
rect -8726 637454 592650 637538
rect -8726 637218 -7734 637454
rect -7498 637218 -7414 637454
rect -7178 637218 24146 637454
rect 24382 637218 24466 637454
rect 24702 637218 60146 637454
rect 60382 637218 60466 637454
rect 60702 637218 96146 637454
rect 96382 637218 96466 637454
rect 96702 637218 132146 637454
rect 132382 637218 132466 637454
rect 132702 637218 168146 637454
rect 168382 637218 168466 637454
rect 168702 637218 204146 637454
rect 204382 637218 204466 637454
rect 204702 637218 240146 637454
rect 240382 637218 240466 637454
rect 240702 637218 276146 637454
rect 276382 637218 276466 637454
rect 276702 637218 312146 637454
rect 312382 637218 312466 637454
rect 312702 637218 348146 637454
rect 348382 637218 348466 637454
rect 348702 637218 384146 637454
rect 384382 637218 384466 637454
rect 384702 637218 420146 637454
rect 420382 637218 420466 637454
rect 420702 637218 456146 637454
rect 456382 637218 456466 637454
rect 456702 637218 492146 637454
rect 492382 637218 492466 637454
rect 492702 637218 564146 637454
rect 564382 637218 564466 637454
rect 564702 637218 591102 637454
rect 591338 637218 591422 637454
rect 591658 637218 592650 637454
rect -8726 637186 592650 637218
rect -8726 634054 592650 634086
rect -8726 633818 -6774 634054
rect -6538 633818 -6454 634054
rect -6218 633818 20426 634054
rect 20662 633818 20746 634054
rect 20982 633818 56426 634054
rect 56662 633818 56746 634054
rect 56982 633818 92426 634054
rect 92662 633818 92746 634054
rect 92982 633818 128426 634054
rect 128662 633818 128746 634054
rect 128982 633818 164426 634054
rect 164662 633818 164746 634054
rect 164982 633818 200426 634054
rect 200662 633818 200746 634054
rect 200982 633818 236426 634054
rect 236662 633818 236746 634054
rect 236982 633818 272426 634054
rect 272662 633818 272746 634054
rect 272982 633818 308426 634054
rect 308662 633818 308746 634054
rect 308982 633818 344426 634054
rect 344662 633818 344746 634054
rect 344982 633818 380426 634054
rect 380662 633818 380746 634054
rect 380982 633818 416426 634054
rect 416662 633818 416746 634054
rect 416982 633818 452426 634054
rect 452662 633818 452746 634054
rect 452982 633818 488426 634054
rect 488662 633818 488746 634054
rect 488982 633818 560426 634054
rect 560662 633818 560746 634054
rect 560982 633818 590142 634054
rect 590378 633818 590462 634054
rect 590698 633818 592650 634054
rect -8726 633734 592650 633818
rect -8726 633498 -6774 633734
rect -6538 633498 -6454 633734
rect -6218 633498 20426 633734
rect 20662 633498 20746 633734
rect 20982 633498 56426 633734
rect 56662 633498 56746 633734
rect 56982 633498 92426 633734
rect 92662 633498 92746 633734
rect 92982 633498 128426 633734
rect 128662 633498 128746 633734
rect 128982 633498 164426 633734
rect 164662 633498 164746 633734
rect 164982 633498 200426 633734
rect 200662 633498 200746 633734
rect 200982 633498 236426 633734
rect 236662 633498 236746 633734
rect 236982 633498 272426 633734
rect 272662 633498 272746 633734
rect 272982 633498 308426 633734
rect 308662 633498 308746 633734
rect 308982 633498 344426 633734
rect 344662 633498 344746 633734
rect 344982 633498 380426 633734
rect 380662 633498 380746 633734
rect 380982 633498 416426 633734
rect 416662 633498 416746 633734
rect 416982 633498 452426 633734
rect 452662 633498 452746 633734
rect 452982 633498 488426 633734
rect 488662 633498 488746 633734
rect 488982 633498 560426 633734
rect 560662 633498 560746 633734
rect 560982 633498 590142 633734
rect 590378 633498 590462 633734
rect 590698 633498 592650 633734
rect -8726 633466 592650 633498
rect -8726 630334 592650 630366
rect -8726 630098 -5814 630334
rect -5578 630098 -5494 630334
rect -5258 630098 16706 630334
rect 16942 630098 17026 630334
rect 17262 630098 52706 630334
rect 52942 630098 53026 630334
rect 53262 630098 160706 630334
rect 160942 630098 161026 630334
rect 161262 630098 268706 630334
rect 268942 630098 269026 630334
rect 269262 630098 376706 630334
rect 376942 630098 377026 630334
rect 377262 630098 412706 630334
rect 412942 630098 413026 630334
rect 413262 630098 448706 630334
rect 448942 630098 449026 630334
rect 449262 630098 484706 630334
rect 484942 630098 485026 630334
rect 485262 630098 556706 630334
rect 556942 630098 557026 630334
rect 557262 630098 589182 630334
rect 589418 630098 589502 630334
rect 589738 630098 592650 630334
rect -8726 630014 592650 630098
rect -8726 629778 -5814 630014
rect -5578 629778 -5494 630014
rect -5258 629778 16706 630014
rect 16942 629778 17026 630014
rect 17262 629778 52706 630014
rect 52942 629778 53026 630014
rect 53262 629778 160706 630014
rect 160942 629778 161026 630014
rect 161262 629778 268706 630014
rect 268942 629778 269026 630014
rect 269262 629778 376706 630014
rect 376942 629778 377026 630014
rect 377262 629778 412706 630014
rect 412942 629778 413026 630014
rect 413262 629778 448706 630014
rect 448942 629778 449026 630014
rect 449262 629778 484706 630014
rect 484942 629778 485026 630014
rect 485262 629778 556706 630014
rect 556942 629778 557026 630014
rect 557262 629778 589182 630014
rect 589418 629778 589502 630014
rect 589738 629778 592650 630014
rect -8726 629746 592650 629778
rect -8726 626614 592650 626646
rect -8726 626378 -4854 626614
rect -4618 626378 -4534 626614
rect -4298 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 588222 626614
rect 588458 626378 588542 626614
rect 588778 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -4854 626294
rect -4618 626058 -4534 626294
rect -4298 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 588222 626294
rect 588458 626058 588542 626294
rect 588778 626058 592650 626294
rect -8726 626026 592650 626058
rect -8726 622894 592650 622926
rect -8726 622658 -3894 622894
rect -3658 622658 -3574 622894
rect -3338 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 587262 622894
rect 587498 622658 587582 622894
rect 587818 622658 592650 622894
rect -8726 622574 592650 622658
rect -8726 622338 -3894 622574
rect -3658 622338 -3574 622574
rect -3338 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 587262 622574
rect 587498 622338 587582 622574
rect 587818 622338 592650 622574
rect -8726 622306 592650 622338
rect -8726 619174 592650 619206
rect -8726 618938 -2934 619174
rect -2698 618938 -2614 619174
rect -2378 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 79610 619174
rect 79846 618938 110330 619174
rect 110566 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 199610 619174
rect 199846 618938 230330 619174
rect 230566 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 319610 619174
rect 319846 618938 350330 619174
rect 350566 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509610 619174
rect 509846 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 586302 619174
rect 586538 618938 586622 619174
rect 586858 618938 592650 619174
rect -8726 618854 592650 618938
rect -8726 618618 -2934 618854
rect -2698 618618 -2614 618854
rect -2378 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 79610 618854
rect 79846 618618 110330 618854
rect 110566 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 199610 618854
rect 199846 618618 230330 618854
rect 230566 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 319610 618854
rect 319846 618618 350330 618854
rect 350566 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509610 618854
rect 509846 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 586302 618854
rect 586538 618618 586622 618854
rect 586858 618618 592650 618854
rect -8726 618586 592650 618618
rect -8726 615454 592650 615486
rect -8726 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 125690 615454
rect 125926 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 184250 615454
rect 184486 615218 214970 615454
rect 215206 615218 245690 615454
rect 245926 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 304250 615454
rect 304486 615218 334970 615454
rect 335206 615218 365690 615454
rect 365926 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 494250 615454
rect 494486 615218 524970 615454
rect 525206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 592650 615454
rect -8726 615134 592650 615218
rect -8726 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 125690 615134
rect 125926 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 184250 615134
rect 184486 614898 214970 615134
rect 215206 614898 245690 615134
rect 245926 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 304250 615134
rect 304486 614898 334970 615134
rect 335206 614898 365690 615134
rect 365926 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 494250 615134
rect 494486 614898 524970 615134
rect 525206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 592650 615134
rect -8726 614866 592650 614898
rect -8726 605494 592650 605526
rect -8726 605258 -8694 605494
rect -8458 605258 -8374 605494
rect -8138 605258 27866 605494
rect 28102 605258 28186 605494
rect 28422 605258 135866 605494
rect 136102 605258 136186 605494
rect 136422 605258 171866 605494
rect 172102 605258 172186 605494
rect 172422 605258 279866 605494
rect 280102 605258 280186 605494
rect 280422 605258 387866 605494
rect 388102 605258 388186 605494
rect 388422 605258 423866 605494
rect 424102 605258 424186 605494
rect 424422 605258 459866 605494
rect 460102 605258 460186 605494
rect 460422 605258 567866 605494
rect 568102 605258 568186 605494
rect 568422 605258 592062 605494
rect 592298 605258 592382 605494
rect 592618 605258 592650 605494
rect -8726 605174 592650 605258
rect -8726 604938 -8694 605174
rect -8458 604938 -8374 605174
rect -8138 604938 27866 605174
rect 28102 604938 28186 605174
rect 28422 604938 135866 605174
rect 136102 604938 136186 605174
rect 136422 604938 171866 605174
rect 172102 604938 172186 605174
rect 172422 604938 279866 605174
rect 280102 604938 280186 605174
rect 280422 604938 387866 605174
rect 388102 604938 388186 605174
rect 388422 604938 423866 605174
rect 424102 604938 424186 605174
rect 424422 604938 459866 605174
rect 460102 604938 460186 605174
rect 460422 604938 567866 605174
rect 568102 604938 568186 605174
rect 568422 604938 592062 605174
rect 592298 604938 592382 605174
rect 592618 604938 592650 605174
rect -8726 604906 592650 604938
rect -8726 601774 592650 601806
rect -8726 601538 -7734 601774
rect -7498 601538 -7414 601774
rect -7178 601538 24146 601774
rect 24382 601538 24466 601774
rect 24702 601538 168146 601774
rect 168382 601538 168466 601774
rect 168702 601538 276146 601774
rect 276382 601538 276466 601774
rect 276702 601538 384146 601774
rect 384382 601538 384466 601774
rect 384702 601538 420146 601774
rect 420382 601538 420466 601774
rect 420702 601538 456146 601774
rect 456382 601538 456466 601774
rect 456702 601538 492146 601774
rect 492382 601538 492466 601774
rect 492702 601538 564146 601774
rect 564382 601538 564466 601774
rect 564702 601538 591102 601774
rect 591338 601538 591422 601774
rect 591658 601538 592650 601774
rect -8726 601454 592650 601538
rect -8726 601218 -7734 601454
rect -7498 601218 -7414 601454
rect -7178 601218 24146 601454
rect 24382 601218 24466 601454
rect 24702 601218 168146 601454
rect 168382 601218 168466 601454
rect 168702 601218 276146 601454
rect 276382 601218 276466 601454
rect 276702 601218 384146 601454
rect 384382 601218 384466 601454
rect 384702 601218 420146 601454
rect 420382 601218 420466 601454
rect 420702 601218 456146 601454
rect 456382 601218 456466 601454
rect 456702 601218 492146 601454
rect 492382 601218 492466 601454
rect 492702 601218 564146 601454
rect 564382 601218 564466 601454
rect 564702 601218 591102 601454
rect 591338 601218 591422 601454
rect 591658 601218 592650 601454
rect -8726 601186 592650 601218
rect -8726 598054 592650 598086
rect -8726 597818 -6774 598054
rect -6538 597818 -6454 598054
rect -6218 597818 20426 598054
rect 20662 597818 20746 598054
rect 20982 597818 56426 598054
rect 56662 597818 56746 598054
rect 56982 597818 164426 598054
rect 164662 597818 164746 598054
rect 164982 597818 272426 598054
rect 272662 597818 272746 598054
rect 272982 597818 380426 598054
rect 380662 597818 380746 598054
rect 380982 597818 416426 598054
rect 416662 597818 416746 598054
rect 416982 597818 452426 598054
rect 452662 597818 452746 598054
rect 452982 597818 488426 598054
rect 488662 597818 488746 598054
rect 488982 597818 524426 598054
rect 524662 597818 524746 598054
rect 524982 597818 560426 598054
rect 560662 597818 560746 598054
rect 560982 597818 590142 598054
rect 590378 597818 590462 598054
rect 590698 597818 592650 598054
rect -8726 597734 592650 597818
rect -8726 597498 -6774 597734
rect -6538 597498 -6454 597734
rect -6218 597498 20426 597734
rect 20662 597498 20746 597734
rect 20982 597498 56426 597734
rect 56662 597498 56746 597734
rect 56982 597498 164426 597734
rect 164662 597498 164746 597734
rect 164982 597498 272426 597734
rect 272662 597498 272746 597734
rect 272982 597498 380426 597734
rect 380662 597498 380746 597734
rect 380982 597498 416426 597734
rect 416662 597498 416746 597734
rect 416982 597498 452426 597734
rect 452662 597498 452746 597734
rect 452982 597498 488426 597734
rect 488662 597498 488746 597734
rect 488982 597498 524426 597734
rect 524662 597498 524746 597734
rect 524982 597498 560426 597734
rect 560662 597498 560746 597734
rect 560982 597498 590142 597734
rect 590378 597498 590462 597734
rect 590698 597498 592650 597734
rect -8726 597466 592650 597498
rect -8726 594334 592650 594366
rect -8726 594098 -5814 594334
rect -5578 594098 -5494 594334
rect -5258 594098 16706 594334
rect 16942 594098 17026 594334
rect 17262 594098 52706 594334
rect 52942 594098 53026 594334
rect 53262 594098 160706 594334
rect 160942 594098 161026 594334
rect 161262 594098 268706 594334
rect 268942 594098 269026 594334
rect 269262 594098 376706 594334
rect 376942 594098 377026 594334
rect 377262 594098 412706 594334
rect 412942 594098 413026 594334
rect 413262 594098 448706 594334
rect 448942 594098 449026 594334
rect 449262 594098 484706 594334
rect 484942 594098 485026 594334
rect 485262 594098 520706 594334
rect 520942 594098 521026 594334
rect 521262 594098 556706 594334
rect 556942 594098 557026 594334
rect 557262 594098 589182 594334
rect 589418 594098 589502 594334
rect 589738 594098 592650 594334
rect -8726 594014 592650 594098
rect -8726 593778 -5814 594014
rect -5578 593778 -5494 594014
rect -5258 593778 16706 594014
rect 16942 593778 17026 594014
rect 17262 593778 52706 594014
rect 52942 593778 53026 594014
rect 53262 593778 160706 594014
rect 160942 593778 161026 594014
rect 161262 593778 268706 594014
rect 268942 593778 269026 594014
rect 269262 593778 376706 594014
rect 376942 593778 377026 594014
rect 377262 593778 412706 594014
rect 412942 593778 413026 594014
rect 413262 593778 448706 594014
rect 448942 593778 449026 594014
rect 449262 593778 484706 594014
rect 484942 593778 485026 594014
rect 485262 593778 520706 594014
rect 520942 593778 521026 594014
rect 521262 593778 556706 594014
rect 556942 593778 557026 594014
rect 557262 593778 589182 594014
rect 589418 593778 589502 594014
rect 589738 593778 592650 594014
rect -8726 593746 592650 593778
rect -8726 590614 592650 590646
rect -8726 590378 -4854 590614
rect -4618 590378 -4534 590614
rect -4298 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 588222 590614
rect 588458 590378 588542 590614
rect 588778 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -4854 590294
rect -4618 590058 -4534 590294
rect -4298 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 588222 590294
rect 588458 590058 588542 590294
rect 588778 590058 592650 590294
rect -8726 590026 592650 590058
rect -8726 586894 592650 586926
rect -8726 586658 -3894 586894
rect -3658 586658 -3574 586894
rect -3338 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 587262 586894
rect 587498 586658 587582 586894
rect 587818 586658 592650 586894
rect -8726 586574 592650 586658
rect -8726 586338 -3894 586574
rect -3658 586338 -3574 586574
rect -3338 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 587262 586574
rect 587498 586338 587582 586574
rect 587818 586338 592650 586574
rect -8726 586306 592650 586338
rect -8726 583174 592650 583206
rect -8726 582938 -2934 583174
rect -2698 582938 -2614 583174
rect -2378 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 79610 583174
rect 79846 582938 110330 583174
rect 110566 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 199610 583174
rect 199846 582938 230330 583174
rect 230566 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 319610 583174
rect 319846 582938 350330 583174
rect 350566 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 586302 583174
rect 586538 582938 586622 583174
rect 586858 582938 592650 583174
rect -8726 582854 592650 582938
rect -8726 582618 -2934 582854
rect -2698 582618 -2614 582854
rect -2378 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 79610 582854
rect 79846 582618 110330 582854
rect 110566 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 199610 582854
rect 199846 582618 230330 582854
rect 230566 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 319610 582854
rect 319846 582618 350330 582854
rect 350566 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 586302 582854
rect 586538 582618 586622 582854
rect 586858 582618 592650 582854
rect -8726 582586 592650 582618
rect -8726 579454 592650 579486
rect -8726 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64250 579454
rect 64486 579218 94970 579454
rect 95206 579218 125690 579454
rect 125926 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 184250 579454
rect 184486 579218 214970 579454
rect 215206 579218 245690 579454
rect 245926 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 304250 579454
rect 304486 579218 334970 579454
rect 335206 579218 365690 579454
rect 365926 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 592650 579454
rect -8726 579134 592650 579218
rect -8726 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64250 579134
rect 64486 578898 94970 579134
rect 95206 578898 125690 579134
rect 125926 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 184250 579134
rect 184486 578898 214970 579134
rect 215206 578898 245690 579134
rect 245926 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 304250 579134
rect 304486 578898 334970 579134
rect 335206 578898 365690 579134
rect 365926 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 592650 579134
rect -8726 578866 592650 578898
rect -8726 569494 592650 569526
rect -8726 569258 -8694 569494
rect -8458 569258 -8374 569494
rect -8138 569258 27866 569494
rect 28102 569258 28186 569494
rect 28422 569258 135866 569494
rect 136102 569258 136186 569494
rect 136422 569258 171866 569494
rect 172102 569258 172186 569494
rect 172422 569258 279866 569494
rect 280102 569258 280186 569494
rect 280422 569258 387866 569494
rect 388102 569258 388186 569494
rect 388422 569258 423866 569494
rect 424102 569258 424186 569494
rect 424422 569258 459866 569494
rect 460102 569258 460186 569494
rect 460422 569258 495866 569494
rect 496102 569258 496186 569494
rect 496422 569258 531866 569494
rect 532102 569258 532186 569494
rect 532422 569258 567866 569494
rect 568102 569258 568186 569494
rect 568422 569258 592062 569494
rect 592298 569258 592382 569494
rect 592618 569258 592650 569494
rect -8726 569174 592650 569258
rect -8726 568938 -8694 569174
rect -8458 568938 -8374 569174
rect -8138 568938 27866 569174
rect 28102 568938 28186 569174
rect 28422 568938 135866 569174
rect 136102 568938 136186 569174
rect 136422 568938 171866 569174
rect 172102 568938 172186 569174
rect 172422 568938 279866 569174
rect 280102 568938 280186 569174
rect 280422 568938 387866 569174
rect 388102 568938 388186 569174
rect 388422 568938 423866 569174
rect 424102 568938 424186 569174
rect 424422 568938 459866 569174
rect 460102 568938 460186 569174
rect 460422 568938 495866 569174
rect 496102 568938 496186 569174
rect 496422 568938 531866 569174
rect 532102 568938 532186 569174
rect 532422 568938 567866 569174
rect 568102 568938 568186 569174
rect 568422 568938 592062 569174
rect 592298 568938 592382 569174
rect 592618 568938 592650 569174
rect -8726 568906 592650 568938
rect -8726 565774 592650 565806
rect -8726 565538 -7734 565774
rect -7498 565538 -7414 565774
rect -7178 565538 24146 565774
rect 24382 565538 24466 565774
rect 24702 565538 168146 565774
rect 168382 565538 168466 565774
rect 168702 565538 276146 565774
rect 276382 565538 276466 565774
rect 276702 565538 384146 565774
rect 384382 565538 384466 565774
rect 384702 565538 420146 565774
rect 420382 565538 420466 565774
rect 420702 565538 456146 565774
rect 456382 565538 456466 565774
rect 456702 565538 492146 565774
rect 492382 565538 492466 565774
rect 492702 565538 528146 565774
rect 528382 565538 528466 565774
rect 528702 565538 564146 565774
rect 564382 565538 564466 565774
rect 564702 565538 591102 565774
rect 591338 565538 591422 565774
rect 591658 565538 592650 565774
rect -8726 565454 592650 565538
rect -8726 565218 -7734 565454
rect -7498 565218 -7414 565454
rect -7178 565218 24146 565454
rect 24382 565218 24466 565454
rect 24702 565218 168146 565454
rect 168382 565218 168466 565454
rect 168702 565218 276146 565454
rect 276382 565218 276466 565454
rect 276702 565218 384146 565454
rect 384382 565218 384466 565454
rect 384702 565218 420146 565454
rect 420382 565218 420466 565454
rect 420702 565218 456146 565454
rect 456382 565218 456466 565454
rect 456702 565218 492146 565454
rect 492382 565218 492466 565454
rect 492702 565218 528146 565454
rect 528382 565218 528466 565454
rect 528702 565218 564146 565454
rect 564382 565218 564466 565454
rect 564702 565218 591102 565454
rect 591338 565218 591422 565454
rect 591658 565218 592650 565454
rect -8726 565186 592650 565218
rect -8726 562054 592650 562086
rect -8726 561818 -6774 562054
rect -6538 561818 -6454 562054
rect -6218 561818 20426 562054
rect 20662 561818 20746 562054
rect 20982 561818 56426 562054
rect 56662 561818 56746 562054
rect 56982 561818 164426 562054
rect 164662 561818 164746 562054
rect 164982 561818 272426 562054
rect 272662 561818 272746 562054
rect 272982 561818 380426 562054
rect 380662 561818 380746 562054
rect 380982 561818 416426 562054
rect 416662 561818 416746 562054
rect 416982 561818 452426 562054
rect 452662 561818 452746 562054
rect 452982 561818 488426 562054
rect 488662 561818 488746 562054
rect 488982 561818 524426 562054
rect 524662 561818 524746 562054
rect 524982 561818 560426 562054
rect 560662 561818 560746 562054
rect 560982 561818 590142 562054
rect 590378 561818 590462 562054
rect 590698 561818 592650 562054
rect -8726 561734 592650 561818
rect -8726 561498 -6774 561734
rect -6538 561498 -6454 561734
rect -6218 561498 20426 561734
rect 20662 561498 20746 561734
rect 20982 561498 56426 561734
rect 56662 561498 56746 561734
rect 56982 561498 164426 561734
rect 164662 561498 164746 561734
rect 164982 561498 272426 561734
rect 272662 561498 272746 561734
rect 272982 561498 380426 561734
rect 380662 561498 380746 561734
rect 380982 561498 416426 561734
rect 416662 561498 416746 561734
rect 416982 561498 452426 561734
rect 452662 561498 452746 561734
rect 452982 561498 488426 561734
rect 488662 561498 488746 561734
rect 488982 561498 524426 561734
rect 524662 561498 524746 561734
rect 524982 561498 560426 561734
rect 560662 561498 560746 561734
rect 560982 561498 590142 561734
rect 590378 561498 590462 561734
rect 590698 561498 592650 561734
rect -8726 561466 592650 561498
rect -8726 558334 592650 558366
rect -8726 558098 -5814 558334
rect -5578 558098 -5494 558334
rect -5258 558098 16706 558334
rect 16942 558098 17026 558334
rect 17262 558098 52706 558334
rect 52942 558098 53026 558334
rect 53262 558098 88706 558334
rect 88942 558098 89026 558334
rect 89262 558098 124706 558334
rect 124942 558098 125026 558334
rect 125262 558098 160706 558334
rect 160942 558098 161026 558334
rect 161262 558098 196706 558334
rect 196942 558098 197026 558334
rect 197262 558098 232706 558334
rect 232942 558098 233026 558334
rect 233262 558098 268706 558334
rect 268942 558098 269026 558334
rect 269262 558098 304706 558334
rect 304942 558098 305026 558334
rect 305262 558098 340706 558334
rect 340942 558098 341026 558334
rect 341262 558098 376706 558334
rect 376942 558098 377026 558334
rect 377262 558098 412706 558334
rect 412942 558098 413026 558334
rect 413262 558098 448706 558334
rect 448942 558098 449026 558334
rect 449262 558098 484706 558334
rect 484942 558098 485026 558334
rect 485262 558098 520706 558334
rect 520942 558098 521026 558334
rect 521262 558098 556706 558334
rect 556942 558098 557026 558334
rect 557262 558098 589182 558334
rect 589418 558098 589502 558334
rect 589738 558098 592650 558334
rect -8726 558014 592650 558098
rect -8726 557778 -5814 558014
rect -5578 557778 -5494 558014
rect -5258 557778 16706 558014
rect 16942 557778 17026 558014
rect 17262 557778 52706 558014
rect 52942 557778 53026 558014
rect 53262 557778 88706 558014
rect 88942 557778 89026 558014
rect 89262 557778 124706 558014
rect 124942 557778 125026 558014
rect 125262 557778 160706 558014
rect 160942 557778 161026 558014
rect 161262 557778 196706 558014
rect 196942 557778 197026 558014
rect 197262 557778 232706 558014
rect 232942 557778 233026 558014
rect 233262 557778 268706 558014
rect 268942 557778 269026 558014
rect 269262 557778 304706 558014
rect 304942 557778 305026 558014
rect 305262 557778 340706 558014
rect 340942 557778 341026 558014
rect 341262 557778 376706 558014
rect 376942 557778 377026 558014
rect 377262 557778 412706 558014
rect 412942 557778 413026 558014
rect 413262 557778 448706 558014
rect 448942 557778 449026 558014
rect 449262 557778 484706 558014
rect 484942 557778 485026 558014
rect 485262 557778 520706 558014
rect 520942 557778 521026 558014
rect 521262 557778 556706 558014
rect 556942 557778 557026 558014
rect 557262 557778 589182 558014
rect 589418 557778 589502 558014
rect 589738 557778 592650 558014
rect -8726 557746 592650 557778
rect -8726 554614 592650 554646
rect -8726 554378 -4854 554614
rect -4618 554378 -4534 554614
rect -4298 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 588222 554614
rect 588458 554378 588542 554614
rect 588778 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -4854 554294
rect -4618 554058 -4534 554294
rect -4298 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 588222 554294
rect 588458 554058 588542 554294
rect 588778 554058 592650 554294
rect -8726 554026 592650 554058
rect -8726 550894 592650 550926
rect -8726 550658 -3894 550894
rect -3658 550658 -3574 550894
rect -3338 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 587262 550894
rect 587498 550658 587582 550894
rect 587818 550658 592650 550894
rect -8726 550574 592650 550658
rect -8726 550338 -3894 550574
rect -3658 550338 -3574 550574
rect -3338 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 587262 550574
rect 587498 550338 587582 550574
rect 587818 550338 592650 550574
rect -8726 550306 592650 550338
rect -8726 547174 592650 547206
rect -8726 546938 -2934 547174
rect -2698 546938 -2614 547174
rect -2378 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 586302 547174
rect 586538 546938 586622 547174
rect 586858 546938 592650 547174
rect -8726 546854 592650 546938
rect -8726 546618 -2934 546854
rect -2698 546618 -2614 546854
rect -2378 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 586302 546854
rect 586538 546618 586622 546854
rect 586858 546618 592650 546854
rect -8726 546586 592650 546618
rect -8726 543454 592650 543486
rect -8726 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 592650 543454
rect -8726 543134 592650 543218
rect -8726 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 592650 543134
rect -8726 542866 592650 542898
rect -8726 533494 592650 533526
rect -8726 533258 -8694 533494
rect -8458 533258 -8374 533494
rect -8138 533258 27866 533494
rect 28102 533258 28186 533494
rect 28422 533258 99866 533494
rect 100102 533258 100186 533494
rect 100422 533258 135866 533494
rect 136102 533258 136186 533494
rect 136422 533258 171866 533494
rect 172102 533258 172186 533494
rect 172422 533258 279866 533494
rect 280102 533258 280186 533494
rect 280422 533258 387866 533494
rect 388102 533258 388186 533494
rect 388422 533258 423866 533494
rect 424102 533258 424186 533494
rect 424422 533258 459866 533494
rect 460102 533258 460186 533494
rect 460422 533258 495866 533494
rect 496102 533258 496186 533494
rect 496422 533258 531866 533494
rect 532102 533258 532186 533494
rect 532422 533258 567866 533494
rect 568102 533258 568186 533494
rect 568422 533258 592062 533494
rect 592298 533258 592382 533494
rect 592618 533258 592650 533494
rect -8726 533174 592650 533258
rect -8726 532938 -8694 533174
rect -8458 532938 -8374 533174
rect -8138 532938 27866 533174
rect 28102 532938 28186 533174
rect 28422 532938 99866 533174
rect 100102 532938 100186 533174
rect 100422 532938 135866 533174
rect 136102 532938 136186 533174
rect 136422 532938 171866 533174
rect 172102 532938 172186 533174
rect 172422 532938 279866 533174
rect 280102 532938 280186 533174
rect 280422 532938 387866 533174
rect 388102 532938 388186 533174
rect 388422 532938 423866 533174
rect 424102 532938 424186 533174
rect 424422 532938 459866 533174
rect 460102 532938 460186 533174
rect 460422 532938 495866 533174
rect 496102 532938 496186 533174
rect 496422 532938 531866 533174
rect 532102 532938 532186 533174
rect 532422 532938 567866 533174
rect 568102 532938 568186 533174
rect 568422 532938 592062 533174
rect 592298 532938 592382 533174
rect 592618 532938 592650 533174
rect -8726 532906 592650 532938
rect -8726 529774 592650 529806
rect -8726 529538 -7734 529774
rect -7498 529538 -7414 529774
rect -7178 529538 24146 529774
rect 24382 529538 24466 529774
rect 24702 529538 60146 529774
rect 60382 529538 60466 529774
rect 60702 529538 96146 529774
rect 96382 529538 96466 529774
rect 96702 529538 132146 529774
rect 132382 529538 132466 529774
rect 132702 529538 168146 529774
rect 168382 529538 168466 529774
rect 168702 529538 276146 529774
rect 276382 529538 276466 529774
rect 276702 529538 384146 529774
rect 384382 529538 384466 529774
rect 384702 529538 420146 529774
rect 420382 529538 420466 529774
rect 420702 529538 456146 529774
rect 456382 529538 456466 529774
rect 456702 529538 492146 529774
rect 492382 529538 492466 529774
rect 492702 529538 528146 529774
rect 528382 529538 528466 529774
rect 528702 529538 564146 529774
rect 564382 529538 564466 529774
rect 564702 529538 591102 529774
rect 591338 529538 591422 529774
rect 591658 529538 592650 529774
rect -8726 529454 592650 529538
rect -8726 529218 -7734 529454
rect -7498 529218 -7414 529454
rect -7178 529218 24146 529454
rect 24382 529218 24466 529454
rect 24702 529218 60146 529454
rect 60382 529218 60466 529454
rect 60702 529218 96146 529454
rect 96382 529218 96466 529454
rect 96702 529218 132146 529454
rect 132382 529218 132466 529454
rect 132702 529218 168146 529454
rect 168382 529218 168466 529454
rect 168702 529218 276146 529454
rect 276382 529218 276466 529454
rect 276702 529218 384146 529454
rect 384382 529218 384466 529454
rect 384702 529218 420146 529454
rect 420382 529218 420466 529454
rect 420702 529218 456146 529454
rect 456382 529218 456466 529454
rect 456702 529218 492146 529454
rect 492382 529218 492466 529454
rect 492702 529218 528146 529454
rect 528382 529218 528466 529454
rect 528702 529218 564146 529454
rect 564382 529218 564466 529454
rect 564702 529218 591102 529454
rect 591338 529218 591422 529454
rect 591658 529218 592650 529454
rect -8726 529186 592650 529218
rect -8726 526054 592650 526086
rect -8726 525818 -6774 526054
rect -6538 525818 -6454 526054
rect -6218 525818 20426 526054
rect 20662 525818 20746 526054
rect 20982 525818 56426 526054
rect 56662 525818 56746 526054
rect 56982 525818 92426 526054
rect 92662 525818 92746 526054
rect 92982 525818 128426 526054
rect 128662 525818 128746 526054
rect 128982 525818 164426 526054
rect 164662 525818 164746 526054
rect 164982 525818 272426 526054
rect 272662 525818 272746 526054
rect 272982 525818 380426 526054
rect 380662 525818 380746 526054
rect 380982 525818 416426 526054
rect 416662 525818 416746 526054
rect 416982 525818 452426 526054
rect 452662 525818 452746 526054
rect 452982 525818 488426 526054
rect 488662 525818 488746 526054
rect 488982 525818 524426 526054
rect 524662 525818 524746 526054
rect 524982 525818 560426 526054
rect 560662 525818 560746 526054
rect 560982 525818 590142 526054
rect 590378 525818 590462 526054
rect 590698 525818 592650 526054
rect -8726 525734 592650 525818
rect -8726 525498 -6774 525734
rect -6538 525498 -6454 525734
rect -6218 525498 20426 525734
rect 20662 525498 20746 525734
rect 20982 525498 56426 525734
rect 56662 525498 56746 525734
rect 56982 525498 92426 525734
rect 92662 525498 92746 525734
rect 92982 525498 128426 525734
rect 128662 525498 128746 525734
rect 128982 525498 164426 525734
rect 164662 525498 164746 525734
rect 164982 525498 272426 525734
rect 272662 525498 272746 525734
rect 272982 525498 380426 525734
rect 380662 525498 380746 525734
rect 380982 525498 416426 525734
rect 416662 525498 416746 525734
rect 416982 525498 452426 525734
rect 452662 525498 452746 525734
rect 452982 525498 488426 525734
rect 488662 525498 488746 525734
rect 488982 525498 524426 525734
rect 524662 525498 524746 525734
rect 524982 525498 560426 525734
rect 560662 525498 560746 525734
rect 560982 525498 590142 525734
rect 590378 525498 590462 525734
rect 590698 525498 592650 525734
rect -8726 525466 592650 525498
rect -8726 522334 592650 522366
rect -8726 522098 -5814 522334
rect -5578 522098 -5494 522334
rect -5258 522098 16706 522334
rect 16942 522098 17026 522334
rect 17262 522098 52706 522334
rect 52942 522098 53026 522334
rect 53262 522098 88706 522334
rect 88942 522098 89026 522334
rect 89262 522098 124706 522334
rect 124942 522098 125026 522334
rect 125262 522098 160706 522334
rect 160942 522098 161026 522334
rect 161262 522098 196706 522334
rect 196942 522098 197026 522334
rect 197262 522098 520706 522334
rect 520942 522098 521026 522334
rect 521262 522098 556706 522334
rect 556942 522098 557026 522334
rect 557262 522098 589182 522334
rect 589418 522098 589502 522334
rect 589738 522098 592650 522334
rect -8726 522014 592650 522098
rect -8726 521778 -5814 522014
rect -5578 521778 -5494 522014
rect -5258 521778 16706 522014
rect 16942 521778 17026 522014
rect 17262 521778 52706 522014
rect 52942 521778 53026 522014
rect 53262 521778 88706 522014
rect 88942 521778 89026 522014
rect 89262 521778 124706 522014
rect 124942 521778 125026 522014
rect 125262 521778 160706 522014
rect 160942 521778 161026 522014
rect 161262 521778 196706 522014
rect 196942 521778 197026 522014
rect 197262 521778 520706 522014
rect 520942 521778 521026 522014
rect 521262 521778 556706 522014
rect 556942 521778 557026 522014
rect 557262 521778 589182 522014
rect 589418 521778 589502 522014
rect 589738 521778 592650 522014
rect -8726 521746 592650 521778
rect -8726 518614 592650 518646
rect -8726 518378 -4854 518614
rect -4618 518378 -4534 518614
rect -4298 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 588222 518614
rect 588458 518378 588542 518614
rect 588778 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -4854 518294
rect -4618 518058 -4534 518294
rect -4298 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 588222 518294
rect 588458 518058 588542 518294
rect 588778 518058 592650 518294
rect -8726 518026 592650 518058
rect -8726 514894 592650 514926
rect -8726 514658 -3894 514894
rect -3658 514658 -3574 514894
rect -3338 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 587262 514894
rect 587498 514658 587582 514894
rect 587818 514658 592650 514894
rect -8726 514574 592650 514658
rect -8726 514338 -3894 514574
rect -3658 514338 -3574 514574
rect -3338 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 587262 514574
rect 587498 514338 587582 514574
rect 587818 514338 592650 514574
rect -8726 514306 592650 514338
rect -8726 511174 592650 511206
rect -8726 510938 -2934 511174
rect -2698 510938 -2614 511174
rect -2378 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 79610 511174
rect 79846 510938 110330 511174
rect 110566 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 141050 511174
rect 141286 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 171770 511174
rect 172006 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 202490 511174
rect 202726 510938 233210 511174
rect 233446 510938 263930 511174
rect 264166 510938 294650 511174
rect 294886 510938 325370 511174
rect 325606 510938 356090 511174
rect 356326 510938 386810 511174
rect 387046 510938 417530 511174
rect 417766 510938 448250 511174
rect 448486 510938 478970 511174
rect 479206 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 586302 511174
rect 586538 510938 586622 511174
rect 586858 510938 592650 511174
rect -8726 510854 592650 510938
rect -8726 510618 -2934 510854
rect -2698 510618 -2614 510854
rect -2378 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 79610 510854
rect 79846 510618 110330 510854
rect 110566 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 141050 510854
rect 141286 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 171770 510854
rect 172006 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 202490 510854
rect 202726 510618 233210 510854
rect 233446 510618 263930 510854
rect 264166 510618 294650 510854
rect 294886 510618 325370 510854
rect 325606 510618 356090 510854
rect 356326 510618 386810 510854
rect 387046 510618 417530 510854
rect 417766 510618 448250 510854
rect 448486 510618 478970 510854
rect 479206 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 586302 510854
rect 586538 510618 586622 510854
rect 586858 510618 592650 510854
rect -8726 510586 592650 510618
rect -8726 507454 592650 507486
rect -8726 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 156410 507454
rect 156646 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 310010 507454
rect 310246 507218 340730 507454
rect 340966 507218 371450 507454
rect 371686 507218 402170 507454
rect 402406 507218 432890 507454
rect 433126 507218 463610 507454
rect 463846 507218 494330 507454
rect 494566 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 592650 507454
rect -8726 507134 592650 507218
rect -8726 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 156410 507134
rect 156646 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 310010 507134
rect 310246 506898 340730 507134
rect 340966 506898 371450 507134
rect 371686 506898 402170 507134
rect 402406 506898 432890 507134
rect 433126 506898 463610 507134
rect 463846 506898 494330 507134
rect 494566 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 592650 507134
rect -8726 506866 592650 506898
rect -8726 497494 592650 497526
rect -8726 497258 -8694 497494
rect -8458 497258 -8374 497494
rect -8138 497258 27866 497494
rect 28102 497258 28186 497494
rect 28422 497258 99866 497494
rect 100102 497258 100186 497494
rect 100422 497258 135866 497494
rect 136102 497258 136186 497494
rect 136422 497258 531866 497494
rect 532102 497258 532186 497494
rect 532422 497258 567866 497494
rect 568102 497258 568186 497494
rect 568422 497258 592062 497494
rect 592298 497258 592382 497494
rect 592618 497258 592650 497494
rect -8726 497174 592650 497258
rect -8726 496938 -8694 497174
rect -8458 496938 -8374 497174
rect -8138 496938 27866 497174
rect 28102 496938 28186 497174
rect 28422 496938 99866 497174
rect 100102 496938 100186 497174
rect 100422 496938 135866 497174
rect 136102 496938 136186 497174
rect 136422 496938 531866 497174
rect 532102 496938 532186 497174
rect 532422 496938 567866 497174
rect 568102 496938 568186 497174
rect 568422 496938 592062 497174
rect 592298 496938 592382 497174
rect 592618 496938 592650 497174
rect -8726 496906 592650 496938
rect -8726 493774 592650 493806
rect -8726 493538 -7734 493774
rect -7498 493538 -7414 493774
rect -7178 493538 24146 493774
rect 24382 493538 24466 493774
rect 24702 493538 60146 493774
rect 60382 493538 60466 493774
rect 60702 493538 96146 493774
rect 96382 493538 96466 493774
rect 96702 493538 132146 493774
rect 132382 493538 132466 493774
rect 132702 493538 168146 493774
rect 168382 493538 168466 493774
rect 168702 493538 528146 493774
rect 528382 493538 528466 493774
rect 528702 493538 564146 493774
rect 564382 493538 564466 493774
rect 564702 493538 591102 493774
rect 591338 493538 591422 493774
rect 591658 493538 592650 493774
rect -8726 493454 592650 493538
rect -8726 493218 -7734 493454
rect -7498 493218 -7414 493454
rect -7178 493218 24146 493454
rect 24382 493218 24466 493454
rect 24702 493218 60146 493454
rect 60382 493218 60466 493454
rect 60702 493218 96146 493454
rect 96382 493218 96466 493454
rect 96702 493218 132146 493454
rect 132382 493218 132466 493454
rect 132702 493218 168146 493454
rect 168382 493218 168466 493454
rect 168702 493218 528146 493454
rect 528382 493218 528466 493454
rect 528702 493218 564146 493454
rect 564382 493218 564466 493454
rect 564702 493218 591102 493454
rect 591338 493218 591422 493454
rect 591658 493218 592650 493454
rect -8726 493186 592650 493218
rect -8726 490054 592650 490086
rect -8726 489818 -6774 490054
rect -6538 489818 -6454 490054
rect -6218 489818 20426 490054
rect 20662 489818 20746 490054
rect 20982 489818 56426 490054
rect 56662 489818 56746 490054
rect 56982 489818 92426 490054
rect 92662 489818 92746 490054
rect 92982 489818 128426 490054
rect 128662 489818 128746 490054
rect 128982 489818 164426 490054
rect 164662 489818 164746 490054
rect 164982 489818 524426 490054
rect 524662 489818 524746 490054
rect 524982 489818 560426 490054
rect 560662 489818 560746 490054
rect 560982 489818 590142 490054
rect 590378 489818 590462 490054
rect 590698 489818 592650 490054
rect -8726 489734 592650 489818
rect -8726 489498 -6774 489734
rect -6538 489498 -6454 489734
rect -6218 489498 20426 489734
rect 20662 489498 20746 489734
rect 20982 489498 56426 489734
rect 56662 489498 56746 489734
rect 56982 489498 92426 489734
rect 92662 489498 92746 489734
rect 92982 489498 128426 489734
rect 128662 489498 128746 489734
rect 128982 489498 164426 489734
rect 164662 489498 164746 489734
rect 164982 489498 524426 489734
rect 524662 489498 524746 489734
rect 524982 489498 560426 489734
rect 560662 489498 560746 489734
rect 560982 489498 590142 489734
rect 590378 489498 590462 489734
rect 590698 489498 592650 489734
rect -8726 489466 592650 489498
rect -8726 486334 592650 486366
rect -8726 486098 -5814 486334
rect -5578 486098 -5494 486334
rect -5258 486098 16706 486334
rect 16942 486098 17026 486334
rect 17262 486098 52706 486334
rect 52942 486098 53026 486334
rect 53262 486098 88706 486334
rect 88942 486098 89026 486334
rect 89262 486098 124706 486334
rect 124942 486098 125026 486334
rect 125262 486098 160706 486334
rect 160942 486098 161026 486334
rect 161262 486098 196706 486334
rect 196942 486098 197026 486334
rect 197262 486098 520706 486334
rect 520942 486098 521026 486334
rect 521262 486098 556706 486334
rect 556942 486098 557026 486334
rect 557262 486098 589182 486334
rect 589418 486098 589502 486334
rect 589738 486098 592650 486334
rect -8726 486014 592650 486098
rect -8726 485778 -5814 486014
rect -5578 485778 -5494 486014
rect -5258 485778 16706 486014
rect 16942 485778 17026 486014
rect 17262 485778 52706 486014
rect 52942 485778 53026 486014
rect 53262 485778 88706 486014
rect 88942 485778 89026 486014
rect 89262 485778 124706 486014
rect 124942 485778 125026 486014
rect 125262 485778 160706 486014
rect 160942 485778 161026 486014
rect 161262 485778 196706 486014
rect 196942 485778 197026 486014
rect 197262 485778 520706 486014
rect 520942 485778 521026 486014
rect 521262 485778 556706 486014
rect 556942 485778 557026 486014
rect 557262 485778 589182 486014
rect 589418 485778 589502 486014
rect 589738 485778 592650 486014
rect -8726 485746 592650 485778
rect -8726 482614 592650 482646
rect -8726 482378 -4854 482614
rect -4618 482378 -4534 482614
rect -4298 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 588222 482614
rect 588458 482378 588542 482614
rect 588778 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -4854 482294
rect -4618 482058 -4534 482294
rect -4298 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 588222 482294
rect 588458 482058 588542 482294
rect 588778 482058 592650 482294
rect -8726 482026 592650 482058
rect -8726 478894 592650 478926
rect -8726 478658 -3894 478894
rect -3658 478658 -3574 478894
rect -3338 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 587262 478894
rect 587498 478658 587582 478894
rect 587818 478658 592650 478894
rect -8726 478574 592650 478658
rect -8726 478338 -3894 478574
rect -3658 478338 -3574 478574
rect -3338 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 587262 478574
rect 587498 478338 587582 478574
rect 587818 478338 592650 478574
rect -8726 478306 592650 478338
rect -8726 475174 592650 475206
rect -8726 474938 -2934 475174
rect -2698 474938 -2614 475174
rect -2378 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 79610 475174
rect 79846 474938 110330 475174
rect 110566 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 141050 475174
rect 141286 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 171770 475174
rect 172006 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 202490 475174
rect 202726 474938 233210 475174
rect 233446 474938 263930 475174
rect 264166 474938 294650 475174
rect 294886 474938 325370 475174
rect 325606 474938 356090 475174
rect 356326 474938 386810 475174
rect 387046 474938 417530 475174
rect 417766 474938 448250 475174
rect 448486 474938 478970 475174
rect 479206 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 586302 475174
rect 586538 474938 586622 475174
rect 586858 474938 592650 475174
rect -8726 474854 592650 474938
rect -8726 474618 -2934 474854
rect -2698 474618 -2614 474854
rect -2378 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 79610 474854
rect 79846 474618 110330 474854
rect 110566 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 141050 474854
rect 141286 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 171770 474854
rect 172006 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 202490 474854
rect 202726 474618 233210 474854
rect 233446 474618 263930 474854
rect 264166 474618 294650 474854
rect 294886 474618 325370 474854
rect 325606 474618 356090 474854
rect 356326 474618 386810 474854
rect 387046 474618 417530 474854
rect 417766 474618 448250 474854
rect 448486 474618 478970 474854
rect 479206 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 586302 474854
rect 586538 474618 586622 474854
rect 586858 474618 592650 474854
rect -8726 474586 592650 474618
rect -8726 471454 592650 471486
rect -8726 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 64250 471454
rect 64486 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 94970 471454
rect 95206 471218 125690 471454
rect 125926 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 156410 471454
rect 156646 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 187130 471454
rect 187366 471218 217850 471454
rect 218086 471218 248570 471454
rect 248806 471218 279290 471454
rect 279526 471218 310010 471454
rect 310246 471218 340730 471454
rect 340966 471218 371450 471454
rect 371686 471218 402170 471454
rect 402406 471218 432890 471454
rect 433126 471218 463610 471454
rect 463846 471218 494330 471454
rect 494566 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 592650 471454
rect -8726 471134 592650 471218
rect -8726 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 64250 471134
rect 64486 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 94970 471134
rect 95206 470898 125690 471134
rect 125926 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 156410 471134
rect 156646 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 187130 471134
rect 187366 470898 217850 471134
rect 218086 470898 248570 471134
rect 248806 470898 279290 471134
rect 279526 470898 310010 471134
rect 310246 470898 340730 471134
rect 340966 470898 371450 471134
rect 371686 470898 402170 471134
rect 402406 470898 432890 471134
rect 433126 470898 463610 471134
rect 463846 470898 494330 471134
rect 494566 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 592650 471134
rect -8726 470866 592650 470898
rect -8726 461494 592650 461526
rect -8726 461258 -8694 461494
rect -8458 461258 -8374 461494
rect -8138 461258 27866 461494
rect 28102 461258 28186 461494
rect 28422 461258 99866 461494
rect 100102 461258 100186 461494
rect 100422 461258 135866 461494
rect 136102 461258 136186 461494
rect 136422 461258 531866 461494
rect 532102 461258 532186 461494
rect 532422 461258 567866 461494
rect 568102 461258 568186 461494
rect 568422 461258 592062 461494
rect 592298 461258 592382 461494
rect 592618 461258 592650 461494
rect -8726 461174 592650 461258
rect -8726 460938 -8694 461174
rect -8458 460938 -8374 461174
rect -8138 460938 27866 461174
rect 28102 460938 28186 461174
rect 28422 460938 99866 461174
rect 100102 460938 100186 461174
rect 100422 460938 135866 461174
rect 136102 460938 136186 461174
rect 136422 460938 531866 461174
rect 532102 460938 532186 461174
rect 532422 460938 567866 461174
rect 568102 460938 568186 461174
rect 568422 460938 592062 461174
rect 592298 460938 592382 461174
rect 592618 460938 592650 461174
rect -8726 460906 592650 460938
rect -8726 457774 592650 457806
rect -8726 457538 -7734 457774
rect -7498 457538 -7414 457774
rect -7178 457538 24146 457774
rect 24382 457538 24466 457774
rect 24702 457538 60146 457774
rect 60382 457538 60466 457774
rect 60702 457538 96146 457774
rect 96382 457538 96466 457774
rect 96702 457538 132146 457774
rect 132382 457538 132466 457774
rect 132702 457538 168146 457774
rect 168382 457538 168466 457774
rect 168702 457538 528146 457774
rect 528382 457538 528466 457774
rect 528702 457538 564146 457774
rect 564382 457538 564466 457774
rect 564702 457538 591102 457774
rect 591338 457538 591422 457774
rect 591658 457538 592650 457774
rect -8726 457454 592650 457538
rect -8726 457218 -7734 457454
rect -7498 457218 -7414 457454
rect -7178 457218 24146 457454
rect 24382 457218 24466 457454
rect 24702 457218 60146 457454
rect 60382 457218 60466 457454
rect 60702 457218 96146 457454
rect 96382 457218 96466 457454
rect 96702 457218 132146 457454
rect 132382 457218 132466 457454
rect 132702 457218 168146 457454
rect 168382 457218 168466 457454
rect 168702 457218 528146 457454
rect 528382 457218 528466 457454
rect 528702 457218 564146 457454
rect 564382 457218 564466 457454
rect 564702 457218 591102 457454
rect 591338 457218 591422 457454
rect 591658 457218 592650 457454
rect -8726 457186 592650 457218
rect -8726 454054 592650 454086
rect -8726 453818 -6774 454054
rect -6538 453818 -6454 454054
rect -6218 453818 20426 454054
rect 20662 453818 20746 454054
rect 20982 453818 56426 454054
rect 56662 453818 56746 454054
rect 56982 453818 92426 454054
rect 92662 453818 92746 454054
rect 92982 453818 128426 454054
rect 128662 453818 128746 454054
rect 128982 453818 164426 454054
rect 164662 453818 164746 454054
rect 164982 453818 524426 454054
rect 524662 453818 524746 454054
rect 524982 453818 560426 454054
rect 560662 453818 560746 454054
rect 560982 453818 590142 454054
rect 590378 453818 590462 454054
rect 590698 453818 592650 454054
rect -8726 453734 592650 453818
rect -8726 453498 -6774 453734
rect -6538 453498 -6454 453734
rect -6218 453498 20426 453734
rect 20662 453498 20746 453734
rect 20982 453498 56426 453734
rect 56662 453498 56746 453734
rect 56982 453498 92426 453734
rect 92662 453498 92746 453734
rect 92982 453498 128426 453734
rect 128662 453498 128746 453734
rect 128982 453498 164426 453734
rect 164662 453498 164746 453734
rect 164982 453498 524426 453734
rect 524662 453498 524746 453734
rect 524982 453498 560426 453734
rect 560662 453498 560746 453734
rect 560982 453498 590142 453734
rect 590378 453498 590462 453734
rect 590698 453498 592650 453734
rect -8726 453466 592650 453498
rect -8726 450334 592650 450366
rect -8726 450098 -5814 450334
rect -5578 450098 -5494 450334
rect -5258 450098 16706 450334
rect 16942 450098 17026 450334
rect 17262 450098 52706 450334
rect 52942 450098 53026 450334
rect 53262 450098 88706 450334
rect 88942 450098 89026 450334
rect 89262 450098 124706 450334
rect 124942 450098 125026 450334
rect 125262 450098 160706 450334
rect 160942 450098 161026 450334
rect 161262 450098 196706 450334
rect 196942 450098 197026 450334
rect 197262 450098 520706 450334
rect 520942 450098 521026 450334
rect 521262 450098 556706 450334
rect 556942 450098 557026 450334
rect 557262 450098 589182 450334
rect 589418 450098 589502 450334
rect 589738 450098 592650 450334
rect -8726 450014 592650 450098
rect -8726 449778 -5814 450014
rect -5578 449778 -5494 450014
rect -5258 449778 16706 450014
rect 16942 449778 17026 450014
rect 17262 449778 52706 450014
rect 52942 449778 53026 450014
rect 53262 449778 88706 450014
rect 88942 449778 89026 450014
rect 89262 449778 124706 450014
rect 124942 449778 125026 450014
rect 125262 449778 160706 450014
rect 160942 449778 161026 450014
rect 161262 449778 196706 450014
rect 196942 449778 197026 450014
rect 197262 449778 520706 450014
rect 520942 449778 521026 450014
rect 521262 449778 556706 450014
rect 556942 449778 557026 450014
rect 557262 449778 589182 450014
rect 589418 449778 589502 450014
rect 589738 449778 592650 450014
rect -8726 449746 592650 449778
rect -8726 446614 592650 446646
rect -8726 446378 -4854 446614
rect -4618 446378 -4534 446614
rect -4298 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 84986 446614
rect 85222 446378 85306 446614
rect 85542 446378 120986 446614
rect 121222 446378 121306 446614
rect 121542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 588222 446614
rect 588458 446378 588542 446614
rect 588778 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -4854 446294
rect -4618 446058 -4534 446294
rect -4298 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 84986 446294
rect 85222 446058 85306 446294
rect 85542 446058 120986 446294
rect 121222 446058 121306 446294
rect 121542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 588222 446294
rect 588458 446058 588542 446294
rect 588778 446058 592650 446294
rect -8726 446026 592650 446058
rect -8726 442894 592650 442926
rect -8726 442658 -3894 442894
rect -3658 442658 -3574 442894
rect -3338 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 81266 442894
rect 81502 442658 81586 442894
rect 81822 442658 117266 442894
rect 117502 442658 117586 442894
rect 117822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 587262 442894
rect 587498 442658 587582 442894
rect 587818 442658 592650 442894
rect -8726 442574 592650 442658
rect -8726 442338 -3894 442574
rect -3658 442338 -3574 442574
rect -3338 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 81266 442574
rect 81502 442338 81586 442574
rect 81822 442338 117266 442574
rect 117502 442338 117586 442574
rect 117822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 587262 442574
rect 587498 442338 587582 442574
rect 587818 442338 592650 442574
rect -8726 442306 592650 442338
rect -8726 439174 592650 439206
rect -8726 438938 -2934 439174
rect -2698 438938 -2614 439174
rect -2378 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 77546 439174
rect 77782 438938 77866 439174
rect 78102 438938 79610 439174
rect 79846 438938 110330 439174
rect 110566 438938 113546 439174
rect 113782 438938 113866 439174
rect 114102 438938 141050 439174
rect 141286 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 171770 439174
rect 172006 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 202490 439174
rect 202726 438938 233210 439174
rect 233446 438938 263930 439174
rect 264166 438938 294650 439174
rect 294886 438938 325370 439174
rect 325606 438938 356090 439174
rect 356326 438938 386810 439174
rect 387046 438938 417530 439174
rect 417766 438938 448250 439174
rect 448486 438938 478970 439174
rect 479206 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 586302 439174
rect 586538 438938 586622 439174
rect 586858 438938 592650 439174
rect -8726 438854 592650 438938
rect -8726 438618 -2934 438854
rect -2698 438618 -2614 438854
rect -2378 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 77546 438854
rect 77782 438618 77866 438854
rect 78102 438618 79610 438854
rect 79846 438618 110330 438854
rect 110566 438618 113546 438854
rect 113782 438618 113866 438854
rect 114102 438618 141050 438854
rect 141286 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 171770 438854
rect 172006 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 202490 438854
rect 202726 438618 233210 438854
rect 233446 438618 263930 438854
rect 264166 438618 294650 438854
rect 294886 438618 325370 438854
rect 325606 438618 356090 438854
rect 356326 438618 386810 438854
rect 387046 438618 417530 438854
rect 417766 438618 448250 438854
rect 448486 438618 478970 438854
rect 479206 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 586302 438854
rect 586538 438618 586622 438854
rect 586858 438618 592650 438854
rect -8726 438586 592650 438618
rect -8726 435454 592650 435486
rect -8726 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 64250 435454
rect 64486 435218 73826 435454
rect 74062 435218 74146 435454
rect 74382 435218 94970 435454
rect 95206 435218 125690 435454
rect 125926 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 156410 435454
rect 156646 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 187130 435454
rect 187366 435218 217850 435454
rect 218086 435218 248570 435454
rect 248806 435218 279290 435454
rect 279526 435218 310010 435454
rect 310246 435218 340730 435454
rect 340966 435218 371450 435454
rect 371686 435218 402170 435454
rect 402406 435218 432890 435454
rect 433126 435218 463610 435454
rect 463846 435218 494330 435454
rect 494566 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 592650 435454
rect -8726 435134 592650 435218
rect -8726 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 64250 435134
rect 64486 434898 73826 435134
rect 74062 434898 74146 435134
rect 74382 434898 94970 435134
rect 95206 434898 125690 435134
rect 125926 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 156410 435134
rect 156646 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 187130 435134
rect 187366 434898 217850 435134
rect 218086 434898 248570 435134
rect 248806 434898 279290 435134
rect 279526 434898 310010 435134
rect 310246 434898 340730 435134
rect 340966 434898 371450 435134
rect 371686 434898 402170 435134
rect 402406 434898 432890 435134
rect 433126 434898 463610 435134
rect 463846 434898 494330 435134
rect 494566 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 592650 435134
rect -8726 434866 592650 434898
rect -8726 425494 592650 425526
rect -8726 425258 -8694 425494
rect -8458 425258 -8374 425494
rect -8138 425258 27866 425494
rect 28102 425258 28186 425494
rect 28422 425258 99866 425494
rect 100102 425258 100186 425494
rect 100422 425258 135866 425494
rect 136102 425258 136186 425494
rect 136422 425258 531866 425494
rect 532102 425258 532186 425494
rect 532422 425258 567866 425494
rect 568102 425258 568186 425494
rect 568422 425258 592062 425494
rect 592298 425258 592382 425494
rect 592618 425258 592650 425494
rect -8726 425174 592650 425258
rect -8726 424938 -8694 425174
rect -8458 424938 -8374 425174
rect -8138 424938 27866 425174
rect 28102 424938 28186 425174
rect 28422 424938 99866 425174
rect 100102 424938 100186 425174
rect 100422 424938 135866 425174
rect 136102 424938 136186 425174
rect 136422 424938 531866 425174
rect 532102 424938 532186 425174
rect 532422 424938 567866 425174
rect 568102 424938 568186 425174
rect 568422 424938 592062 425174
rect 592298 424938 592382 425174
rect 592618 424938 592650 425174
rect -8726 424906 592650 424938
rect -8726 421774 592650 421806
rect -8726 421538 -7734 421774
rect -7498 421538 -7414 421774
rect -7178 421538 24146 421774
rect 24382 421538 24466 421774
rect 24702 421538 60146 421774
rect 60382 421538 60466 421774
rect 60702 421538 96146 421774
rect 96382 421538 96466 421774
rect 96702 421538 132146 421774
rect 132382 421538 132466 421774
rect 132702 421538 168146 421774
rect 168382 421538 168466 421774
rect 168702 421538 528146 421774
rect 528382 421538 528466 421774
rect 528702 421538 564146 421774
rect 564382 421538 564466 421774
rect 564702 421538 591102 421774
rect 591338 421538 591422 421774
rect 591658 421538 592650 421774
rect -8726 421454 592650 421538
rect -8726 421218 -7734 421454
rect -7498 421218 -7414 421454
rect -7178 421218 24146 421454
rect 24382 421218 24466 421454
rect 24702 421218 60146 421454
rect 60382 421218 60466 421454
rect 60702 421218 96146 421454
rect 96382 421218 96466 421454
rect 96702 421218 132146 421454
rect 132382 421218 132466 421454
rect 132702 421218 168146 421454
rect 168382 421218 168466 421454
rect 168702 421218 528146 421454
rect 528382 421218 528466 421454
rect 528702 421218 564146 421454
rect 564382 421218 564466 421454
rect 564702 421218 591102 421454
rect 591338 421218 591422 421454
rect 591658 421218 592650 421454
rect -8726 421186 592650 421218
rect -8726 418054 592650 418086
rect -8726 417818 -6774 418054
rect -6538 417818 -6454 418054
rect -6218 417818 20426 418054
rect 20662 417818 20746 418054
rect 20982 417818 56426 418054
rect 56662 417818 56746 418054
rect 56982 417818 92426 418054
rect 92662 417818 92746 418054
rect 92982 417818 128426 418054
rect 128662 417818 128746 418054
rect 128982 417818 164426 418054
rect 164662 417818 164746 418054
rect 164982 417818 524426 418054
rect 524662 417818 524746 418054
rect 524982 417818 560426 418054
rect 560662 417818 560746 418054
rect 560982 417818 590142 418054
rect 590378 417818 590462 418054
rect 590698 417818 592650 418054
rect -8726 417734 592650 417818
rect -8726 417498 -6774 417734
rect -6538 417498 -6454 417734
rect -6218 417498 20426 417734
rect 20662 417498 20746 417734
rect 20982 417498 56426 417734
rect 56662 417498 56746 417734
rect 56982 417498 92426 417734
rect 92662 417498 92746 417734
rect 92982 417498 128426 417734
rect 128662 417498 128746 417734
rect 128982 417498 164426 417734
rect 164662 417498 164746 417734
rect 164982 417498 524426 417734
rect 524662 417498 524746 417734
rect 524982 417498 560426 417734
rect 560662 417498 560746 417734
rect 560982 417498 590142 417734
rect 590378 417498 590462 417734
rect 590698 417498 592650 417734
rect -8726 417466 592650 417498
rect -8726 414334 592650 414366
rect -8726 414098 -5814 414334
rect -5578 414098 -5494 414334
rect -5258 414098 16706 414334
rect 16942 414098 17026 414334
rect 17262 414098 52706 414334
rect 52942 414098 53026 414334
rect 53262 414098 88706 414334
rect 88942 414098 89026 414334
rect 89262 414098 124706 414334
rect 124942 414098 125026 414334
rect 125262 414098 160706 414334
rect 160942 414098 161026 414334
rect 161262 414098 196706 414334
rect 196942 414098 197026 414334
rect 197262 414098 520706 414334
rect 520942 414098 521026 414334
rect 521262 414098 556706 414334
rect 556942 414098 557026 414334
rect 557262 414098 589182 414334
rect 589418 414098 589502 414334
rect 589738 414098 592650 414334
rect -8726 414014 592650 414098
rect -8726 413778 -5814 414014
rect -5578 413778 -5494 414014
rect -5258 413778 16706 414014
rect 16942 413778 17026 414014
rect 17262 413778 52706 414014
rect 52942 413778 53026 414014
rect 53262 413778 88706 414014
rect 88942 413778 89026 414014
rect 89262 413778 124706 414014
rect 124942 413778 125026 414014
rect 125262 413778 160706 414014
rect 160942 413778 161026 414014
rect 161262 413778 196706 414014
rect 196942 413778 197026 414014
rect 197262 413778 520706 414014
rect 520942 413778 521026 414014
rect 521262 413778 556706 414014
rect 556942 413778 557026 414014
rect 557262 413778 589182 414014
rect 589418 413778 589502 414014
rect 589738 413778 592650 414014
rect -8726 413746 592650 413778
rect -8726 410614 592650 410646
rect -8726 410378 -4854 410614
rect -4618 410378 -4534 410614
rect -4298 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 84986 410614
rect 85222 410378 85306 410614
rect 85542 410378 120986 410614
rect 121222 410378 121306 410614
rect 121542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 588222 410614
rect 588458 410378 588542 410614
rect 588778 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -4854 410294
rect -4618 410058 -4534 410294
rect -4298 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 84986 410294
rect 85222 410058 85306 410294
rect 85542 410058 120986 410294
rect 121222 410058 121306 410294
rect 121542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 588222 410294
rect 588458 410058 588542 410294
rect 588778 410058 592650 410294
rect -8726 410026 592650 410058
rect -8726 406894 592650 406926
rect -8726 406658 -3894 406894
rect -3658 406658 -3574 406894
rect -3338 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 81266 406894
rect 81502 406658 81586 406894
rect 81822 406658 117266 406894
rect 117502 406658 117586 406894
rect 117822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 587262 406894
rect 587498 406658 587582 406894
rect 587818 406658 592650 406894
rect -8726 406574 592650 406658
rect -8726 406338 -3894 406574
rect -3658 406338 -3574 406574
rect -3338 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 81266 406574
rect 81502 406338 81586 406574
rect 81822 406338 117266 406574
rect 117502 406338 117586 406574
rect 117822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 587262 406574
rect 587498 406338 587582 406574
rect 587818 406338 592650 406574
rect -8726 406306 592650 406338
rect -8726 403174 592650 403206
rect -8726 402938 -2934 403174
rect -2698 402938 -2614 403174
rect -2378 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 77546 403174
rect 77782 402938 77866 403174
rect 78102 402938 79610 403174
rect 79846 402938 110330 403174
rect 110566 402938 113546 403174
rect 113782 402938 113866 403174
rect 114102 402938 141050 403174
rect 141286 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 171770 403174
rect 172006 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 202490 403174
rect 202726 402938 233210 403174
rect 233446 402938 263930 403174
rect 264166 402938 294650 403174
rect 294886 402938 325370 403174
rect 325606 402938 356090 403174
rect 356326 402938 386810 403174
rect 387046 402938 417530 403174
rect 417766 402938 448250 403174
rect 448486 402938 478970 403174
rect 479206 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 586302 403174
rect 586538 402938 586622 403174
rect 586858 402938 592650 403174
rect -8726 402854 592650 402938
rect -8726 402618 -2934 402854
rect -2698 402618 -2614 402854
rect -2378 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 77546 402854
rect 77782 402618 77866 402854
rect 78102 402618 79610 402854
rect 79846 402618 110330 402854
rect 110566 402618 113546 402854
rect 113782 402618 113866 402854
rect 114102 402618 141050 402854
rect 141286 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 171770 402854
rect 172006 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 202490 402854
rect 202726 402618 233210 402854
rect 233446 402618 263930 402854
rect 264166 402618 294650 402854
rect 294886 402618 325370 402854
rect 325606 402618 356090 402854
rect 356326 402618 386810 402854
rect 387046 402618 417530 402854
rect 417766 402618 448250 402854
rect 448486 402618 478970 402854
rect 479206 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 586302 402854
rect 586538 402618 586622 402854
rect 586858 402618 592650 402854
rect -8726 402586 592650 402618
rect -8726 399454 592650 399486
rect -8726 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 64250 399454
rect 64486 399218 73826 399454
rect 74062 399218 74146 399454
rect 74382 399218 94970 399454
rect 95206 399218 125690 399454
rect 125926 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 156410 399454
rect 156646 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 187130 399454
rect 187366 399218 217850 399454
rect 218086 399218 248570 399454
rect 248806 399218 279290 399454
rect 279526 399218 310010 399454
rect 310246 399218 340730 399454
rect 340966 399218 371450 399454
rect 371686 399218 402170 399454
rect 402406 399218 432890 399454
rect 433126 399218 463610 399454
rect 463846 399218 494330 399454
rect 494566 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 592650 399454
rect -8726 399134 592650 399218
rect -8726 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 64250 399134
rect 64486 398898 73826 399134
rect 74062 398898 74146 399134
rect 74382 398898 94970 399134
rect 95206 398898 125690 399134
rect 125926 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 156410 399134
rect 156646 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 187130 399134
rect 187366 398898 217850 399134
rect 218086 398898 248570 399134
rect 248806 398898 279290 399134
rect 279526 398898 310010 399134
rect 310246 398898 340730 399134
rect 340966 398898 371450 399134
rect 371686 398898 402170 399134
rect 402406 398898 432890 399134
rect 433126 398898 463610 399134
rect 463846 398898 494330 399134
rect 494566 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 592650 399134
rect -8726 398866 592650 398898
rect -8726 389494 592650 389526
rect -8726 389258 -8694 389494
rect -8458 389258 -8374 389494
rect -8138 389258 27866 389494
rect 28102 389258 28186 389494
rect 28422 389258 63866 389494
rect 64102 389258 64186 389494
rect 64422 389258 99866 389494
rect 100102 389258 100186 389494
rect 100422 389258 135866 389494
rect 136102 389258 136186 389494
rect 136422 389258 171866 389494
rect 172102 389258 172186 389494
rect 172422 389258 531866 389494
rect 532102 389258 532186 389494
rect 532422 389258 567866 389494
rect 568102 389258 568186 389494
rect 568422 389258 592062 389494
rect 592298 389258 592382 389494
rect 592618 389258 592650 389494
rect -8726 389174 592650 389258
rect -8726 388938 -8694 389174
rect -8458 388938 -8374 389174
rect -8138 388938 27866 389174
rect 28102 388938 28186 389174
rect 28422 388938 63866 389174
rect 64102 388938 64186 389174
rect 64422 388938 99866 389174
rect 100102 388938 100186 389174
rect 100422 388938 135866 389174
rect 136102 388938 136186 389174
rect 136422 388938 171866 389174
rect 172102 388938 172186 389174
rect 172422 388938 531866 389174
rect 532102 388938 532186 389174
rect 532422 388938 567866 389174
rect 568102 388938 568186 389174
rect 568422 388938 592062 389174
rect 592298 388938 592382 389174
rect 592618 388938 592650 389174
rect -8726 388906 592650 388938
rect -8726 385774 592650 385806
rect -8726 385538 -7734 385774
rect -7498 385538 -7414 385774
rect -7178 385538 24146 385774
rect 24382 385538 24466 385774
rect 24702 385538 60146 385774
rect 60382 385538 60466 385774
rect 60702 385538 96146 385774
rect 96382 385538 96466 385774
rect 96702 385538 132146 385774
rect 132382 385538 132466 385774
rect 132702 385538 168146 385774
rect 168382 385538 168466 385774
rect 168702 385538 204146 385774
rect 204382 385538 204466 385774
rect 204702 385538 240146 385774
rect 240382 385538 240466 385774
rect 240702 385538 276146 385774
rect 276382 385538 276466 385774
rect 276702 385538 312146 385774
rect 312382 385538 312466 385774
rect 312702 385538 348146 385774
rect 348382 385538 348466 385774
rect 348702 385538 384146 385774
rect 384382 385538 384466 385774
rect 384702 385538 420146 385774
rect 420382 385538 420466 385774
rect 420702 385538 456146 385774
rect 456382 385538 456466 385774
rect 456702 385538 492146 385774
rect 492382 385538 492466 385774
rect 492702 385538 528146 385774
rect 528382 385538 528466 385774
rect 528702 385538 564146 385774
rect 564382 385538 564466 385774
rect 564702 385538 591102 385774
rect 591338 385538 591422 385774
rect 591658 385538 592650 385774
rect -8726 385454 592650 385538
rect -8726 385218 -7734 385454
rect -7498 385218 -7414 385454
rect -7178 385218 24146 385454
rect 24382 385218 24466 385454
rect 24702 385218 60146 385454
rect 60382 385218 60466 385454
rect 60702 385218 96146 385454
rect 96382 385218 96466 385454
rect 96702 385218 132146 385454
rect 132382 385218 132466 385454
rect 132702 385218 168146 385454
rect 168382 385218 168466 385454
rect 168702 385218 204146 385454
rect 204382 385218 204466 385454
rect 204702 385218 240146 385454
rect 240382 385218 240466 385454
rect 240702 385218 276146 385454
rect 276382 385218 276466 385454
rect 276702 385218 312146 385454
rect 312382 385218 312466 385454
rect 312702 385218 348146 385454
rect 348382 385218 348466 385454
rect 348702 385218 384146 385454
rect 384382 385218 384466 385454
rect 384702 385218 420146 385454
rect 420382 385218 420466 385454
rect 420702 385218 456146 385454
rect 456382 385218 456466 385454
rect 456702 385218 492146 385454
rect 492382 385218 492466 385454
rect 492702 385218 528146 385454
rect 528382 385218 528466 385454
rect 528702 385218 564146 385454
rect 564382 385218 564466 385454
rect 564702 385218 591102 385454
rect 591338 385218 591422 385454
rect 591658 385218 592650 385454
rect -8726 385186 592650 385218
rect -8726 382054 592650 382086
rect -8726 381818 -6774 382054
rect -6538 381818 -6454 382054
rect -6218 381818 20426 382054
rect 20662 381818 20746 382054
rect 20982 381818 56426 382054
rect 56662 381818 56746 382054
rect 56982 381818 92426 382054
rect 92662 381818 92746 382054
rect 92982 381818 128426 382054
rect 128662 381818 128746 382054
rect 128982 381818 164426 382054
rect 164662 381818 164746 382054
rect 164982 381818 200426 382054
rect 200662 381818 200746 382054
rect 200982 381818 236426 382054
rect 236662 381818 236746 382054
rect 236982 381818 272426 382054
rect 272662 381818 272746 382054
rect 272982 381818 308426 382054
rect 308662 381818 308746 382054
rect 308982 381818 344426 382054
rect 344662 381818 344746 382054
rect 344982 381818 524426 382054
rect 524662 381818 524746 382054
rect 524982 381818 560426 382054
rect 560662 381818 560746 382054
rect 560982 381818 590142 382054
rect 590378 381818 590462 382054
rect 590698 381818 592650 382054
rect -8726 381734 592650 381818
rect -8726 381498 -6774 381734
rect -6538 381498 -6454 381734
rect -6218 381498 20426 381734
rect 20662 381498 20746 381734
rect 20982 381498 56426 381734
rect 56662 381498 56746 381734
rect 56982 381498 92426 381734
rect 92662 381498 92746 381734
rect 92982 381498 128426 381734
rect 128662 381498 128746 381734
rect 128982 381498 164426 381734
rect 164662 381498 164746 381734
rect 164982 381498 200426 381734
rect 200662 381498 200746 381734
rect 200982 381498 236426 381734
rect 236662 381498 236746 381734
rect 236982 381498 272426 381734
rect 272662 381498 272746 381734
rect 272982 381498 308426 381734
rect 308662 381498 308746 381734
rect 308982 381498 344426 381734
rect 344662 381498 344746 381734
rect 344982 381498 524426 381734
rect 524662 381498 524746 381734
rect 524982 381498 560426 381734
rect 560662 381498 560746 381734
rect 560982 381498 590142 381734
rect 590378 381498 590462 381734
rect 590698 381498 592650 381734
rect -8726 381466 592650 381498
rect -8726 378334 592650 378366
rect -8726 378098 -5814 378334
rect -5578 378098 -5494 378334
rect -5258 378098 16706 378334
rect 16942 378098 17026 378334
rect 17262 378098 52706 378334
rect 52942 378098 53026 378334
rect 53262 378098 88706 378334
rect 88942 378098 89026 378334
rect 89262 378098 124706 378334
rect 124942 378098 125026 378334
rect 125262 378098 160706 378334
rect 160942 378098 161026 378334
rect 161262 378098 196706 378334
rect 196942 378098 197026 378334
rect 197262 378098 232706 378334
rect 232942 378098 233026 378334
rect 233262 378098 268706 378334
rect 268942 378098 269026 378334
rect 269262 378098 304706 378334
rect 304942 378098 305026 378334
rect 305262 378098 340706 378334
rect 340942 378098 341026 378334
rect 341262 378098 520706 378334
rect 520942 378098 521026 378334
rect 521262 378098 556706 378334
rect 556942 378098 557026 378334
rect 557262 378098 589182 378334
rect 589418 378098 589502 378334
rect 589738 378098 592650 378334
rect -8726 378014 592650 378098
rect -8726 377778 -5814 378014
rect -5578 377778 -5494 378014
rect -5258 377778 16706 378014
rect 16942 377778 17026 378014
rect 17262 377778 52706 378014
rect 52942 377778 53026 378014
rect 53262 377778 88706 378014
rect 88942 377778 89026 378014
rect 89262 377778 124706 378014
rect 124942 377778 125026 378014
rect 125262 377778 160706 378014
rect 160942 377778 161026 378014
rect 161262 377778 196706 378014
rect 196942 377778 197026 378014
rect 197262 377778 232706 378014
rect 232942 377778 233026 378014
rect 233262 377778 268706 378014
rect 268942 377778 269026 378014
rect 269262 377778 304706 378014
rect 304942 377778 305026 378014
rect 305262 377778 340706 378014
rect 340942 377778 341026 378014
rect 341262 377778 520706 378014
rect 520942 377778 521026 378014
rect 521262 377778 556706 378014
rect 556942 377778 557026 378014
rect 557262 377778 589182 378014
rect 589418 377778 589502 378014
rect 589738 377778 592650 378014
rect -8726 377746 592650 377778
rect -8726 374614 592650 374646
rect -8726 374378 -4854 374614
rect -4618 374378 -4534 374614
rect -4298 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 588222 374614
rect 588458 374378 588542 374614
rect 588778 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -4854 374294
rect -4618 374058 -4534 374294
rect -4298 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 588222 374294
rect 588458 374058 588542 374294
rect 588778 374058 592650 374294
rect -8726 374026 592650 374058
rect -8726 370894 592650 370926
rect -8726 370658 -3894 370894
rect -3658 370658 -3574 370894
rect -3338 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 587262 370894
rect 587498 370658 587582 370894
rect 587818 370658 592650 370894
rect -8726 370574 592650 370658
rect -8726 370338 -3894 370574
rect -3658 370338 -3574 370574
rect -3338 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 587262 370574
rect 587498 370338 587582 370574
rect 587818 370338 592650 370574
rect -8726 370306 592650 370338
rect -8726 367174 592650 367206
rect -8726 366938 -2934 367174
rect -2698 366938 -2614 367174
rect -2378 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 586302 367174
rect 586538 366938 586622 367174
rect 586858 366938 592650 367174
rect -8726 366854 592650 366938
rect -8726 366618 -2934 366854
rect -2698 366618 -2614 366854
rect -2378 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 586302 366854
rect 586538 366618 586622 366854
rect 586858 366618 592650 366854
rect -8726 366586 592650 366618
rect -8726 363454 592650 363486
rect -8726 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 592650 363454
rect -8726 363134 592650 363218
rect -8726 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 592650 363134
rect -8726 362866 592650 362898
rect -8726 353494 592650 353526
rect -8726 353258 -8694 353494
rect -8458 353258 -8374 353494
rect -8138 353258 27866 353494
rect 28102 353258 28186 353494
rect 28422 353258 63866 353494
rect 64102 353258 64186 353494
rect 64422 353258 99866 353494
rect 100102 353258 100186 353494
rect 100422 353258 135866 353494
rect 136102 353258 136186 353494
rect 136422 353258 171866 353494
rect 172102 353258 172186 353494
rect 172422 353258 207866 353494
rect 208102 353258 208186 353494
rect 208422 353258 315866 353494
rect 316102 353258 316186 353494
rect 316422 353258 351866 353494
rect 352102 353258 352186 353494
rect 352422 353258 531866 353494
rect 532102 353258 532186 353494
rect 532422 353258 567866 353494
rect 568102 353258 568186 353494
rect 568422 353258 592062 353494
rect 592298 353258 592382 353494
rect 592618 353258 592650 353494
rect -8726 353174 592650 353258
rect -8726 352938 -8694 353174
rect -8458 352938 -8374 353174
rect -8138 352938 27866 353174
rect 28102 352938 28186 353174
rect 28422 352938 63866 353174
rect 64102 352938 64186 353174
rect 64422 352938 99866 353174
rect 100102 352938 100186 353174
rect 100422 352938 135866 353174
rect 136102 352938 136186 353174
rect 136422 352938 171866 353174
rect 172102 352938 172186 353174
rect 172422 352938 207866 353174
rect 208102 352938 208186 353174
rect 208422 352938 315866 353174
rect 316102 352938 316186 353174
rect 316422 352938 351866 353174
rect 352102 352938 352186 353174
rect 352422 352938 531866 353174
rect 532102 352938 532186 353174
rect 532422 352938 567866 353174
rect 568102 352938 568186 353174
rect 568422 352938 592062 353174
rect 592298 352938 592382 353174
rect 592618 352938 592650 353174
rect -8726 352906 592650 352938
rect -8726 349774 592650 349806
rect -8726 349538 -7734 349774
rect -7498 349538 -7414 349774
rect -7178 349538 24146 349774
rect 24382 349538 24466 349774
rect 24702 349538 60146 349774
rect 60382 349538 60466 349774
rect 60702 349538 96146 349774
rect 96382 349538 96466 349774
rect 96702 349538 132146 349774
rect 132382 349538 132466 349774
rect 132702 349538 168146 349774
rect 168382 349538 168466 349774
rect 168702 349538 204146 349774
rect 204382 349538 204466 349774
rect 204702 349538 240146 349774
rect 240382 349538 240466 349774
rect 240702 349538 276146 349774
rect 276382 349538 276466 349774
rect 276702 349538 312146 349774
rect 312382 349538 312466 349774
rect 312702 349538 348146 349774
rect 348382 349538 348466 349774
rect 348702 349538 384146 349774
rect 384382 349538 384466 349774
rect 384702 349538 420146 349774
rect 420382 349538 420466 349774
rect 420702 349538 492146 349774
rect 492382 349538 492466 349774
rect 492702 349538 528146 349774
rect 528382 349538 528466 349774
rect 528702 349538 564146 349774
rect 564382 349538 564466 349774
rect 564702 349538 591102 349774
rect 591338 349538 591422 349774
rect 591658 349538 592650 349774
rect -8726 349454 592650 349538
rect -8726 349218 -7734 349454
rect -7498 349218 -7414 349454
rect -7178 349218 24146 349454
rect 24382 349218 24466 349454
rect 24702 349218 60146 349454
rect 60382 349218 60466 349454
rect 60702 349218 96146 349454
rect 96382 349218 96466 349454
rect 96702 349218 132146 349454
rect 132382 349218 132466 349454
rect 132702 349218 168146 349454
rect 168382 349218 168466 349454
rect 168702 349218 204146 349454
rect 204382 349218 204466 349454
rect 204702 349218 240146 349454
rect 240382 349218 240466 349454
rect 240702 349218 276146 349454
rect 276382 349218 276466 349454
rect 276702 349218 312146 349454
rect 312382 349218 312466 349454
rect 312702 349218 348146 349454
rect 348382 349218 348466 349454
rect 348702 349218 384146 349454
rect 384382 349218 384466 349454
rect 384702 349218 420146 349454
rect 420382 349218 420466 349454
rect 420702 349218 492146 349454
rect 492382 349218 492466 349454
rect 492702 349218 528146 349454
rect 528382 349218 528466 349454
rect 528702 349218 564146 349454
rect 564382 349218 564466 349454
rect 564702 349218 591102 349454
rect 591338 349218 591422 349454
rect 591658 349218 592650 349454
rect -8726 349186 592650 349218
rect -8726 346054 592650 346086
rect -8726 345818 -6774 346054
rect -6538 345818 -6454 346054
rect -6218 345818 20426 346054
rect 20662 345818 20746 346054
rect 20982 345818 56426 346054
rect 56662 345818 56746 346054
rect 56982 345818 92426 346054
rect 92662 345818 92746 346054
rect 92982 345818 128426 346054
rect 128662 345818 128746 346054
rect 128982 345818 164426 346054
rect 164662 345818 164746 346054
rect 164982 345818 200426 346054
rect 200662 345818 200746 346054
rect 200982 345818 236426 346054
rect 236662 345818 236746 346054
rect 236982 345818 272426 346054
rect 272662 345818 272746 346054
rect 272982 345818 308426 346054
rect 308662 345818 308746 346054
rect 308982 345818 344426 346054
rect 344662 345818 344746 346054
rect 344982 345818 524426 346054
rect 524662 345818 524746 346054
rect 524982 345818 560426 346054
rect 560662 345818 560746 346054
rect 560982 345818 590142 346054
rect 590378 345818 590462 346054
rect 590698 345818 592650 346054
rect -8726 345734 592650 345818
rect -8726 345498 -6774 345734
rect -6538 345498 -6454 345734
rect -6218 345498 20426 345734
rect 20662 345498 20746 345734
rect 20982 345498 56426 345734
rect 56662 345498 56746 345734
rect 56982 345498 92426 345734
rect 92662 345498 92746 345734
rect 92982 345498 128426 345734
rect 128662 345498 128746 345734
rect 128982 345498 164426 345734
rect 164662 345498 164746 345734
rect 164982 345498 200426 345734
rect 200662 345498 200746 345734
rect 200982 345498 236426 345734
rect 236662 345498 236746 345734
rect 236982 345498 272426 345734
rect 272662 345498 272746 345734
rect 272982 345498 308426 345734
rect 308662 345498 308746 345734
rect 308982 345498 344426 345734
rect 344662 345498 344746 345734
rect 344982 345498 524426 345734
rect 524662 345498 524746 345734
rect 524982 345498 560426 345734
rect 560662 345498 560746 345734
rect 560982 345498 590142 345734
rect 590378 345498 590462 345734
rect 590698 345498 592650 345734
rect -8726 345466 592650 345498
rect -8726 342334 592650 342366
rect -8726 342098 -5814 342334
rect -5578 342098 -5494 342334
rect -5258 342098 16706 342334
rect 16942 342098 17026 342334
rect 17262 342098 52706 342334
rect 52942 342098 53026 342334
rect 53262 342098 88706 342334
rect 88942 342098 89026 342334
rect 89262 342098 124706 342334
rect 124942 342098 125026 342334
rect 125262 342098 160706 342334
rect 160942 342098 161026 342334
rect 161262 342098 196706 342334
rect 196942 342098 197026 342334
rect 197262 342098 232706 342334
rect 232942 342098 233026 342334
rect 233262 342098 268706 342334
rect 268942 342098 269026 342334
rect 269262 342098 304706 342334
rect 304942 342098 305026 342334
rect 305262 342098 340706 342334
rect 340942 342098 341026 342334
rect 341262 342098 520706 342334
rect 520942 342098 521026 342334
rect 521262 342098 556706 342334
rect 556942 342098 557026 342334
rect 557262 342098 589182 342334
rect 589418 342098 589502 342334
rect 589738 342098 592650 342334
rect -8726 342014 592650 342098
rect -8726 341778 -5814 342014
rect -5578 341778 -5494 342014
rect -5258 341778 16706 342014
rect 16942 341778 17026 342014
rect 17262 341778 52706 342014
rect 52942 341778 53026 342014
rect 53262 341778 88706 342014
rect 88942 341778 89026 342014
rect 89262 341778 124706 342014
rect 124942 341778 125026 342014
rect 125262 341778 160706 342014
rect 160942 341778 161026 342014
rect 161262 341778 196706 342014
rect 196942 341778 197026 342014
rect 197262 341778 232706 342014
rect 232942 341778 233026 342014
rect 233262 341778 268706 342014
rect 268942 341778 269026 342014
rect 269262 341778 304706 342014
rect 304942 341778 305026 342014
rect 305262 341778 340706 342014
rect 340942 341778 341026 342014
rect 341262 341778 520706 342014
rect 520942 341778 521026 342014
rect 521262 341778 556706 342014
rect 556942 341778 557026 342014
rect 557262 341778 589182 342014
rect 589418 341778 589502 342014
rect 589738 341778 592650 342014
rect -8726 341746 592650 341778
rect -8726 338614 592650 338646
rect -8726 338378 -4854 338614
rect -4618 338378 -4534 338614
rect -4298 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 588222 338614
rect 588458 338378 588542 338614
rect 588778 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -4854 338294
rect -4618 338058 -4534 338294
rect -4298 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 588222 338294
rect 588458 338058 588542 338294
rect 588778 338058 592650 338294
rect -8726 338026 592650 338058
rect -8726 334894 592650 334926
rect -8726 334658 -3894 334894
rect -3658 334658 -3574 334894
rect -3338 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 587262 334894
rect 587498 334658 587582 334894
rect 587818 334658 592650 334894
rect -8726 334574 592650 334658
rect -8726 334338 -3894 334574
rect -3658 334338 -3574 334574
rect -3338 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 587262 334574
rect 587498 334338 587582 334574
rect 587818 334338 592650 334574
rect -8726 334306 592650 334338
rect -8726 331174 592650 331206
rect -8726 330938 -2934 331174
rect -2698 330938 -2614 331174
rect -2378 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 259610 331174
rect 259846 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 379610 331174
rect 379846 330938 410330 331174
rect 410566 330938 441050 331174
rect 441286 330938 471770 331174
rect 472006 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 586302 331174
rect 586538 330938 586622 331174
rect 586858 330938 592650 331174
rect -8726 330854 592650 330938
rect -8726 330618 -2934 330854
rect -2698 330618 -2614 330854
rect -2378 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 259610 330854
rect 259846 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 379610 330854
rect 379846 330618 410330 330854
rect 410566 330618 441050 330854
rect 441286 330618 471770 330854
rect 472006 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 586302 330854
rect 586538 330618 586622 330854
rect 586858 330618 592650 330854
rect -8726 330586 592650 330618
rect -8726 327454 592650 327486
rect -8726 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 244250 327454
rect 244486 327218 274970 327454
rect 275206 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 364250 327454
rect 364486 327218 394970 327454
rect 395206 327218 425690 327454
rect 425926 327218 456410 327454
rect 456646 327218 487130 327454
rect 487366 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 592650 327454
rect -8726 327134 592650 327218
rect -8726 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 244250 327134
rect 244486 326898 274970 327134
rect 275206 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 364250 327134
rect 364486 326898 394970 327134
rect 395206 326898 425690 327134
rect 425926 326898 456410 327134
rect 456646 326898 487130 327134
rect 487366 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 592650 327134
rect -8726 326866 592650 326898
rect -8726 317494 592650 317526
rect -8726 317258 -8694 317494
rect -8458 317258 -8374 317494
rect -8138 317258 27866 317494
rect 28102 317258 28186 317494
rect 28422 317258 63866 317494
rect 64102 317258 64186 317494
rect 64422 317258 99866 317494
rect 100102 317258 100186 317494
rect 100422 317258 135866 317494
rect 136102 317258 136186 317494
rect 136422 317258 171866 317494
rect 172102 317258 172186 317494
rect 172422 317258 207866 317494
rect 208102 317258 208186 317494
rect 208422 317258 315866 317494
rect 316102 317258 316186 317494
rect 316422 317258 351866 317494
rect 352102 317258 352186 317494
rect 352422 317258 531866 317494
rect 532102 317258 532186 317494
rect 532422 317258 567866 317494
rect 568102 317258 568186 317494
rect 568422 317258 592062 317494
rect 592298 317258 592382 317494
rect 592618 317258 592650 317494
rect -8726 317174 592650 317258
rect -8726 316938 -8694 317174
rect -8458 316938 -8374 317174
rect -8138 316938 27866 317174
rect 28102 316938 28186 317174
rect 28422 316938 63866 317174
rect 64102 316938 64186 317174
rect 64422 316938 99866 317174
rect 100102 316938 100186 317174
rect 100422 316938 135866 317174
rect 136102 316938 136186 317174
rect 136422 316938 171866 317174
rect 172102 316938 172186 317174
rect 172422 316938 207866 317174
rect 208102 316938 208186 317174
rect 208422 316938 315866 317174
rect 316102 316938 316186 317174
rect 316422 316938 351866 317174
rect 352102 316938 352186 317174
rect 352422 316938 531866 317174
rect 532102 316938 532186 317174
rect 532422 316938 567866 317174
rect 568102 316938 568186 317174
rect 568422 316938 592062 317174
rect 592298 316938 592382 317174
rect 592618 316938 592650 317174
rect -8726 316906 592650 316938
rect -8726 313774 592650 313806
rect -8726 313538 -7734 313774
rect -7498 313538 -7414 313774
rect -7178 313538 24146 313774
rect 24382 313538 24466 313774
rect 24702 313538 60146 313774
rect 60382 313538 60466 313774
rect 60702 313538 96146 313774
rect 96382 313538 96466 313774
rect 96702 313538 132146 313774
rect 132382 313538 132466 313774
rect 132702 313538 168146 313774
rect 168382 313538 168466 313774
rect 168702 313538 204146 313774
rect 204382 313538 204466 313774
rect 204702 313538 312146 313774
rect 312382 313538 312466 313774
rect 312702 313538 348146 313774
rect 348382 313538 348466 313774
rect 348702 313538 528146 313774
rect 528382 313538 528466 313774
rect 528702 313538 564146 313774
rect 564382 313538 564466 313774
rect 564702 313538 591102 313774
rect 591338 313538 591422 313774
rect 591658 313538 592650 313774
rect -8726 313454 592650 313538
rect -8726 313218 -7734 313454
rect -7498 313218 -7414 313454
rect -7178 313218 24146 313454
rect 24382 313218 24466 313454
rect 24702 313218 60146 313454
rect 60382 313218 60466 313454
rect 60702 313218 96146 313454
rect 96382 313218 96466 313454
rect 96702 313218 132146 313454
rect 132382 313218 132466 313454
rect 132702 313218 168146 313454
rect 168382 313218 168466 313454
rect 168702 313218 204146 313454
rect 204382 313218 204466 313454
rect 204702 313218 312146 313454
rect 312382 313218 312466 313454
rect 312702 313218 348146 313454
rect 348382 313218 348466 313454
rect 348702 313218 528146 313454
rect 528382 313218 528466 313454
rect 528702 313218 564146 313454
rect 564382 313218 564466 313454
rect 564702 313218 591102 313454
rect 591338 313218 591422 313454
rect 591658 313218 592650 313454
rect -8726 313186 592650 313218
rect -8726 310054 592650 310086
rect -8726 309818 -6774 310054
rect -6538 309818 -6454 310054
rect -6218 309818 20426 310054
rect 20662 309818 20746 310054
rect 20982 309818 56426 310054
rect 56662 309818 56746 310054
rect 56982 309818 92426 310054
rect 92662 309818 92746 310054
rect 92982 309818 128426 310054
rect 128662 309818 128746 310054
rect 128982 309818 164426 310054
rect 164662 309818 164746 310054
rect 164982 309818 200426 310054
rect 200662 309818 200746 310054
rect 200982 309818 236426 310054
rect 236662 309818 236746 310054
rect 236982 309818 308426 310054
rect 308662 309818 308746 310054
rect 308982 309818 344426 310054
rect 344662 309818 344746 310054
rect 344982 309818 524426 310054
rect 524662 309818 524746 310054
rect 524982 309818 560426 310054
rect 560662 309818 560746 310054
rect 560982 309818 590142 310054
rect 590378 309818 590462 310054
rect 590698 309818 592650 310054
rect -8726 309734 592650 309818
rect -8726 309498 -6774 309734
rect -6538 309498 -6454 309734
rect -6218 309498 20426 309734
rect 20662 309498 20746 309734
rect 20982 309498 56426 309734
rect 56662 309498 56746 309734
rect 56982 309498 92426 309734
rect 92662 309498 92746 309734
rect 92982 309498 128426 309734
rect 128662 309498 128746 309734
rect 128982 309498 164426 309734
rect 164662 309498 164746 309734
rect 164982 309498 200426 309734
rect 200662 309498 200746 309734
rect 200982 309498 236426 309734
rect 236662 309498 236746 309734
rect 236982 309498 308426 309734
rect 308662 309498 308746 309734
rect 308982 309498 344426 309734
rect 344662 309498 344746 309734
rect 344982 309498 524426 309734
rect 524662 309498 524746 309734
rect 524982 309498 560426 309734
rect 560662 309498 560746 309734
rect 560982 309498 590142 309734
rect 590378 309498 590462 309734
rect 590698 309498 592650 309734
rect -8726 309466 592650 309498
rect -8726 306334 592650 306366
rect -8726 306098 -5814 306334
rect -5578 306098 -5494 306334
rect -5258 306098 16706 306334
rect 16942 306098 17026 306334
rect 17262 306098 52706 306334
rect 52942 306098 53026 306334
rect 53262 306098 88706 306334
rect 88942 306098 89026 306334
rect 89262 306098 124706 306334
rect 124942 306098 125026 306334
rect 125262 306098 160706 306334
rect 160942 306098 161026 306334
rect 161262 306098 196706 306334
rect 196942 306098 197026 306334
rect 197262 306098 232706 306334
rect 232942 306098 233026 306334
rect 233262 306098 304706 306334
rect 304942 306098 305026 306334
rect 305262 306098 340706 306334
rect 340942 306098 341026 306334
rect 341262 306098 520706 306334
rect 520942 306098 521026 306334
rect 521262 306098 556706 306334
rect 556942 306098 557026 306334
rect 557262 306098 589182 306334
rect 589418 306098 589502 306334
rect 589738 306098 592650 306334
rect -8726 306014 592650 306098
rect -8726 305778 -5814 306014
rect -5578 305778 -5494 306014
rect -5258 305778 16706 306014
rect 16942 305778 17026 306014
rect 17262 305778 52706 306014
rect 52942 305778 53026 306014
rect 53262 305778 88706 306014
rect 88942 305778 89026 306014
rect 89262 305778 124706 306014
rect 124942 305778 125026 306014
rect 125262 305778 160706 306014
rect 160942 305778 161026 306014
rect 161262 305778 196706 306014
rect 196942 305778 197026 306014
rect 197262 305778 232706 306014
rect 232942 305778 233026 306014
rect 233262 305778 304706 306014
rect 304942 305778 305026 306014
rect 305262 305778 340706 306014
rect 340942 305778 341026 306014
rect 341262 305778 520706 306014
rect 520942 305778 521026 306014
rect 521262 305778 556706 306014
rect 556942 305778 557026 306014
rect 557262 305778 589182 306014
rect 589418 305778 589502 306014
rect 589738 305778 592650 306014
rect -8726 305746 592650 305778
rect -8726 302614 592650 302646
rect -8726 302378 -4854 302614
rect -4618 302378 -4534 302614
rect -4298 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 588222 302614
rect 588458 302378 588542 302614
rect 588778 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -4854 302294
rect -4618 302058 -4534 302294
rect -4298 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 588222 302294
rect 588458 302058 588542 302294
rect 588778 302058 592650 302294
rect -8726 302026 592650 302058
rect -8726 298894 592650 298926
rect -8726 298658 -3894 298894
rect -3658 298658 -3574 298894
rect -3338 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 587262 298894
rect 587498 298658 587582 298894
rect 587818 298658 592650 298894
rect -8726 298574 592650 298658
rect -8726 298338 -3894 298574
rect -3658 298338 -3574 298574
rect -3338 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 587262 298574
rect 587498 298338 587582 298574
rect 587818 298338 592650 298574
rect -8726 298306 592650 298338
rect -8726 295174 592650 295206
rect -8726 294938 -2934 295174
rect -2698 294938 -2614 295174
rect -2378 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 69610 295174
rect 69846 294938 100330 295174
rect 100566 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 259610 295174
rect 259846 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 379610 295174
rect 379846 294938 410330 295174
rect 410566 294938 441050 295174
rect 441286 294938 471770 295174
rect 472006 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 586302 295174
rect 586538 294938 586622 295174
rect 586858 294938 592650 295174
rect -8726 294854 592650 294938
rect -8726 294618 -2934 294854
rect -2698 294618 -2614 294854
rect -2378 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 69610 294854
rect 69846 294618 100330 294854
rect 100566 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 259610 294854
rect 259846 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 379610 294854
rect 379846 294618 410330 294854
rect 410566 294618 441050 294854
rect 441286 294618 471770 294854
rect 472006 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 586302 294854
rect 586538 294618 586622 294854
rect 586858 294618 592650 294854
rect -8726 294586 592650 294618
rect -8726 291454 592650 291486
rect -8726 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 54250 291454
rect 54486 291218 84970 291454
rect 85206 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 244250 291454
rect 244486 291218 274970 291454
rect 275206 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 364250 291454
rect 364486 291218 394970 291454
rect 395206 291218 425690 291454
rect 425926 291218 456410 291454
rect 456646 291218 487130 291454
rect 487366 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 592650 291454
rect -8726 291134 592650 291218
rect -8726 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 54250 291134
rect 54486 290898 84970 291134
rect 85206 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 244250 291134
rect 244486 290898 274970 291134
rect 275206 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 364250 291134
rect 364486 290898 394970 291134
rect 395206 290898 425690 291134
rect 425926 290898 456410 291134
rect 456646 290898 487130 291134
rect 487366 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 592650 291134
rect -8726 290866 592650 290898
rect -8726 281494 592650 281526
rect -8726 281258 -8694 281494
rect -8458 281258 -8374 281494
rect -8138 281258 27866 281494
rect 28102 281258 28186 281494
rect 28422 281258 135866 281494
rect 136102 281258 136186 281494
rect 136422 281258 171866 281494
rect 172102 281258 172186 281494
rect 172422 281258 207866 281494
rect 208102 281258 208186 281494
rect 208422 281258 315866 281494
rect 316102 281258 316186 281494
rect 316422 281258 351866 281494
rect 352102 281258 352186 281494
rect 352422 281258 531866 281494
rect 532102 281258 532186 281494
rect 532422 281258 567866 281494
rect 568102 281258 568186 281494
rect 568422 281258 592062 281494
rect 592298 281258 592382 281494
rect 592618 281258 592650 281494
rect -8726 281174 592650 281258
rect -8726 280938 -8694 281174
rect -8458 280938 -8374 281174
rect -8138 280938 27866 281174
rect 28102 280938 28186 281174
rect 28422 280938 135866 281174
rect 136102 280938 136186 281174
rect 136422 280938 171866 281174
rect 172102 280938 172186 281174
rect 172422 280938 207866 281174
rect 208102 280938 208186 281174
rect 208422 280938 315866 281174
rect 316102 280938 316186 281174
rect 316422 280938 351866 281174
rect 352102 280938 352186 281174
rect 352422 280938 531866 281174
rect 532102 280938 532186 281174
rect 532422 280938 567866 281174
rect 568102 280938 568186 281174
rect 568422 280938 592062 281174
rect 592298 280938 592382 281174
rect 592618 280938 592650 281174
rect -8726 280906 592650 280938
rect -8726 277774 592650 277806
rect -8726 277538 -7734 277774
rect -7498 277538 -7414 277774
rect -7178 277538 24146 277774
rect 24382 277538 24466 277774
rect 24702 277538 132146 277774
rect 132382 277538 132466 277774
rect 132702 277538 168146 277774
rect 168382 277538 168466 277774
rect 168702 277538 204146 277774
rect 204382 277538 204466 277774
rect 204702 277538 312146 277774
rect 312382 277538 312466 277774
rect 312702 277538 348146 277774
rect 348382 277538 348466 277774
rect 348702 277538 528146 277774
rect 528382 277538 528466 277774
rect 528702 277538 564146 277774
rect 564382 277538 564466 277774
rect 564702 277538 591102 277774
rect 591338 277538 591422 277774
rect 591658 277538 592650 277774
rect -8726 277454 592650 277538
rect -8726 277218 -7734 277454
rect -7498 277218 -7414 277454
rect -7178 277218 24146 277454
rect 24382 277218 24466 277454
rect 24702 277218 132146 277454
rect 132382 277218 132466 277454
rect 132702 277218 168146 277454
rect 168382 277218 168466 277454
rect 168702 277218 204146 277454
rect 204382 277218 204466 277454
rect 204702 277218 312146 277454
rect 312382 277218 312466 277454
rect 312702 277218 348146 277454
rect 348382 277218 348466 277454
rect 348702 277218 528146 277454
rect 528382 277218 528466 277454
rect 528702 277218 564146 277454
rect 564382 277218 564466 277454
rect 564702 277218 591102 277454
rect 591338 277218 591422 277454
rect 591658 277218 592650 277454
rect -8726 277186 592650 277218
rect -8726 274054 592650 274086
rect -8726 273818 -6774 274054
rect -6538 273818 -6454 274054
rect -6218 273818 20426 274054
rect 20662 273818 20746 274054
rect 20982 273818 56426 274054
rect 56662 273818 56746 274054
rect 56982 273818 128426 274054
rect 128662 273818 128746 274054
rect 128982 273818 164426 274054
rect 164662 273818 164746 274054
rect 164982 273818 200426 274054
rect 200662 273818 200746 274054
rect 200982 273818 236426 274054
rect 236662 273818 236746 274054
rect 236982 273818 308426 274054
rect 308662 273818 308746 274054
rect 308982 273818 344426 274054
rect 344662 273818 344746 274054
rect 344982 273818 524426 274054
rect 524662 273818 524746 274054
rect 524982 273818 560426 274054
rect 560662 273818 560746 274054
rect 560982 273818 590142 274054
rect 590378 273818 590462 274054
rect 590698 273818 592650 274054
rect -8726 273734 592650 273818
rect -8726 273498 -6774 273734
rect -6538 273498 -6454 273734
rect -6218 273498 20426 273734
rect 20662 273498 20746 273734
rect 20982 273498 56426 273734
rect 56662 273498 56746 273734
rect 56982 273498 128426 273734
rect 128662 273498 128746 273734
rect 128982 273498 164426 273734
rect 164662 273498 164746 273734
rect 164982 273498 200426 273734
rect 200662 273498 200746 273734
rect 200982 273498 236426 273734
rect 236662 273498 236746 273734
rect 236982 273498 308426 273734
rect 308662 273498 308746 273734
rect 308982 273498 344426 273734
rect 344662 273498 344746 273734
rect 344982 273498 524426 273734
rect 524662 273498 524746 273734
rect 524982 273498 560426 273734
rect 560662 273498 560746 273734
rect 560982 273498 590142 273734
rect 590378 273498 590462 273734
rect 590698 273498 592650 273734
rect -8726 273466 592650 273498
rect -8726 270334 592650 270366
rect -8726 270098 -5814 270334
rect -5578 270098 -5494 270334
rect -5258 270098 16706 270334
rect 16942 270098 17026 270334
rect 17262 270098 52706 270334
rect 52942 270098 53026 270334
rect 53262 270098 124706 270334
rect 124942 270098 125026 270334
rect 125262 270098 160706 270334
rect 160942 270098 161026 270334
rect 161262 270098 196706 270334
rect 196942 270098 197026 270334
rect 197262 270098 232706 270334
rect 232942 270098 233026 270334
rect 233262 270098 304706 270334
rect 304942 270098 305026 270334
rect 305262 270098 340706 270334
rect 340942 270098 341026 270334
rect 341262 270098 520706 270334
rect 520942 270098 521026 270334
rect 521262 270098 556706 270334
rect 556942 270098 557026 270334
rect 557262 270098 589182 270334
rect 589418 270098 589502 270334
rect 589738 270098 592650 270334
rect -8726 270014 592650 270098
rect -8726 269778 -5814 270014
rect -5578 269778 -5494 270014
rect -5258 269778 16706 270014
rect 16942 269778 17026 270014
rect 17262 269778 52706 270014
rect 52942 269778 53026 270014
rect 53262 269778 124706 270014
rect 124942 269778 125026 270014
rect 125262 269778 160706 270014
rect 160942 269778 161026 270014
rect 161262 269778 196706 270014
rect 196942 269778 197026 270014
rect 197262 269778 232706 270014
rect 232942 269778 233026 270014
rect 233262 269778 304706 270014
rect 304942 269778 305026 270014
rect 305262 269778 340706 270014
rect 340942 269778 341026 270014
rect 341262 269778 520706 270014
rect 520942 269778 521026 270014
rect 521262 269778 556706 270014
rect 556942 269778 557026 270014
rect 557262 269778 589182 270014
rect 589418 269778 589502 270014
rect 589738 269778 592650 270014
rect -8726 269746 592650 269778
rect -8726 266614 592650 266646
rect -8726 266378 -4854 266614
rect -4618 266378 -4534 266614
rect -4298 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 588222 266614
rect 588458 266378 588542 266614
rect 588778 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -4854 266294
rect -4618 266058 -4534 266294
rect -4298 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 588222 266294
rect 588458 266058 588542 266294
rect 588778 266058 592650 266294
rect -8726 266026 592650 266058
rect -8726 262894 592650 262926
rect -8726 262658 -3894 262894
rect -3658 262658 -3574 262894
rect -3338 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 587262 262894
rect 587498 262658 587582 262894
rect 587818 262658 592650 262894
rect -8726 262574 592650 262658
rect -8726 262338 -3894 262574
rect -3658 262338 -3574 262574
rect -3338 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 587262 262574
rect 587498 262338 587582 262574
rect 587818 262338 592650 262574
rect -8726 262306 592650 262338
rect -8726 259174 592650 259206
rect -8726 258938 -2934 259174
rect -2698 258938 -2614 259174
rect -2378 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 69610 259174
rect 69846 258938 100330 259174
rect 100566 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 259610 259174
rect 259846 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 379610 259174
rect 379846 258938 410330 259174
rect 410566 258938 441050 259174
rect 441286 258938 471770 259174
rect 472006 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 586302 259174
rect 586538 258938 586622 259174
rect 586858 258938 592650 259174
rect -8726 258854 592650 258938
rect -8726 258618 -2934 258854
rect -2698 258618 -2614 258854
rect -2378 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 69610 258854
rect 69846 258618 100330 258854
rect 100566 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 259610 258854
rect 259846 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 379610 258854
rect 379846 258618 410330 258854
rect 410566 258618 441050 258854
rect 441286 258618 471770 258854
rect 472006 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 586302 258854
rect 586538 258618 586622 258854
rect 586858 258618 592650 258854
rect -8726 258586 592650 258618
rect -8726 255454 592650 255486
rect -8726 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 54250 255454
rect 54486 255218 84970 255454
rect 85206 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 244250 255454
rect 244486 255218 274970 255454
rect 275206 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 364250 255454
rect 364486 255218 394970 255454
rect 395206 255218 425690 255454
rect 425926 255218 456410 255454
rect 456646 255218 487130 255454
rect 487366 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 592650 255454
rect -8726 255134 592650 255218
rect -8726 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 54250 255134
rect 54486 254898 84970 255134
rect 85206 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 244250 255134
rect 244486 254898 274970 255134
rect 275206 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 364250 255134
rect 364486 254898 394970 255134
rect 395206 254898 425690 255134
rect 425926 254898 456410 255134
rect 456646 254898 487130 255134
rect 487366 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 592650 255134
rect -8726 254866 592650 254898
rect -8726 245494 592650 245526
rect -8726 245258 -8694 245494
rect -8458 245258 -8374 245494
rect -8138 245258 27866 245494
rect 28102 245258 28186 245494
rect 28422 245258 135866 245494
rect 136102 245258 136186 245494
rect 136422 245258 171866 245494
rect 172102 245258 172186 245494
rect 172422 245258 207866 245494
rect 208102 245258 208186 245494
rect 208422 245258 315866 245494
rect 316102 245258 316186 245494
rect 316422 245258 351866 245494
rect 352102 245258 352186 245494
rect 352422 245258 531866 245494
rect 532102 245258 532186 245494
rect 532422 245258 567866 245494
rect 568102 245258 568186 245494
rect 568422 245258 592062 245494
rect 592298 245258 592382 245494
rect 592618 245258 592650 245494
rect -8726 245174 592650 245258
rect -8726 244938 -8694 245174
rect -8458 244938 -8374 245174
rect -8138 244938 27866 245174
rect 28102 244938 28186 245174
rect 28422 244938 135866 245174
rect 136102 244938 136186 245174
rect 136422 244938 171866 245174
rect 172102 244938 172186 245174
rect 172422 244938 207866 245174
rect 208102 244938 208186 245174
rect 208422 244938 315866 245174
rect 316102 244938 316186 245174
rect 316422 244938 351866 245174
rect 352102 244938 352186 245174
rect 352422 244938 531866 245174
rect 532102 244938 532186 245174
rect 532422 244938 567866 245174
rect 568102 244938 568186 245174
rect 568422 244938 592062 245174
rect 592298 244938 592382 245174
rect 592618 244938 592650 245174
rect -8726 244906 592650 244938
rect -8726 241774 592650 241806
rect -8726 241538 -7734 241774
rect -7498 241538 -7414 241774
rect -7178 241538 24146 241774
rect 24382 241538 24466 241774
rect 24702 241538 132146 241774
rect 132382 241538 132466 241774
rect 132702 241538 168146 241774
rect 168382 241538 168466 241774
rect 168702 241538 204146 241774
rect 204382 241538 204466 241774
rect 204702 241538 312146 241774
rect 312382 241538 312466 241774
rect 312702 241538 348146 241774
rect 348382 241538 348466 241774
rect 348702 241538 528146 241774
rect 528382 241538 528466 241774
rect 528702 241538 564146 241774
rect 564382 241538 564466 241774
rect 564702 241538 591102 241774
rect 591338 241538 591422 241774
rect 591658 241538 592650 241774
rect -8726 241454 592650 241538
rect -8726 241218 -7734 241454
rect -7498 241218 -7414 241454
rect -7178 241218 24146 241454
rect 24382 241218 24466 241454
rect 24702 241218 132146 241454
rect 132382 241218 132466 241454
rect 132702 241218 168146 241454
rect 168382 241218 168466 241454
rect 168702 241218 204146 241454
rect 204382 241218 204466 241454
rect 204702 241218 312146 241454
rect 312382 241218 312466 241454
rect 312702 241218 348146 241454
rect 348382 241218 348466 241454
rect 348702 241218 528146 241454
rect 528382 241218 528466 241454
rect 528702 241218 564146 241454
rect 564382 241218 564466 241454
rect 564702 241218 591102 241454
rect 591338 241218 591422 241454
rect 591658 241218 592650 241454
rect -8726 241186 592650 241218
rect -8726 238054 592650 238086
rect -8726 237818 -6774 238054
rect -6538 237818 -6454 238054
rect -6218 237818 20426 238054
rect 20662 237818 20746 238054
rect 20982 237818 56426 238054
rect 56662 237818 56746 238054
rect 56982 237818 92426 238054
rect 92662 237818 92746 238054
rect 92982 237818 128426 238054
rect 128662 237818 128746 238054
rect 128982 237818 164426 238054
rect 164662 237818 164746 238054
rect 164982 237818 200426 238054
rect 200662 237818 200746 238054
rect 200982 237818 236426 238054
rect 236662 237818 236746 238054
rect 236982 237818 308426 238054
rect 308662 237818 308746 238054
rect 308982 237818 344426 238054
rect 344662 237818 344746 238054
rect 344982 237818 524426 238054
rect 524662 237818 524746 238054
rect 524982 237818 560426 238054
rect 560662 237818 560746 238054
rect 560982 237818 590142 238054
rect 590378 237818 590462 238054
rect 590698 237818 592650 238054
rect -8726 237734 592650 237818
rect -8726 237498 -6774 237734
rect -6538 237498 -6454 237734
rect -6218 237498 20426 237734
rect 20662 237498 20746 237734
rect 20982 237498 56426 237734
rect 56662 237498 56746 237734
rect 56982 237498 92426 237734
rect 92662 237498 92746 237734
rect 92982 237498 128426 237734
rect 128662 237498 128746 237734
rect 128982 237498 164426 237734
rect 164662 237498 164746 237734
rect 164982 237498 200426 237734
rect 200662 237498 200746 237734
rect 200982 237498 236426 237734
rect 236662 237498 236746 237734
rect 236982 237498 308426 237734
rect 308662 237498 308746 237734
rect 308982 237498 344426 237734
rect 344662 237498 344746 237734
rect 344982 237498 524426 237734
rect 524662 237498 524746 237734
rect 524982 237498 560426 237734
rect 560662 237498 560746 237734
rect 560982 237498 590142 237734
rect 590378 237498 590462 237734
rect 590698 237498 592650 237734
rect -8726 237466 592650 237498
rect -8726 234334 592650 234366
rect -8726 234098 -5814 234334
rect -5578 234098 -5494 234334
rect -5258 234098 16706 234334
rect 16942 234098 17026 234334
rect 17262 234098 52706 234334
rect 52942 234098 53026 234334
rect 53262 234098 88706 234334
rect 88942 234098 89026 234334
rect 89262 234098 124706 234334
rect 124942 234098 125026 234334
rect 125262 234098 160706 234334
rect 160942 234098 161026 234334
rect 161262 234098 196706 234334
rect 196942 234098 197026 234334
rect 197262 234098 232706 234334
rect 232942 234098 233026 234334
rect 233262 234098 304706 234334
rect 304942 234098 305026 234334
rect 305262 234098 340706 234334
rect 340942 234098 341026 234334
rect 341262 234098 520706 234334
rect 520942 234098 521026 234334
rect 521262 234098 556706 234334
rect 556942 234098 557026 234334
rect 557262 234098 589182 234334
rect 589418 234098 589502 234334
rect 589738 234098 592650 234334
rect -8726 234014 592650 234098
rect -8726 233778 -5814 234014
rect -5578 233778 -5494 234014
rect -5258 233778 16706 234014
rect 16942 233778 17026 234014
rect 17262 233778 52706 234014
rect 52942 233778 53026 234014
rect 53262 233778 88706 234014
rect 88942 233778 89026 234014
rect 89262 233778 124706 234014
rect 124942 233778 125026 234014
rect 125262 233778 160706 234014
rect 160942 233778 161026 234014
rect 161262 233778 196706 234014
rect 196942 233778 197026 234014
rect 197262 233778 232706 234014
rect 232942 233778 233026 234014
rect 233262 233778 304706 234014
rect 304942 233778 305026 234014
rect 305262 233778 340706 234014
rect 340942 233778 341026 234014
rect 341262 233778 520706 234014
rect 520942 233778 521026 234014
rect 521262 233778 556706 234014
rect 556942 233778 557026 234014
rect 557262 233778 589182 234014
rect 589418 233778 589502 234014
rect 589738 233778 592650 234014
rect -8726 233746 592650 233778
rect -8726 230614 592650 230646
rect -8726 230378 -4854 230614
rect -4618 230378 -4534 230614
rect -4298 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 588222 230614
rect 588458 230378 588542 230614
rect 588778 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -4854 230294
rect -4618 230058 -4534 230294
rect -4298 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 588222 230294
rect 588458 230058 588542 230294
rect 588778 230058 592650 230294
rect -8726 230026 592650 230058
rect -8726 226894 592650 226926
rect -8726 226658 -3894 226894
rect -3658 226658 -3574 226894
rect -3338 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 587262 226894
rect 587498 226658 587582 226894
rect 587818 226658 592650 226894
rect -8726 226574 592650 226658
rect -8726 226338 -3894 226574
rect -3658 226338 -3574 226574
rect -3338 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 587262 226574
rect 587498 226338 587582 226574
rect 587818 226338 592650 226574
rect -8726 226306 592650 226338
rect -8726 223174 592650 223206
rect -8726 222938 -2934 223174
rect -2698 222938 -2614 223174
rect -2378 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 259610 223174
rect 259846 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 379610 223174
rect 379846 222938 410330 223174
rect 410566 222938 441050 223174
rect 441286 222938 471770 223174
rect 472006 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 586302 223174
rect 586538 222938 586622 223174
rect 586858 222938 592650 223174
rect -8726 222854 592650 222938
rect -8726 222618 -2934 222854
rect -2698 222618 -2614 222854
rect -2378 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 259610 222854
rect 259846 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 379610 222854
rect 379846 222618 410330 222854
rect 410566 222618 441050 222854
rect 441286 222618 471770 222854
rect 472006 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 586302 222854
rect 586538 222618 586622 222854
rect 586858 222618 592650 222854
rect -8726 222586 592650 222618
rect -8726 219454 592650 219486
rect -8726 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 244250 219454
rect 244486 219218 274970 219454
rect 275206 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 364250 219454
rect 364486 219218 394970 219454
rect 395206 219218 425690 219454
rect 425926 219218 456410 219454
rect 456646 219218 487130 219454
rect 487366 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 592650 219454
rect -8726 219134 592650 219218
rect -8726 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 244250 219134
rect 244486 218898 274970 219134
rect 275206 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 364250 219134
rect 364486 218898 394970 219134
rect 395206 218898 425690 219134
rect 425926 218898 456410 219134
rect 456646 218898 487130 219134
rect 487366 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 592650 219134
rect -8726 218866 592650 218898
rect -8726 209494 592650 209526
rect -8726 209258 -8694 209494
rect -8458 209258 -8374 209494
rect -8138 209258 27866 209494
rect 28102 209258 28186 209494
rect 28422 209258 135866 209494
rect 136102 209258 136186 209494
rect 136422 209258 171866 209494
rect 172102 209258 172186 209494
rect 172422 209258 207866 209494
rect 208102 209258 208186 209494
rect 208422 209258 315866 209494
rect 316102 209258 316186 209494
rect 316422 209258 351866 209494
rect 352102 209258 352186 209494
rect 352422 209258 531866 209494
rect 532102 209258 532186 209494
rect 532422 209258 567866 209494
rect 568102 209258 568186 209494
rect 568422 209258 592062 209494
rect 592298 209258 592382 209494
rect 592618 209258 592650 209494
rect -8726 209174 592650 209258
rect -8726 208938 -8694 209174
rect -8458 208938 -8374 209174
rect -8138 208938 27866 209174
rect 28102 208938 28186 209174
rect 28422 208938 135866 209174
rect 136102 208938 136186 209174
rect 136422 208938 171866 209174
rect 172102 208938 172186 209174
rect 172422 208938 207866 209174
rect 208102 208938 208186 209174
rect 208422 208938 315866 209174
rect 316102 208938 316186 209174
rect 316422 208938 351866 209174
rect 352102 208938 352186 209174
rect 352422 208938 531866 209174
rect 532102 208938 532186 209174
rect 532422 208938 567866 209174
rect 568102 208938 568186 209174
rect 568422 208938 592062 209174
rect 592298 208938 592382 209174
rect 592618 208938 592650 209174
rect -8726 208906 592650 208938
rect -8726 205774 592650 205806
rect -8726 205538 -7734 205774
rect -7498 205538 -7414 205774
rect -7178 205538 24146 205774
rect 24382 205538 24466 205774
rect 24702 205538 132146 205774
rect 132382 205538 132466 205774
rect 132702 205538 168146 205774
rect 168382 205538 168466 205774
rect 168702 205538 204146 205774
rect 204382 205538 204466 205774
rect 204702 205538 312146 205774
rect 312382 205538 312466 205774
rect 312702 205538 348146 205774
rect 348382 205538 348466 205774
rect 348702 205538 528146 205774
rect 528382 205538 528466 205774
rect 528702 205538 564146 205774
rect 564382 205538 564466 205774
rect 564702 205538 591102 205774
rect 591338 205538 591422 205774
rect 591658 205538 592650 205774
rect -8726 205454 592650 205538
rect -8726 205218 -7734 205454
rect -7498 205218 -7414 205454
rect -7178 205218 24146 205454
rect 24382 205218 24466 205454
rect 24702 205218 132146 205454
rect 132382 205218 132466 205454
rect 132702 205218 168146 205454
rect 168382 205218 168466 205454
rect 168702 205218 204146 205454
rect 204382 205218 204466 205454
rect 204702 205218 312146 205454
rect 312382 205218 312466 205454
rect 312702 205218 348146 205454
rect 348382 205218 348466 205454
rect 348702 205218 528146 205454
rect 528382 205218 528466 205454
rect 528702 205218 564146 205454
rect 564382 205218 564466 205454
rect 564702 205218 591102 205454
rect 591338 205218 591422 205454
rect 591658 205218 592650 205454
rect -8726 205186 592650 205218
rect -8726 202054 592650 202086
rect -8726 201818 -6774 202054
rect -6538 201818 -6454 202054
rect -6218 201818 20426 202054
rect 20662 201818 20746 202054
rect 20982 201818 56426 202054
rect 56662 201818 56746 202054
rect 56982 201818 92426 202054
rect 92662 201818 92746 202054
rect 92982 201818 128426 202054
rect 128662 201818 128746 202054
rect 128982 201818 164426 202054
rect 164662 201818 164746 202054
rect 164982 201818 200426 202054
rect 200662 201818 200746 202054
rect 200982 201818 236426 202054
rect 236662 201818 236746 202054
rect 236982 201818 308426 202054
rect 308662 201818 308746 202054
rect 308982 201818 344426 202054
rect 344662 201818 344746 202054
rect 344982 201818 524426 202054
rect 524662 201818 524746 202054
rect 524982 201818 560426 202054
rect 560662 201818 560746 202054
rect 560982 201818 590142 202054
rect 590378 201818 590462 202054
rect 590698 201818 592650 202054
rect -8726 201734 592650 201818
rect -8726 201498 -6774 201734
rect -6538 201498 -6454 201734
rect -6218 201498 20426 201734
rect 20662 201498 20746 201734
rect 20982 201498 56426 201734
rect 56662 201498 56746 201734
rect 56982 201498 92426 201734
rect 92662 201498 92746 201734
rect 92982 201498 128426 201734
rect 128662 201498 128746 201734
rect 128982 201498 164426 201734
rect 164662 201498 164746 201734
rect 164982 201498 200426 201734
rect 200662 201498 200746 201734
rect 200982 201498 236426 201734
rect 236662 201498 236746 201734
rect 236982 201498 308426 201734
rect 308662 201498 308746 201734
rect 308982 201498 344426 201734
rect 344662 201498 344746 201734
rect 344982 201498 524426 201734
rect 524662 201498 524746 201734
rect 524982 201498 560426 201734
rect 560662 201498 560746 201734
rect 560982 201498 590142 201734
rect 590378 201498 590462 201734
rect 590698 201498 592650 201734
rect -8726 201466 592650 201498
rect -8726 198334 592650 198366
rect -8726 198098 -5814 198334
rect -5578 198098 -5494 198334
rect -5258 198098 16706 198334
rect 16942 198098 17026 198334
rect 17262 198098 52706 198334
rect 52942 198098 53026 198334
rect 53262 198098 88706 198334
rect 88942 198098 89026 198334
rect 89262 198098 124706 198334
rect 124942 198098 125026 198334
rect 125262 198098 160706 198334
rect 160942 198098 161026 198334
rect 161262 198098 196706 198334
rect 196942 198098 197026 198334
rect 197262 198098 232706 198334
rect 232942 198098 233026 198334
rect 233262 198098 304706 198334
rect 304942 198098 305026 198334
rect 305262 198098 340706 198334
rect 340942 198098 341026 198334
rect 341262 198098 520706 198334
rect 520942 198098 521026 198334
rect 521262 198098 556706 198334
rect 556942 198098 557026 198334
rect 557262 198098 589182 198334
rect 589418 198098 589502 198334
rect 589738 198098 592650 198334
rect -8726 198014 592650 198098
rect -8726 197778 -5814 198014
rect -5578 197778 -5494 198014
rect -5258 197778 16706 198014
rect 16942 197778 17026 198014
rect 17262 197778 52706 198014
rect 52942 197778 53026 198014
rect 53262 197778 88706 198014
rect 88942 197778 89026 198014
rect 89262 197778 124706 198014
rect 124942 197778 125026 198014
rect 125262 197778 160706 198014
rect 160942 197778 161026 198014
rect 161262 197778 196706 198014
rect 196942 197778 197026 198014
rect 197262 197778 232706 198014
rect 232942 197778 233026 198014
rect 233262 197778 304706 198014
rect 304942 197778 305026 198014
rect 305262 197778 340706 198014
rect 340942 197778 341026 198014
rect 341262 197778 520706 198014
rect 520942 197778 521026 198014
rect 521262 197778 556706 198014
rect 556942 197778 557026 198014
rect 557262 197778 589182 198014
rect 589418 197778 589502 198014
rect 589738 197778 592650 198014
rect -8726 197746 592650 197778
rect -8726 194614 592650 194646
rect -8726 194378 -4854 194614
rect -4618 194378 -4534 194614
rect -4298 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 588222 194614
rect 588458 194378 588542 194614
rect 588778 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -4854 194294
rect -4618 194058 -4534 194294
rect -4298 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 588222 194294
rect 588458 194058 588542 194294
rect 588778 194058 592650 194294
rect -8726 194026 592650 194058
rect -8726 190894 592650 190926
rect -8726 190658 -3894 190894
rect -3658 190658 -3574 190894
rect -3338 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 587262 190894
rect 587498 190658 587582 190894
rect 587818 190658 592650 190894
rect -8726 190574 592650 190658
rect -8726 190338 -3894 190574
rect -3658 190338 -3574 190574
rect -3338 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 587262 190574
rect 587498 190338 587582 190574
rect 587818 190338 592650 190574
rect -8726 190306 592650 190338
rect -8726 187174 592650 187206
rect -8726 186938 -2934 187174
rect -2698 186938 -2614 187174
rect -2378 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 259610 187174
rect 259846 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 379610 187174
rect 379846 186938 410330 187174
rect 410566 186938 441050 187174
rect 441286 186938 471770 187174
rect 472006 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 586302 187174
rect 586538 186938 586622 187174
rect 586858 186938 592650 187174
rect -8726 186854 592650 186938
rect -8726 186618 -2934 186854
rect -2698 186618 -2614 186854
rect -2378 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 259610 186854
rect 259846 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 379610 186854
rect 379846 186618 410330 186854
rect 410566 186618 441050 186854
rect 441286 186618 471770 186854
rect 472006 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 586302 186854
rect 586538 186618 586622 186854
rect 586858 186618 592650 186854
rect -8726 186586 592650 186618
rect -8726 183454 592650 183486
rect -8726 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 244250 183454
rect 244486 183218 274970 183454
rect 275206 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 364250 183454
rect 364486 183218 394970 183454
rect 395206 183218 425690 183454
rect 425926 183218 456410 183454
rect 456646 183218 487130 183454
rect 487366 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 592650 183454
rect -8726 183134 592650 183218
rect -8726 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 244250 183134
rect 244486 182898 274970 183134
rect 275206 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 364250 183134
rect 364486 182898 394970 183134
rect 395206 182898 425690 183134
rect 425926 182898 456410 183134
rect 456646 182898 487130 183134
rect 487366 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 592650 183134
rect -8726 182866 592650 182898
rect -8726 173494 592650 173526
rect -8726 173258 -8694 173494
rect -8458 173258 -8374 173494
rect -8138 173258 27866 173494
rect 28102 173258 28186 173494
rect 28422 173258 135866 173494
rect 136102 173258 136186 173494
rect 136422 173258 171866 173494
rect 172102 173258 172186 173494
rect 172422 173258 207866 173494
rect 208102 173258 208186 173494
rect 208422 173258 315866 173494
rect 316102 173258 316186 173494
rect 316422 173258 351866 173494
rect 352102 173258 352186 173494
rect 352422 173258 423866 173494
rect 424102 173258 424186 173494
rect 424422 173258 459866 173494
rect 460102 173258 460186 173494
rect 460422 173258 495866 173494
rect 496102 173258 496186 173494
rect 496422 173258 531866 173494
rect 532102 173258 532186 173494
rect 532422 173258 567866 173494
rect 568102 173258 568186 173494
rect 568422 173258 592062 173494
rect 592298 173258 592382 173494
rect 592618 173258 592650 173494
rect -8726 173174 592650 173258
rect -8726 172938 -8694 173174
rect -8458 172938 -8374 173174
rect -8138 172938 27866 173174
rect 28102 172938 28186 173174
rect 28422 172938 135866 173174
rect 136102 172938 136186 173174
rect 136422 172938 171866 173174
rect 172102 172938 172186 173174
rect 172422 172938 207866 173174
rect 208102 172938 208186 173174
rect 208422 172938 315866 173174
rect 316102 172938 316186 173174
rect 316422 172938 351866 173174
rect 352102 172938 352186 173174
rect 352422 172938 423866 173174
rect 424102 172938 424186 173174
rect 424422 172938 459866 173174
rect 460102 172938 460186 173174
rect 460422 172938 495866 173174
rect 496102 172938 496186 173174
rect 496422 172938 531866 173174
rect 532102 172938 532186 173174
rect 532422 172938 567866 173174
rect 568102 172938 568186 173174
rect 568422 172938 592062 173174
rect 592298 172938 592382 173174
rect 592618 172938 592650 173174
rect -8726 172906 592650 172938
rect -8726 169774 592650 169806
rect -8726 169538 -7734 169774
rect -7498 169538 -7414 169774
rect -7178 169538 24146 169774
rect 24382 169538 24466 169774
rect 24702 169538 132146 169774
rect 132382 169538 132466 169774
rect 132702 169538 168146 169774
rect 168382 169538 168466 169774
rect 168702 169538 204146 169774
rect 204382 169538 204466 169774
rect 204702 169538 312146 169774
rect 312382 169538 312466 169774
rect 312702 169538 348146 169774
rect 348382 169538 348466 169774
rect 348702 169538 420146 169774
rect 420382 169538 420466 169774
rect 420702 169538 456146 169774
rect 456382 169538 456466 169774
rect 456702 169538 492146 169774
rect 492382 169538 492466 169774
rect 492702 169538 528146 169774
rect 528382 169538 528466 169774
rect 528702 169538 564146 169774
rect 564382 169538 564466 169774
rect 564702 169538 591102 169774
rect 591338 169538 591422 169774
rect 591658 169538 592650 169774
rect -8726 169454 592650 169538
rect -8726 169218 -7734 169454
rect -7498 169218 -7414 169454
rect -7178 169218 24146 169454
rect 24382 169218 24466 169454
rect 24702 169218 132146 169454
rect 132382 169218 132466 169454
rect 132702 169218 168146 169454
rect 168382 169218 168466 169454
rect 168702 169218 204146 169454
rect 204382 169218 204466 169454
rect 204702 169218 312146 169454
rect 312382 169218 312466 169454
rect 312702 169218 348146 169454
rect 348382 169218 348466 169454
rect 348702 169218 420146 169454
rect 420382 169218 420466 169454
rect 420702 169218 456146 169454
rect 456382 169218 456466 169454
rect 456702 169218 492146 169454
rect 492382 169218 492466 169454
rect 492702 169218 528146 169454
rect 528382 169218 528466 169454
rect 528702 169218 564146 169454
rect 564382 169218 564466 169454
rect 564702 169218 591102 169454
rect 591338 169218 591422 169454
rect 591658 169218 592650 169454
rect -8726 169186 592650 169218
rect -8726 166054 592650 166086
rect -8726 165818 -6774 166054
rect -6538 165818 -6454 166054
rect -6218 165818 20426 166054
rect 20662 165818 20746 166054
rect 20982 165818 56426 166054
rect 56662 165818 56746 166054
rect 56982 165818 128426 166054
rect 128662 165818 128746 166054
rect 128982 165818 164426 166054
rect 164662 165818 164746 166054
rect 164982 165818 200426 166054
rect 200662 165818 200746 166054
rect 200982 165818 236426 166054
rect 236662 165818 236746 166054
rect 236982 165818 308426 166054
rect 308662 165818 308746 166054
rect 308982 165818 344426 166054
rect 344662 165818 344746 166054
rect 344982 165818 416426 166054
rect 416662 165818 416746 166054
rect 416982 165818 452426 166054
rect 452662 165818 452746 166054
rect 452982 165818 488426 166054
rect 488662 165818 488746 166054
rect 488982 165818 524426 166054
rect 524662 165818 524746 166054
rect 524982 165818 560426 166054
rect 560662 165818 560746 166054
rect 560982 165818 590142 166054
rect 590378 165818 590462 166054
rect 590698 165818 592650 166054
rect -8726 165734 592650 165818
rect -8726 165498 -6774 165734
rect -6538 165498 -6454 165734
rect -6218 165498 20426 165734
rect 20662 165498 20746 165734
rect 20982 165498 56426 165734
rect 56662 165498 56746 165734
rect 56982 165498 128426 165734
rect 128662 165498 128746 165734
rect 128982 165498 164426 165734
rect 164662 165498 164746 165734
rect 164982 165498 200426 165734
rect 200662 165498 200746 165734
rect 200982 165498 236426 165734
rect 236662 165498 236746 165734
rect 236982 165498 308426 165734
rect 308662 165498 308746 165734
rect 308982 165498 344426 165734
rect 344662 165498 344746 165734
rect 344982 165498 416426 165734
rect 416662 165498 416746 165734
rect 416982 165498 452426 165734
rect 452662 165498 452746 165734
rect 452982 165498 488426 165734
rect 488662 165498 488746 165734
rect 488982 165498 524426 165734
rect 524662 165498 524746 165734
rect 524982 165498 560426 165734
rect 560662 165498 560746 165734
rect 560982 165498 590142 165734
rect 590378 165498 590462 165734
rect 590698 165498 592650 165734
rect -8726 165466 592650 165498
rect -8726 162334 592650 162366
rect -8726 162098 -5814 162334
rect -5578 162098 -5494 162334
rect -5258 162098 16706 162334
rect 16942 162098 17026 162334
rect 17262 162098 52706 162334
rect 52942 162098 53026 162334
rect 53262 162098 124706 162334
rect 124942 162098 125026 162334
rect 125262 162098 160706 162334
rect 160942 162098 161026 162334
rect 161262 162098 196706 162334
rect 196942 162098 197026 162334
rect 197262 162098 232706 162334
rect 232942 162098 233026 162334
rect 233262 162098 304706 162334
rect 304942 162098 305026 162334
rect 305262 162098 340706 162334
rect 340942 162098 341026 162334
rect 341262 162098 412706 162334
rect 412942 162098 413026 162334
rect 413262 162098 448706 162334
rect 448942 162098 449026 162334
rect 449262 162098 484706 162334
rect 484942 162098 485026 162334
rect 485262 162098 520706 162334
rect 520942 162098 521026 162334
rect 521262 162098 556706 162334
rect 556942 162098 557026 162334
rect 557262 162098 589182 162334
rect 589418 162098 589502 162334
rect 589738 162098 592650 162334
rect -8726 162014 592650 162098
rect -8726 161778 -5814 162014
rect -5578 161778 -5494 162014
rect -5258 161778 16706 162014
rect 16942 161778 17026 162014
rect 17262 161778 52706 162014
rect 52942 161778 53026 162014
rect 53262 161778 124706 162014
rect 124942 161778 125026 162014
rect 125262 161778 160706 162014
rect 160942 161778 161026 162014
rect 161262 161778 196706 162014
rect 196942 161778 197026 162014
rect 197262 161778 232706 162014
rect 232942 161778 233026 162014
rect 233262 161778 304706 162014
rect 304942 161778 305026 162014
rect 305262 161778 340706 162014
rect 340942 161778 341026 162014
rect 341262 161778 412706 162014
rect 412942 161778 413026 162014
rect 413262 161778 448706 162014
rect 448942 161778 449026 162014
rect 449262 161778 484706 162014
rect 484942 161778 485026 162014
rect 485262 161778 520706 162014
rect 520942 161778 521026 162014
rect 521262 161778 556706 162014
rect 556942 161778 557026 162014
rect 557262 161778 589182 162014
rect 589418 161778 589502 162014
rect 589738 161778 592650 162014
rect -8726 161746 592650 161778
rect -8726 158614 592650 158646
rect -8726 158378 -4854 158614
rect -4618 158378 -4534 158614
rect -4298 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 588222 158614
rect 588458 158378 588542 158614
rect 588778 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -4854 158294
rect -4618 158058 -4534 158294
rect -4298 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 588222 158294
rect 588458 158058 588542 158294
rect 588778 158058 592650 158294
rect -8726 158026 592650 158058
rect -8726 154894 592650 154926
rect -8726 154658 -3894 154894
rect -3658 154658 -3574 154894
rect -3338 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 587262 154894
rect 587498 154658 587582 154894
rect 587818 154658 592650 154894
rect -8726 154574 592650 154658
rect -8726 154338 -3894 154574
rect -3658 154338 -3574 154574
rect -3338 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 587262 154574
rect 587498 154338 587582 154574
rect 587818 154338 592650 154574
rect -8726 154306 592650 154338
rect -8726 151174 592650 151206
rect -8726 150938 -2934 151174
rect -2698 150938 -2614 151174
rect -2378 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 79610 151174
rect 79846 150938 110330 151174
rect 110566 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 259610 151174
rect 259846 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 586302 151174
rect 586538 150938 586622 151174
rect 586858 150938 592650 151174
rect -8726 150854 592650 150938
rect -8726 150618 -2934 150854
rect -2698 150618 -2614 150854
rect -2378 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 79610 150854
rect 79846 150618 110330 150854
rect 110566 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 259610 150854
rect 259846 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 586302 150854
rect 586538 150618 586622 150854
rect 586858 150618 592650 150854
rect -8726 150586 592650 150618
rect -8726 147454 592650 147486
rect -8726 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 244250 147454
rect 244486 147218 274970 147454
rect 275206 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 592650 147454
rect -8726 147134 592650 147218
rect -8726 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 244250 147134
rect 244486 146898 274970 147134
rect 275206 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 592650 147134
rect -8726 146866 592650 146898
rect -8726 137494 592650 137526
rect -8726 137258 -8694 137494
rect -8458 137258 -8374 137494
rect -8138 137258 27866 137494
rect 28102 137258 28186 137494
rect 28422 137258 135866 137494
rect 136102 137258 136186 137494
rect 136422 137258 171866 137494
rect 172102 137258 172186 137494
rect 172422 137258 207866 137494
rect 208102 137258 208186 137494
rect 208422 137258 315866 137494
rect 316102 137258 316186 137494
rect 316422 137258 351866 137494
rect 352102 137258 352186 137494
rect 352422 137258 423866 137494
rect 424102 137258 424186 137494
rect 424422 137258 459866 137494
rect 460102 137258 460186 137494
rect 460422 137258 495866 137494
rect 496102 137258 496186 137494
rect 496422 137258 531866 137494
rect 532102 137258 532186 137494
rect 532422 137258 567866 137494
rect 568102 137258 568186 137494
rect 568422 137258 592062 137494
rect 592298 137258 592382 137494
rect 592618 137258 592650 137494
rect -8726 137174 592650 137258
rect -8726 136938 -8694 137174
rect -8458 136938 -8374 137174
rect -8138 136938 27866 137174
rect 28102 136938 28186 137174
rect 28422 136938 135866 137174
rect 136102 136938 136186 137174
rect 136422 136938 171866 137174
rect 172102 136938 172186 137174
rect 172422 136938 207866 137174
rect 208102 136938 208186 137174
rect 208422 136938 315866 137174
rect 316102 136938 316186 137174
rect 316422 136938 351866 137174
rect 352102 136938 352186 137174
rect 352422 136938 423866 137174
rect 424102 136938 424186 137174
rect 424422 136938 459866 137174
rect 460102 136938 460186 137174
rect 460422 136938 495866 137174
rect 496102 136938 496186 137174
rect 496422 136938 531866 137174
rect 532102 136938 532186 137174
rect 532422 136938 567866 137174
rect 568102 136938 568186 137174
rect 568422 136938 592062 137174
rect 592298 136938 592382 137174
rect 592618 136938 592650 137174
rect -8726 136906 592650 136938
rect -8726 133774 592650 133806
rect -8726 133538 -7734 133774
rect -7498 133538 -7414 133774
rect -7178 133538 24146 133774
rect 24382 133538 24466 133774
rect 24702 133538 132146 133774
rect 132382 133538 132466 133774
rect 132702 133538 168146 133774
rect 168382 133538 168466 133774
rect 168702 133538 204146 133774
rect 204382 133538 204466 133774
rect 204702 133538 312146 133774
rect 312382 133538 312466 133774
rect 312702 133538 348146 133774
rect 348382 133538 348466 133774
rect 348702 133538 420146 133774
rect 420382 133538 420466 133774
rect 420702 133538 456146 133774
rect 456382 133538 456466 133774
rect 456702 133538 492146 133774
rect 492382 133538 492466 133774
rect 492702 133538 528146 133774
rect 528382 133538 528466 133774
rect 528702 133538 564146 133774
rect 564382 133538 564466 133774
rect 564702 133538 591102 133774
rect 591338 133538 591422 133774
rect 591658 133538 592650 133774
rect -8726 133454 592650 133538
rect -8726 133218 -7734 133454
rect -7498 133218 -7414 133454
rect -7178 133218 24146 133454
rect 24382 133218 24466 133454
rect 24702 133218 132146 133454
rect 132382 133218 132466 133454
rect 132702 133218 168146 133454
rect 168382 133218 168466 133454
rect 168702 133218 204146 133454
rect 204382 133218 204466 133454
rect 204702 133218 312146 133454
rect 312382 133218 312466 133454
rect 312702 133218 348146 133454
rect 348382 133218 348466 133454
rect 348702 133218 420146 133454
rect 420382 133218 420466 133454
rect 420702 133218 456146 133454
rect 456382 133218 456466 133454
rect 456702 133218 492146 133454
rect 492382 133218 492466 133454
rect 492702 133218 528146 133454
rect 528382 133218 528466 133454
rect 528702 133218 564146 133454
rect 564382 133218 564466 133454
rect 564702 133218 591102 133454
rect 591338 133218 591422 133454
rect 591658 133218 592650 133454
rect -8726 133186 592650 133218
rect -8726 130054 592650 130086
rect -8726 129818 -6774 130054
rect -6538 129818 -6454 130054
rect -6218 129818 20426 130054
rect 20662 129818 20746 130054
rect 20982 129818 56426 130054
rect 56662 129818 56746 130054
rect 56982 129818 128426 130054
rect 128662 129818 128746 130054
rect 128982 129818 164426 130054
rect 164662 129818 164746 130054
rect 164982 129818 200426 130054
rect 200662 129818 200746 130054
rect 200982 129818 236426 130054
rect 236662 129818 236746 130054
rect 236982 129818 272426 130054
rect 272662 129818 272746 130054
rect 272982 129818 308426 130054
rect 308662 129818 308746 130054
rect 308982 129818 344426 130054
rect 344662 129818 344746 130054
rect 344982 129818 416426 130054
rect 416662 129818 416746 130054
rect 416982 129818 452426 130054
rect 452662 129818 452746 130054
rect 452982 129818 488426 130054
rect 488662 129818 488746 130054
rect 488982 129818 524426 130054
rect 524662 129818 524746 130054
rect 524982 129818 560426 130054
rect 560662 129818 560746 130054
rect 560982 129818 590142 130054
rect 590378 129818 590462 130054
rect 590698 129818 592650 130054
rect -8726 129734 592650 129818
rect -8726 129498 -6774 129734
rect -6538 129498 -6454 129734
rect -6218 129498 20426 129734
rect 20662 129498 20746 129734
rect 20982 129498 56426 129734
rect 56662 129498 56746 129734
rect 56982 129498 128426 129734
rect 128662 129498 128746 129734
rect 128982 129498 164426 129734
rect 164662 129498 164746 129734
rect 164982 129498 200426 129734
rect 200662 129498 200746 129734
rect 200982 129498 236426 129734
rect 236662 129498 236746 129734
rect 236982 129498 272426 129734
rect 272662 129498 272746 129734
rect 272982 129498 308426 129734
rect 308662 129498 308746 129734
rect 308982 129498 344426 129734
rect 344662 129498 344746 129734
rect 344982 129498 416426 129734
rect 416662 129498 416746 129734
rect 416982 129498 452426 129734
rect 452662 129498 452746 129734
rect 452982 129498 488426 129734
rect 488662 129498 488746 129734
rect 488982 129498 524426 129734
rect 524662 129498 524746 129734
rect 524982 129498 560426 129734
rect 560662 129498 560746 129734
rect 560982 129498 590142 129734
rect 590378 129498 590462 129734
rect 590698 129498 592650 129734
rect -8726 129466 592650 129498
rect -8726 126334 592650 126366
rect -8726 126098 -5814 126334
rect -5578 126098 -5494 126334
rect -5258 126098 16706 126334
rect 16942 126098 17026 126334
rect 17262 126098 52706 126334
rect 52942 126098 53026 126334
rect 53262 126098 124706 126334
rect 124942 126098 125026 126334
rect 125262 126098 160706 126334
rect 160942 126098 161026 126334
rect 161262 126098 196706 126334
rect 196942 126098 197026 126334
rect 197262 126098 232706 126334
rect 232942 126098 233026 126334
rect 233262 126098 268706 126334
rect 268942 126098 269026 126334
rect 269262 126098 304706 126334
rect 304942 126098 305026 126334
rect 305262 126098 340706 126334
rect 340942 126098 341026 126334
rect 341262 126098 412706 126334
rect 412942 126098 413026 126334
rect 413262 126098 448706 126334
rect 448942 126098 449026 126334
rect 449262 126098 484706 126334
rect 484942 126098 485026 126334
rect 485262 126098 520706 126334
rect 520942 126098 521026 126334
rect 521262 126098 556706 126334
rect 556942 126098 557026 126334
rect 557262 126098 589182 126334
rect 589418 126098 589502 126334
rect 589738 126098 592650 126334
rect -8726 126014 592650 126098
rect -8726 125778 -5814 126014
rect -5578 125778 -5494 126014
rect -5258 125778 16706 126014
rect 16942 125778 17026 126014
rect 17262 125778 52706 126014
rect 52942 125778 53026 126014
rect 53262 125778 124706 126014
rect 124942 125778 125026 126014
rect 125262 125778 160706 126014
rect 160942 125778 161026 126014
rect 161262 125778 196706 126014
rect 196942 125778 197026 126014
rect 197262 125778 232706 126014
rect 232942 125778 233026 126014
rect 233262 125778 268706 126014
rect 268942 125778 269026 126014
rect 269262 125778 304706 126014
rect 304942 125778 305026 126014
rect 305262 125778 340706 126014
rect 340942 125778 341026 126014
rect 341262 125778 412706 126014
rect 412942 125778 413026 126014
rect 413262 125778 448706 126014
rect 448942 125778 449026 126014
rect 449262 125778 484706 126014
rect 484942 125778 485026 126014
rect 485262 125778 520706 126014
rect 520942 125778 521026 126014
rect 521262 125778 556706 126014
rect 556942 125778 557026 126014
rect 557262 125778 589182 126014
rect 589418 125778 589502 126014
rect 589738 125778 592650 126014
rect -8726 125746 592650 125778
rect -8726 122614 592650 122646
rect -8726 122378 -4854 122614
rect -4618 122378 -4534 122614
rect -4298 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 120986 122614
rect 121222 122378 121306 122614
rect 121542 122378 156986 122614
rect 157222 122378 157306 122614
rect 157542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 588222 122614
rect 588458 122378 588542 122614
rect 588778 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -4854 122294
rect -4618 122058 -4534 122294
rect -4298 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 120986 122294
rect 121222 122058 121306 122294
rect 121542 122058 156986 122294
rect 157222 122058 157306 122294
rect 157542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 588222 122294
rect 588458 122058 588542 122294
rect 588778 122058 592650 122294
rect -8726 122026 592650 122058
rect -8726 118894 592650 118926
rect -8726 118658 -3894 118894
rect -3658 118658 -3574 118894
rect -3338 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 81266 118894
rect 81502 118658 81586 118894
rect 81822 118658 117266 118894
rect 117502 118658 117586 118894
rect 117822 118658 153266 118894
rect 153502 118658 153586 118894
rect 153822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 225266 118894
rect 225502 118658 225586 118894
rect 225822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 587262 118894
rect 587498 118658 587582 118894
rect 587818 118658 592650 118894
rect -8726 118574 592650 118658
rect -8726 118338 -3894 118574
rect -3658 118338 -3574 118574
rect -3338 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 81266 118574
rect 81502 118338 81586 118574
rect 81822 118338 117266 118574
rect 117502 118338 117586 118574
rect 117822 118338 153266 118574
rect 153502 118338 153586 118574
rect 153822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 225266 118574
rect 225502 118338 225586 118574
rect 225822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 587262 118574
rect 587498 118338 587582 118574
rect 587818 118338 592650 118574
rect -8726 118306 592650 118338
rect -8726 115174 592650 115206
rect -8726 114938 -2934 115174
rect -2698 114938 -2614 115174
rect -2378 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 77546 115174
rect 77782 114938 77866 115174
rect 78102 114938 113546 115174
rect 113782 114938 113866 115174
rect 114102 114938 149546 115174
rect 149782 114938 149866 115174
rect 150102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 221546 115174
rect 221782 114938 221866 115174
rect 222102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 379610 115174
rect 379846 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 586302 115174
rect 586538 114938 586622 115174
rect 586858 114938 592650 115174
rect -8726 114854 592650 114938
rect -8726 114618 -2934 114854
rect -2698 114618 -2614 114854
rect -2378 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 77546 114854
rect 77782 114618 77866 114854
rect 78102 114618 113546 114854
rect 113782 114618 113866 114854
rect 114102 114618 149546 114854
rect 149782 114618 149866 114854
rect 150102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 221546 114854
rect 221782 114618 221866 114854
rect 222102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 379610 114854
rect 379846 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 586302 114854
rect 586538 114618 586622 114854
rect 586858 114618 592650 114854
rect -8726 114586 592650 114618
rect -8726 111454 592650 111486
rect -8726 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 73826 111454
rect 74062 111218 74146 111454
rect 74382 111218 109826 111454
rect 110062 111218 110146 111454
rect 110382 111218 145826 111454
rect 146062 111218 146146 111454
rect 146382 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 217826 111454
rect 218062 111218 218146 111454
rect 218382 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 364250 111454
rect 364486 111218 394970 111454
rect 395206 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 592650 111454
rect -8726 111134 592650 111218
rect -8726 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 73826 111134
rect 74062 110898 74146 111134
rect 74382 110898 109826 111134
rect 110062 110898 110146 111134
rect 110382 110898 145826 111134
rect 146062 110898 146146 111134
rect 146382 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 217826 111134
rect 218062 110898 218146 111134
rect 218382 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 364250 111134
rect 364486 110898 394970 111134
rect 395206 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 592650 111134
rect -8726 110866 592650 110898
rect -8726 101494 592650 101526
rect -8726 101258 -8694 101494
rect -8458 101258 -8374 101494
rect -8138 101258 27866 101494
rect 28102 101258 28186 101494
rect 28422 101258 63866 101494
rect 64102 101258 64186 101494
rect 64422 101258 99866 101494
rect 100102 101258 100186 101494
rect 100422 101258 135866 101494
rect 136102 101258 136186 101494
rect 136422 101258 171866 101494
rect 172102 101258 172186 101494
rect 172422 101258 207866 101494
rect 208102 101258 208186 101494
rect 208422 101258 243866 101494
rect 244102 101258 244186 101494
rect 244422 101258 279866 101494
rect 280102 101258 280186 101494
rect 280422 101258 315866 101494
rect 316102 101258 316186 101494
rect 316422 101258 351866 101494
rect 352102 101258 352186 101494
rect 352422 101258 423866 101494
rect 424102 101258 424186 101494
rect 424422 101258 459866 101494
rect 460102 101258 460186 101494
rect 460422 101258 495866 101494
rect 496102 101258 496186 101494
rect 496422 101258 531866 101494
rect 532102 101258 532186 101494
rect 532422 101258 567866 101494
rect 568102 101258 568186 101494
rect 568422 101258 592062 101494
rect 592298 101258 592382 101494
rect 592618 101258 592650 101494
rect -8726 101174 592650 101258
rect -8726 100938 -8694 101174
rect -8458 100938 -8374 101174
rect -8138 100938 27866 101174
rect 28102 100938 28186 101174
rect 28422 100938 63866 101174
rect 64102 100938 64186 101174
rect 64422 100938 99866 101174
rect 100102 100938 100186 101174
rect 100422 100938 135866 101174
rect 136102 100938 136186 101174
rect 136422 100938 171866 101174
rect 172102 100938 172186 101174
rect 172422 100938 207866 101174
rect 208102 100938 208186 101174
rect 208422 100938 243866 101174
rect 244102 100938 244186 101174
rect 244422 100938 279866 101174
rect 280102 100938 280186 101174
rect 280422 100938 315866 101174
rect 316102 100938 316186 101174
rect 316422 100938 351866 101174
rect 352102 100938 352186 101174
rect 352422 100938 423866 101174
rect 424102 100938 424186 101174
rect 424422 100938 459866 101174
rect 460102 100938 460186 101174
rect 460422 100938 495866 101174
rect 496102 100938 496186 101174
rect 496422 100938 531866 101174
rect 532102 100938 532186 101174
rect 532422 100938 567866 101174
rect 568102 100938 568186 101174
rect 568422 100938 592062 101174
rect 592298 100938 592382 101174
rect 592618 100938 592650 101174
rect -8726 100906 592650 100938
rect -8726 97774 592650 97806
rect -8726 97538 -7734 97774
rect -7498 97538 -7414 97774
rect -7178 97538 24146 97774
rect 24382 97538 24466 97774
rect 24702 97538 60146 97774
rect 60382 97538 60466 97774
rect 60702 97538 96146 97774
rect 96382 97538 96466 97774
rect 96702 97538 132146 97774
rect 132382 97538 132466 97774
rect 132702 97538 168146 97774
rect 168382 97538 168466 97774
rect 168702 97538 204146 97774
rect 204382 97538 204466 97774
rect 204702 97538 240146 97774
rect 240382 97538 240466 97774
rect 240702 97538 276146 97774
rect 276382 97538 276466 97774
rect 276702 97538 312146 97774
rect 312382 97538 312466 97774
rect 312702 97538 348146 97774
rect 348382 97538 348466 97774
rect 348702 97538 384146 97774
rect 384382 97538 384466 97774
rect 384702 97538 420146 97774
rect 420382 97538 420466 97774
rect 420702 97538 456146 97774
rect 456382 97538 456466 97774
rect 456702 97538 492146 97774
rect 492382 97538 492466 97774
rect 492702 97538 528146 97774
rect 528382 97538 528466 97774
rect 528702 97538 564146 97774
rect 564382 97538 564466 97774
rect 564702 97538 591102 97774
rect 591338 97538 591422 97774
rect 591658 97538 592650 97774
rect -8726 97454 592650 97538
rect -8726 97218 -7734 97454
rect -7498 97218 -7414 97454
rect -7178 97218 24146 97454
rect 24382 97218 24466 97454
rect 24702 97218 60146 97454
rect 60382 97218 60466 97454
rect 60702 97218 96146 97454
rect 96382 97218 96466 97454
rect 96702 97218 132146 97454
rect 132382 97218 132466 97454
rect 132702 97218 168146 97454
rect 168382 97218 168466 97454
rect 168702 97218 204146 97454
rect 204382 97218 204466 97454
rect 204702 97218 240146 97454
rect 240382 97218 240466 97454
rect 240702 97218 276146 97454
rect 276382 97218 276466 97454
rect 276702 97218 312146 97454
rect 312382 97218 312466 97454
rect 312702 97218 348146 97454
rect 348382 97218 348466 97454
rect 348702 97218 384146 97454
rect 384382 97218 384466 97454
rect 384702 97218 420146 97454
rect 420382 97218 420466 97454
rect 420702 97218 456146 97454
rect 456382 97218 456466 97454
rect 456702 97218 492146 97454
rect 492382 97218 492466 97454
rect 492702 97218 528146 97454
rect 528382 97218 528466 97454
rect 528702 97218 564146 97454
rect 564382 97218 564466 97454
rect 564702 97218 591102 97454
rect 591338 97218 591422 97454
rect 591658 97218 592650 97454
rect -8726 97186 592650 97218
rect -8726 94054 592650 94086
rect -8726 93818 -6774 94054
rect -6538 93818 -6454 94054
rect -6218 93818 20426 94054
rect 20662 93818 20746 94054
rect 20982 93818 56426 94054
rect 56662 93818 56746 94054
rect 56982 93818 92426 94054
rect 92662 93818 92746 94054
rect 92982 93818 128426 94054
rect 128662 93818 128746 94054
rect 128982 93818 164426 94054
rect 164662 93818 164746 94054
rect 164982 93818 200426 94054
rect 200662 93818 200746 94054
rect 200982 93818 236426 94054
rect 236662 93818 236746 94054
rect 236982 93818 272426 94054
rect 272662 93818 272746 94054
rect 272982 93818 308426 94054
rect 308662 93818 308746 94054
rect 308982 93818 344426 94054
rect 344662 93818 344746 94054
rect 344982 93818 380426 94054
rect 380662 93818 380746 94054
rect 380982 93818 416426 94054
rect 416662 93818 416746 94054
rect 416982 93818 452426 94054
rect 452662 93818 452746 94054
rect 452982 93818 488426 94054
rect 488662 93818 488746 94054
rect 488982 93818 524426 94054
rect 524662 93818 524746 94054
rect 524982 93818 560426 94054
rect 560662 93818 560746 94054
rect 560982 93818 590142 94054
rect 590378 93818 590462 94054
rect 590698 93818 592650 94054
rect -8726 93734 592650 93818
rect -8726 93498 -6774 93734
rect -6538 93498 -6454 93734
rect -6218 93498 20426 93734
rect 20662 93498 20746 93734
rect 20982 93498 56426 93734
rect 56662 93498 56746 93734
rect 56982 93498 92426 93734
rect 92662 93498 92746 93734
rect 92982 93498 128426 93734
rect 128662 93498 128746 93734
rect 128982 93498 164426 93734
rect 164662 93498 164746 93734
rect 164982 93498 200426 93734
rect 200662 93498 200746 93734
rect 200982 93498 236426 93734
rect 236662 93498 236746 93734
rect 236982 93498 272426 93734
rect 272662 93498 272746 93734
rect 272982 93498 308426 93734
rect 308662 93498 308746 93734
rect 308982 93498 344426 93734
rect 344662 93498 344746 93734
rect 344982 93498 380426 93734
rect 380662 93498 380746 93734
rect 380982 93498 416426 93734
rect 416662 93498 416746 93734
rect 416982 93498 452426 93734
rect 452662 93498 452746 93734
rect 452982 93498 488426 93734
rect 488662 93498 488746 93734
rect 488982 93498 524426 93734
rect 524662 93498 524746 93734
rect 524982 93498 560426 93734
rect 560662 93498 560746 93734
rect 560982 93498 590142 93734
rect 590378 93498 590462 93734
rect 590698 93498 592650 93734
rect -8726 93466 592650 93498
rect -8726 90334 592650 90366
rect -8726 90098 -5814 90334
rect -5578 90098 -5494 90334
rect -5258 90098 16706 90334
rect 16942 90098 17026 90334
rect 17262 90098 52706 90334
rect 52942 90098 53026 90334
rect 53262 90098 88706 90334
rect 88942 90098 89026 90334
rect 89262 90098 124706 90334
rect 124942 90098 125026 90334
rect 125262 90098 160706 90334
rect 160942 90098 161026 90334
rect 161262 90098 196706 90334
rect 196942 90098 197026 90334
rect 197262 90098 232706 90334
rect 232942 90098 233026 90334
rect 233262 90098 268706 90334
rect 268942 90098 269026 90334
rect 269262 90098 304706 90334
rect 304942 90098 305026 90334
rect 305262 90098 340706 90334
rect 340942 90098 341026 90334
rect 341262 90098 376706 90334
rect 376942 90098 377026 90334
rect 377262 90098 412706 90334
rect 412942 90098 413026 90334
rect 413262 90098 448706 90334
rect 448942 90098 449026 90334
rect 449262 90098 484706 90334
rect 484942 90098 485026 90334
rect 485262 90098 520706 90334
rect 520942 90098 521026 90334
rect 521262 90098 556706 90334
rect 556942 90098 557026 90334
rect 557262 90098 589182 90334
rect 589418 90098 589502 90334
rect 589738 90098 592650 90334
rect -8726 90014 592650 90098
rect -8726 89778 -5814 90014
rect -5578 89778 -5494 90014
rect -5258 89778 16706 90014
rect 16942 89778 17026 90014
rect 17262 89778 52706 90014
rect 52942 89778 53026 90014
rect 53262 89778 88706 90014
rect 88942 89778 89026 90014
rect 89262 89778 124706 90014
rect 124942 89778 125026 90014
rect 125262 89778 160706 90014
rect 160942 89778 161026 90014
rect 161262 89778 196706 90014
rect 196942 89778 197026 90014
rect 197262 89778 232706 90014
rect 232942 89778 233026 90014
rect 233262 89778 268706 90014
rect 268942 89778 269026 90014
rect 269262 89778 304706 90014
rect 304942 89778 305026 90014
rect 305262 89778 340706 90014
rect 340942 89778 341026 90014
rect 341262 89778 376706 90014
rect 376942 89778 377026 90014
rect 377262 89778 412706 90014
rect 412942 89778 413026 90014
rect 413262 89778 448706 90014
rect 448942 89778 449026 90014
rect 449262 89778 484706 90014
rect 484942 89778 485026 90014
rect 485262 89778 520706 90014
rect 520942 89778 521026 90014
rect 521262 89778 556706 90014
rect 556942 89778 557026 90014
rect 557262 89778 589182 90014
rect 589418 89778 589502 90014
rect 589738 89778 592650 90014
rect -8726 89746 592650 89778
rect -8726 86614 592650 86646
rect -8726 86378 -4854 86614
rect -4618 86378 -4534 86614
rect -4298 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 588222 86614
rect 588458 86378 588542 86614
rect 588778 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -4854 86294
rect -4618 86058 -4534 86294
rect -4298 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 588222 86294
rect 588458 86058 588542 86294
rect 588778 86058 592650 86294
rect -8726 86026 592650 86058
rect -8726 82894 592650 82926
rect -8726 82658 -3894 82894
rect -3658 82658 -3574 82894
rect -3338 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 587262 82894
rect 587498 82658 587582 82894
rect 587818 82658 592650 82894
rect -8726 82574 592650 82658
rect -8726 82338 -3894 82574
rect -3658 82338 -3574 82574
rect -3338 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 587262 82574
rect 587498 82338 587582 82574
rect 587818 82338 592650 82574
rect -8726 82306 592650 82338
rect -8726 79174 592650 79206
rect -8726 78938 -2934 79174
rect -2698 78938 -2614 79174
rect -2378 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 59174 79174
rect 59410 78938 67362 79174
rect 67598 78938 75550 79174
rect 75786 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 83738 79174
rect 83974 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 586302 79174
rect 586538 78938 586622 79174
rect 586858 78938 592650 79174
rect -8726 78854 592650 78938
rect -8726 78618 -2934 78854
rect -2698 78618 -2614 78854
rect -2378 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 59174 78854
rect 59410 78618 67362 78854
rect 67598 78618 75550 78854
rect 75786 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 83738 78854
rect 83974 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 586302 78854
rect 586538 78618 586622 78854
rect 586858 78618 592650 78854
rect -8726 78586 592650 78618
rect -8726 75454 592650 75486
rect -8726 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 55080 75454
rect 55316 75218 63268 75454
rect 63504 75218 71456 75454
rect 71692 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 79644 75454
rect 79880 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 592650 75454
rect -8726 75134 592650 75218
rect -8726 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 55080 75134
rect 55316 74898 63268 75134
rect 63504 74898 71456 75134
rect 71692 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 79644 75134
rect 79880 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 592650 75134
rect -8726 74866 592650 74898
rect -8726 65494 592650 65526
rect -8726 65258 -8694 65494
rect -8458 65258 -8374 65494
rect -8138 65258 27866 65494
rect 28102 65258 28186 65494
rect 28422 65258 63866 65494
rect 64102 65258 64186 65494
rect 64422 65258 99866 65494
rect 100102 65258 100186 65494
rect 100422 65258 135866 65494
rect 136102 65258 136186 65494
rect 136422 65258 171866 65494
rect 172102 65258 172186 65494
rect 172422 65258 207866 65494
rect 208102 65258 208186 65494
rect 208422 65258 243866 65494
rect 244102 65258 244186 65494
rect 244422 65258 279866 65494
rect 280102 65258 280186 65494
rect 280422 65258 315866 65494
rect 316102 65258 316186 65494
rect 316422 65258 351866 65494
rect 352102 65258 352186 65494
rect 352422 65258 387866 65494
rect 388102 65258 388186 65494
rect 388422 65258 423866 65494
rect 424102 65258 424186 65494
rect 424422 65258 459866 65494
rect 460102 65258 460186 65494
rect 460422 65258 495866 65494
rect 496102 65258 496186 65494
rect 496422 65258 531866 65494
rect 532102 65258 532186 65494
rect 532422 65258 567866 65494
rect 568102 65258 568186 65494
rect 568422 65258 592062 65494
rect 592298 65258 592382 65494
rect 592618 65258 592650 65494
rect -8726 65174 592650 65258
rect -8726 64938 -8694 65174
rect -8458 64938 -8374 65174
rect -8138 64938 27866 65174
rect 28102 64938 28186 65174
rect 28422 64938 63866 65174
rect 64102 64938 64186 65174
rect 64422 64938 99866 65174
rect 100102 64938 100186 65174
rect 100422 64938 135866 65174
rect 136102 64938 136186 65174
rect 136422 64938 171866 65174
rect 172102 64938 172186 65174
rect 172422 64938 207866 65174
rect 208102 64938 208186 65174
rect 208422 64938 243866 65174
rect 244102 64938 244186 65174
rect 244422 64938 279866 65174
rect 280102 64938 280186 65174
rect 280422 64938 315866 65174
rect 316102 64938 316186 65174
rect 316422 64938 351866 65174
rect 352102 64938 352186 65174
rect 352422 64938 387866 65174
rect 388102 64938 388186 65174
rect 388422 64938 423866 65174
rect 424102 64938 424186 65174
rect 424422 64938 459866 65174
rect 460102 64938 460186 65174
rect 460422 64938 495866 65174
rect 496102 64938 496186 65174
rect 496422 64938 531866 65174
rect 532102 64938 532186 65174
rect 532422 64938 567866 65174
rect 568102 64938 568186 65174
rect 568422 64938 592062 65174
rect 592298 64938 592382 65174
rect 592618 64938 592650 65174
rect -8726 64906 592650 64938
rect -8726 61774 592650 61806
rect -8726 61538 -7734 61774
rect -7498 61538 -7414 61774
rect -7178 61538 24146 61774
rect 24382 61538 24466 61774
rect 24702 61538 60146 61774
rect 60382 61538 60466 61774
rect 60702 61538 96146 61774
rect 96382 61538 96466 61774
rect 96702 61538 132146 61774
rect 132382 61538 132466 61774
rect 132702 61538 168146 61774
rect 168382 61538 168466 61774
rect 168702 61538 204146 61774
rect 204382 61538 204466 61774
rect 204702 61538 240146 61774
rect 240382 61538 240466 61774
rect 240702 61538 276146 61774
rect 276382 61538 276466 61774
rect 276702 61538 312146 61774
rect 312382 61538 312466 61774
rect 312702 61538 348146 61774
rect 348382 61538 348466 61774
rect 348702 61538 384146 61774
rect 384382 61538 384466 61774
rect 384702 61538 420146 61774
rect 420382 61538 420466 61774
rect 420702 61538 456146 61774
rect 456382 61538 456466 61774
rect 456702 61538 492146 61774
rect 492382 61538 492466 61774
rect 492702 61538 528146 61774
rect 528382 61538 528466 61774
rect 528702 61538 564146 61774
rect 564382 61538 564466 61774
rect 564702 61538 591102 61774
rect 591338 61538 591422 61774
rect 591658 61538 592650 61774
rect -8726 61454 592650 61538
rect -8726 61218 -7734 61454
rect -7498 61218 -7414 61454
rect -7178 61218 24146 61454
rect 24382 61218 24466 61454
rect 24702 61218 60146 61454
rect 60382 61218 60466 61454
rect 60702 61218 96146 61454
rect 96382 61218 96466 61454
rect 96702 61218 132146 61454
rect 132382 61218 132466 61454
rect 132702 61218 168146 61454
rect 168382 61218 168466 61454
rect 168702 61218 204146 61454
rect 204382 61218 204466 61454
rect 204702 61218 240146 61454
rect 240382 61218 240466 61454
rect 240702 61218 276146 61454
rect 276382 61218 276466 61454
rect 276702 61218 312146 61454
rect 312382 61218 312466 61454
rect 312702 61218 348146 61454
rect 348382 61218 348466 61454
rect 348702 61218 384146 61454
rect 384382 61218 384466 61454
rect 384702 61218 420146 61454
rect 420382 61218 420466 61454
rect 420702 61218 456146 61454
rect 456382 61218 456466 61454
rect 456702 61218 492146 61454
rect 492382 61218 492466 61454
rect 492702 61218 528146 61454
rect 528382 61218 528466 61454
rect 528702 61218 564146 61454
rect 564382 61218 564466 61454
rect 564702 61218 591102 61454
rect 591338 61218 591422 61454
rect 591658 61218 592650 61454
rect -8726 61186 592650 61218
rect -8726 58054 592650 58086
rect -8726 57818 -6774 58054
rect -6538 57818 -6454 58054
rect -6218 57818 20426 58054
rect 20662 57818 20746 58054
rect 20982 57818 56426 58054
rect 56662 57818 56746 58054
rect 56982 57818 92426 58054
rect 92662 57818 92746 58054
rect 92982 57818 128426 58054
rect 128662 57818 128746 58054
rect 128982 57818 164426 58054
rect 164662 57818 164746 58054
rect 164982 57818 200426 58054
rect 200662 57818 200746 58054
rect 200982 57818 236426 58054
rect 236662 57818 236746 58054
rect 236982 57818 272426 58054
rect 272662 57818 272746 58054
rect 272982 57818 308426 58054
rect 308662 57818 308746 58054
rect 308982 57818 344426 58054
rect 344662 57818 344746 58054
rect 344982 57818 380426 58054
rect 380662 57818 380746 58054
rect 380982 57818 416426 58054
rect 416662 57818 416746 58054
rect 416982 57818 452426 58054
rect 452662 57818 452746 58054
rect 452982 57818 488426 58054
rect 488662 57818 488746 58054
rect 488982 57818 524426 58054
rect 524662 57818 524746 58054
rect 524982 57818 560426 58054
rect 560662 57818 560746 58054
rect 560982 57818 590142 58054
rect 590378 57818 590462 58054
rect 590698 57818 592650 58054
rect -8726 57734 592650 57818
rect -8726 57498 -6774 57734
rect -6538 57498 -6454 57734
rect -6218 57498 20426 57734
rect 20662 57498 20746 57734
rect 20982 57498 56426 57734
rect 56662 57498 56746 57734
rect 56982 57498 92426 57734
rect 92662 57498 92746 57734
rect 92982 57498 128426 57734
rect 128662 57498 128746 57734
rect 128982 57498 164426 57734
rect 164662 57498 164746 57734
rect 164982 57498 200426 57734
rect 200662 57498 200746 57734
rect 200982 57498 236426 57734
rect 236662 57498 236746 57734
rect 236982 57498 272426 57734
rect 272662 57498 272746 57734
rect 272982 57498 308426 57734
rect 308662 57498 308746 57734
rect 308982 57498 344426 57734
rect 344662 57498 344746 57734
rect 344982 57498 380426 57734
rect 380662 57498 380746 57734
rect 380982 57498 416426 57734
rect 416662 57498 416746 57734
rect 416982 57498 452426 57734
rect 452662 57498 452746 57734
rect 452982 57498 488426 57734
rect 488662 57498 488746 57734
rect 488982 57498 524426 57734
rect 524662 57498 524746 57734
rect 524982 57498 560426 57734
rect 560662 57498 560746 57734
rect 560982 57498 590142 57734
rect 590378 57498 590462 57734
rect 590698 57498 592650 57734
rect -8726 57466 592650 57498
rect -8726 54334 592650 54366
rect -8726 54098 -5814 54334
rect -5578 54098 -5494 54334
rect -5258 54098 16706 54334
rect 16942 54098 17026 54334
rect 17262 54098 52706 54334
rect 52942 54098 53026 54334
rect 53262 54098 88706 54334
rect 88942 54098 89026 54334
rect 89262 54098 124706 54334
rect 124942 54098 125026 54334
rect 125262 54098 160706 54334
rect 160942 54098 161026 54334
rect 161262 54098 196706 54334
rect 196942 54098 197026 54334
rect 197262 54098 232706 54334
rect 232942 54098 233026 54334
rect 233262 54098 268706 54334
rect 268942 54098 269026 54334
rect 269262 54098 304706 54334
rect 304942 54098 305026 54334
rect 305262 54098 340706 54334
rect 340942 54098 341026 54334
rect 341262 54098 376706 54334
rect 376942 54098 377026 54334
rect 377262 54098 412706 54334
rect 412942 54098 413026 54334
rect 413262 54098 448706 54334
rect 448942 54098 449026 54334
rect 449262 54098 484706 54334
rect 484942 54098 485026 54334
rect 485262 54098 520706 54334
rect 520942 54098 521026 54334
rect 521262 54098 556706 54334
rect 556942 54098 557026 54334
rect 557262 54098 589182 54334
rect 589418 54098 589502 54334
rect 589738 54098 592650 54334
rect -8726 54014 592650 54098
rect -8726 53778 -5814 54014
rect -5578 53778 -5494 54014
rect -5258 53778 16706 54014
rect 16942 53778 17026 54014
rect 17262 53778 52706 54014
rect 52942 53778 53026 54014
rect 53262 53778 88706 54014
rect 88942 53778 89026 54014
rect 89262 53778 124706 54014
rect 124942 53778 125026 54014
rect 125262 53778 160706 54014
rect 160942 53778 161026 54014
rect 161262 53778 196706 54014
rect 196942 53778 197026 54014
rect 197262 53778 232706 54014
rect 232942 53778 233026 54014
rect 233262 53778 268706 54014
rect 268942 53778 269026 54014
rect 269262 53778 304706 54014
rect 304942 53778 305026 54014
rect 305262 53778 340706 54014
rect 340942 53778 341026 54014
rect 341262 53778 376706 54014
rect 376942 53778 377026 54014
rect 377262 53778 412706 54014
rect 412942 53778 413026 54014
rect 413262 53778 448706 54014
rect 448942 53778 449026 54014
rect 449262 53778 484706 54014
rect 484942 53778 485026 54014
rect 485262 53778 520706 54014
rect 520942 53778 521026 54014
rect 521262 53778 556706 54014
rect 556942 53778 557026 54014
rect 557262 53778 589182 54014
rect 589418 53778 589502 54014
rect 589738 53778 592650 54014
rect -8726 53746 592650 53778
rect -8726 50614 592650 50646
rect -8726 50378 -4854 50614
rect -4618 50378 -4534 50614
rect -4298 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 588222 50614
rect 588458 50378 588542 50614
rect 588778 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -4854 50294
rect -4618 50058 -4534 50294
rect -4298 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 588222 50294
rect 588458 50058 588542 50294
rect 588778 50058 592650 50294
rect -8726 50026 592650 50058
rect -8726 46894 592650 46926
rect -8726 46658 -3894 46894
rect -3658 46658 -3574 46894
rect -3338 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 587262 46894
rect 587498 46658 587582 46894
rect 587818 46658 592650 46894
rect -8726 46574 592650 46658
rect -8726 46338 -3894 46574
rect -3658 46338 -3574 46574
rect -3338 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 587262 46574
rect 587498 46338 587582 46574
rect 587818 46338 592650 46574
rect -8726 46306 592650 46338
rect -8726 43174 592650 43206
rect -8726 42938 -2934 43174
rect -2698 42938 -2614 43174
rect -2378 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 586302 43174
rect 586538 42938 586622 43174
rect 586858 42938 592650 43174
rect -8726 42854 592650 42938
rect -8726 42618 -2934 42854
rect -2698 42618 -2614 42854
rect -2378 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 586302 42854
rect 586538 42618 586622 42854
rect 586858 42618 592650 42854
rect -8726 42586 592650 42618
rect -8726 39454 592650 39486
rect -8726 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 592650 39454
rect -8726 39134 592650 39218
rect -8726 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 592650 39134
rect -8726 38866 592650 38898
rect -8726 29494 592650 29526
rect -8726 29258 -8694 29494
rect -8458 29258 -8374 29494
rect -8138 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 63866 29494
rect 64102 29258 64186 29494
rect 64422 29258 99866 29494
rect 100102 29258 100186 29494
rect 100422 29258 135866 29494
rect 136102 29258 136186 29494
rect 136422 29258 171866 29494
rect 172102 29258 172186 29494
rect 172422 29258 207866 29494
rect 208102 29258 208186 29494
rect 208422 29258 243866 29494
rect 244102 29258 244186 29494
rect 244422 29258 279866 29494
rect 280102 29258 280186 29494
rect 280422 29258 315866 29494
rect 316102 29258 316186 29494
rect 316422 29258 351866 29494
rect 352102 29258 352186 29494
rect 352422 29258 387866 29494
rect 388102 29258 388186 29494
rect 388422 29258 423866 29494
rect 424102 29258 424186 29494
rect 424422 29258 459866 29494
rect 460102 29258 460186 29494
rect 460422 29258 495866 29494
rect 496102 29258 496186 29494
rect 496422 29258 531866 29494
rect 532102 29258 532186 29494
rect 532422 29258 567866 29494
rect 568102 29258 568186 29494
rect 568422 29258 592062 29494
rect 592298 29258 592382 29494
rect 592618 29258 592650 29494
rect -8726 29174 592650 29258
rect -8726 28938 -8694 29174
rect -8458 28938 -8374 29174
rect -8138 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 63866 29174
rect 64102 28938 64186 29174
rect 64422 28938 99866 29174
rect 100102 28938 100186 29174
rect 100422 28938 135866 29174
rect 136102 28938 136186 29174
rect 136422 28938 171866 29174
rect 172102 28938 172186 29174
rect 172422 28938 207866 29174
rect 208102 28938 208186 29174
rect 208422 28938 243866 29174
rect 244102 28938 244186 29174
rect 244422 28938 279866 29174
rect 280102 28938 280186 29174
rect 280422 28938 315866 29174
rect 316102 28938 316186 29174
rect 316422 28938 351866 29174
rect 352102 28938 352186 29174
rect 352422 28938 387866 29174
rect 388102 28938 388186 29174
rect 388422 28938 423866 29174
rect 424102 28938 424186 29174
rect 424422 28938 459866 29174
rect 460102 28938 460186 29174
rect 460422 28938 495866 29174
rect 496102 28938 496186 29174
rect 496422 28938 531866 29174
rect 532102 28938 532186 29174
rect 532422 28938 567866 29174
rect 568102 28938 568186 29174
rect 568422 28938 592062 29174
rect 592298 28938 592382 29174
rect 592618 28938 592650 29174
rect -8726 28906 592650 28938
rect -8726 25774 592650 25806
rect -8726 25538 -7734 25774
rect -7498 25538 -7414 25774
rect -7178 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 60146 25774
rect 60382 25538 60466 25774
rect 60702 25538 96146 25774
rect 96382 25538 96466 25774
rect 96702 25538 132146 25774
rect 132382 25538 132466 25774
rect 132702 25538 168146 25774
rect 168382 25538 168466 25774
rect 168702 25538 204146 25774
rect 204382 25538 204466 25774
rect 204702 25538 240146 25774
rect 240382 25538 240466 25774
rect 240702 25538 276146 25774
rect 276382 25538 276466 25774
rect 276702 25538 312146 25774
rect 312382 25538 312466 25774
rect 312702 25538 348146 25774
rect 348382 25538 348466 25774
rect 348702 25538 384146 25774
rect 384382 25538 384466 25774
rect 384702 25538 420146 25774
rect 420382 25538 420466 25774
rect 420702 25538 456146 25774
rect 456382 25538 456466 25774
rect 456702 25538 492146 25774
rect 492382 25538 492466 25774
rect 492702 25538 528146 25774
rect 528382 25538 528466 25774
rect 528702 25538 564146 25774
rect 564382 25538 564466 25774
rect 564702 25538 591102 25774
rect 591338 25538 591422 25774
rect 591658 25538 592650 25774
rect -8726 25454 592650 25538
rect -8726 25218 -7734 25454
rect -7498 25218 -7414 25454
rect -7178 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 60146 25454
rect 60382 25218 60466 25454
rect 60702 25218 96146 25454
rect 96382 25218 96466 25454
rect 96702 25218 132146 25454
rect 132382 25218 132466 25454
rect 132702 25218 168146 25454
rect 168382 25218 168466 25454
rect 168702 25218 204146 25454
rect 204382 25218 204466 25454
rect 204702 25218 240146 25454
rect 240382 25218 240466 25454
rect 240702 25218 276146 25454
rect 276382 25218 276466 25454
rect 276702 25218 312146 25454
rect 312382 25218 312466 25454
rect 312702 25218 348146 25454
rect 348382 25218 348466 25454
rect 348702 25218 384146 25454
rect 384382 25218 384466 25454
rect 384702 25218 420146 25454
rect 420382 25218 420466 25454
rect 420702 25218 456146 25454
rect 456382 25218 456466 25454
rect 456702 25218 492146 25454
rect 492382 25218 492466 25454
rect 492702 25218 528146 25454
rect 528382 25218 528466 25454
rect 528702 25218 564146 25454
rect 564382 25218 564466 25454
rect 564702 25218 591102 25454
rect 591338 25218 591422 25454
rect 591658 25218 592650 25454
rect -8726 25186 592650 25218
rect -8726 22054 592650 22086
rect -8726 21818 -6774 22054
rect -6538 21818 -6454 22054
rect -6218 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 56426 22054
rect 56662 21818 56746 22054
rect 56982 21818 92426 22054
rect 92662 21818 92746 22054
rect 92982 21818 128426 22054
rect 128662 21818 128746 22054
rect 128982 21818 164426 22054
rect 164662 21818 164746 22054
rect 164982 21818 200426 22054
rect 200662 21818 200746 22054
rect 200982 21818 236426 22054
rect 236662 21818 236746 22054
rect 236982 21818 272426 22054
rect 272662 21818 272746 22054
rect 272982 21818 308426 22054
rect 308662 21818 308746 22054
rect 308982 21818 344426 22054
rect 344662 21818 344746 22054
rect 344982 21818 380426 22054
rect 380662 21818 380746 22054
rect 380982 21818 416426 22054
rect 416662 21818 416746 22054
rect 416982 21818 452426 22054
rect 452662 21818 452746 22054
rect 452982 21818 488426 22054
rect 488662 21818 488746 22054
rect 488982 21818 524426 22054
rect 524662 21818 524746 22054
rect 524982 21818 560426 22054
rect 560662 21818 560746 22054
rect 560982 21818 590142 22054
rect 590378 21818 590462 22054
rect 590698 21818 592650 22054
rect -8726 21734 592650 21818
rect -8726 21498 -6774 21734
rect -6538 21498 -6454 21734
rect -6218 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 56426 21734
rect 56662 21498 56746 21734
rect 56982 21498 92426 21734
rect 92662 21498 92746 21734
rect 92982 21498 128426 21734
rect 128662 21498 128746 21734
rect 128982 21498 164426 21734
rect 164662 21498 164746 21734
rect 164982 21498 200426 21734
rect 200662 21498 200746 21734
rect 200982 21498 236426 21734
rect 236662 21498 236746 21734
rect 236982 21498 272426 21734
rect 272662 21498 272746 21734
rect 272982 21498 308426 21734
rect 308662 21498 308746 21734
rect 308982 21498 344426 21734
rect 344662 21498 344746 21734
rect 344982 21498 380426 21734
rect 380662 21498 380746 21734
rect 380982 21498 416426 21734
rect 416662 21498 416746 21734
rect 416982 21498 452426 21734
rect 452662 21498 452746 21734
rect 452982 21498 488426 21734
rect 488662 21498 488746 21734
rect 488982 21498 524426 21734
rect 524662 21498 524746 21734
rect 524982 21498 560426 21734
rect 560662 21498 560746 21734
rect 560982 21498 590142 21734
rect 590378 21498 590462 21734
rect 590698 21498 592650 21734
rect -8726 21466 592650 21498
rect -8726 18334 592650 18366
rect -8726 18098 -5814 18334
rect -5578 18098 -5494 18334
rect -5258 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 52706 18334
rect 52942 18098 53026 18334
rect 53262 18098 88706 18334
rect 88942 18098 89026 18334
rect 89262 18098 124706 18334
rect 124942 18098 125026 18334
rect 125262 18098 160706 18334
rect 160942 18098 161026 18334
rect 161262 18098 196706 18334
rect 196942 18098 197026 18334
rect 197262 18098 232706 18334
rect 232942 18098 233026 18334
rect 233262 18098 268706 18334
rect 268942 18098 269026 18334
rect 269262 18098 304706 18334
rect 304942 18098 305026 18334
rect 305262 18098 340706 18334
rect 340942 18098 341026 18334
rect 341262 18098 376706 18334
rect 376942 18098 377026 18334
rect 377262 18098 412706 18334
rect 412942 18098 413026 18334
rect 413262 18098 448706 18334
rect 448942 18098 449026 18334
rect 449262 18098 484706 18334
rect 484942 18098 485026 18334
rect 485262 18098 520706 18334
rect 520942 18098 521026 18334
rect 521262 18098 556706 18334
rect 556942 18098 557026 18334
rect 557262 18098 589182 18334
rect 589418 18098 589502 18334
rect 589738 18098 592650 18334
rect -8726 18014 592650 18098
rect -8726 17778 -5814 18014
rect -5578 17778 -5494 18014
rect -5258 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 52706 18014
rect 52942 17778 53026 18014
rect 53262 17778 88706 18014
rect 88942 17778 89026 18014
rect 89262 17778 124706 18014
rect 124942 17778 125026 18014
rect 125262 17778 160706 18014
rect 160942 17778 161026 18014
rect 161262 17778 196706 18014
rect 196942 17778 197026 18014
rect 197262 17778 232706 18014
rect 232942 17778 233026 18014
rect 233262 17778 268706 18014
rect 268942 17778 269026 18014
rect 269262 17778 304706 18014
rect 304942 17778 305026 18014
rect 305262 17778 340706 18014
rect 340942 17778 341026 18014
rect 341262 17778 376706 18014
rect 376942 17778 377026 18014
rect 377262 17778 412706 18014
rect 412942 17778 413026 18014
rect 413262 17778 448706 18014
rect 448942 17778 449026 18014
rect 449262 17778 484706 18014
rect 484942 17778 485026 18014
rect 485262 17778 520706 18014
rect 520942 17778 521026 18014
rect 521262 17778 556706 18014
rect 556942 17778 557026 18014
rect 557262 17778 589182 18014
rect 589418 17778 589502 18014
rect 589738 17778 592650 18014
rect -8726 17746 592650 17778
rect -8726 14614 592650 14646
rect -8726 14378 -4854 14614
rect -4618 14378 -4534 14614
rect -4298 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 588222 14614
rect 588458 14378 588542 14614
rect 588778 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -4854 14294
rect -4618 14058 -4534 14294
rect -4298 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 588222 14294
rect 588458 14058 588542 14294
rect 588778 14058 592650 14294
rect -8726 14026 592650 14058
rect -8726 10894 592650 10926
rect -8726 10658 -3894 10894
rect -3658 10658 -3574 10894
rect -3338 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 587262 10894
rect 587498 10658 587582 10894
rect 587818 10658 592650 10894
rect -8726 10574 592650 10658
rect -8726 10338 -3894 10574
rect -3658 10338 -3574 10574
rect -3338 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 587262 10574
rect 587498 10338 587582 10574
rect 587818 10338 592650 10574
rect -8726 10306 592650 10338
rect -8726 7174 592650 7206
rect -8726 6938 -2934 7174
rect -2698 6938 -2614 7174
rect -2378 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 586302 7174
rect 586538 6938 586622 7174
rect 586858 6938 592650 7174
rect -8726 6854 592650 6938
rect -8726 6618 -2934 6854
rect -2698 6618 -2614 6854
rect -2378 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 586302 6854
rect 586538 6618 586622 6854
rect 586858 6618 592650 6854
rect -8726 6586 592650 6618
rect -8726 3454 592650 3486
rect -8726 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 592650 3454
rect -8726 3134 592650 3218
rect -8726 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 592650 3134
rect -8726 2866 592650 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 5546 -1306
rect 5782 -1542 5866 -1306
rect 6102 -1542 41546 -1306
rect 41782 -1542 41866 -1306
rect 42102 -1542 77546 -1306
rect 77782 -1542 77866 -1306
rect 78102 -1542 113546 -1306
rect 113782 -1542 113866 -1306
rect 114102 -1542 149546 -1306
rect 149782 -1542 149866 -1306
rect 150102 -1542 185546 -1306
rect 185782 -1542 185866 -1306
rect 186102 -1542 221546 -1306
rect 221782 -1542 221866 -1306
rect 222102 -1542 257546 -1306
rect 257782 -1542 257866 -1306
rect 258102 -1542 293546 -1306
rect 293782 -1542 293866 -1306
rect 294102 -1542 329546 -1306
rect 329782 -1542 329866 -1306
rect 330102 -1542 365546 -1306
rect 365782 -1542 365866 -1306
rect 366102 -1542 401546 -1306
rect 401782 -1542 401866 -1306
rect 402102 -1542 437546 -1306
rect 437782 -1542 437866 -1306
rect 438102 -1542 473546 -1306
rect 473782 -1542 473866 -1306
rect 474102 -1542 509546 -1306
rect 509782 -1542 509866 -1306
rect 510102 -1542 545546 -1306
rect 545782 -1542 545866 -1306
rect 546102 -1542 581546 -1306
rect 581782 -1542 581866 -1306
rect 582102 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 5546 -1626
rect 5782 -1862 5866 -1626
rect 6102 -1862 41546 -1626
rect 41782 -1862 41866 -1626
rect 42102 -1862 77546 -1626
rect 77782 -1862 77866 -1626
rect 78102 -1862 113546 -1626
rect 113782 -1862 113866 -1626
rect 114102 -1862 149546 -1626
rect 149782 -1862 149866 -1626
rect 150102 -1862 185546 -1626
rect 185782 -1862 185866 -1626
rect 186102 -1862 221546 -1626
rect 221782 -1862 221866 -1626
rect 222102 -1862 257546 -1626
rect 257782 -1862 257866 -1626
rect 258102 -1862 293546 -1626
rect 293782 -1862 293866 -1626
rect 294102 -1862 329546 -1626
rect 329782 -1862 329866 -1626
rect 330102 -1862 365546 -1626
rect 365782 -1862 365866 -1626
rect 366102 -1862 401546 -1626
rect 401782 -1862 401866 -1626
rect 402102 -1862 437546 -1626
rect 437782 -1862 437866 -1626
rect 438102 -1862 473546 -1626
rect 473782 -1862 473866 -1626
rect 474102 -1862 509546 -1626
rect 509782 -1862 509866 -1626
rect 510102 -1862 545546 -1626
rect 545782 -1862 545866 -1626
rect 546102 -1862 581546 -1626
rect 581782 -1862 581866 -1626
rect 582102 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 9266 -2266
rect 9502 -2502 9586 -2266
rect 9822 -2502 45266 -2266
rect 45502 -2502 45586 -2266
rect 45822 -2502 81266 -2266
rect 81502 -2502 81586 -2266
rect 81822 -2502 117266 -2266
rect 117502 -2502 117586 -2266
rect 117822 -2502 153266 -2266
rect 153502 -2502 153586 -2266
rect 153822 -2502 189266 -2266
rect 189502 -2502 189586 -2266
rect 189822 -2502 225266 -2266
rect 225502 -2502 225586 -2266
rect 225822 -2502 261266 -2266
rect 261502 -2502 261586 -2266
rect 261822 -2502 297266 -2266
rect 297502 -2502 297586 -2266
rect 297822 -2502 333266 -2266
rect 333502 -2502 333586 -2266
rect 333822 -2502 369266 -2266
rect 369502 -2502 369586 -2266
rect 369822 -2502 405266 -2266
rect 405502 -2502 405586 -2266
rect 405822 -2502 441266 -2266
rect 441502 -2502 441586 -2266
rect 441822 -2502 477266 -2266
rect 477502 -2502 477586 -2266
rect 477822 -2502 513266 -2266
rect 513502 -2502 513586 -2266
rect 513822 -2502 549266 -2266
rect 549502 -2502 549586 -2266
rect 549822 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 9266 -2586
rect 9502 -2822 9586 -2586
rect 9822 -2822 45266 -2586
rect 45502 -2822 45586 -2586
rect 45822 -2822 81266 -2586
rect 81502 -2822 81586 -2586
rect 81822 -2822 117266 -2586
rect 117502 -2822 117586 -2586
rect 117822 -2822 153266 -2586
rect 153502 -2822 153586 -2586
rect 153822 -2822 189266 -2586
rect 189502 -2822 189586 -2586
rect 189822 -2822 225266 -2586
rect 225502 -2822 225586 -2586
rect 225822 -2822 261266 -2586
rect 261502 -2822 261586 -2586
rect 261822 -2822 297266 -2586
rect 297502 -2822 297586 -2586
rect 297822 -2822 333266 -2586
rect 333502 -2822 333586 -2586
rect 333822 -2822 369266 -2586
rect 369502 -2822 369586 -2586
rect 369822 -2822 405266 -2586
rect 405502 -2822 405586 -2586
rect 405822 -2822 441266 -2586
rect 441502 -2822 441586 -2586
rect 441822 -2822 477266 -2586
rect 477502 -2822 477586 -2586
rect 477822 -2822 513266 -2586
rect 513502 -2822 513586 -2586
rect 513822 -2822 549266 -2586
rect 549502 -2822 549586 -2586
rect 549822 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 12986 -3226
rect 13222 -3462 13306 -3226
rect 13542 -3462 48986 -3226
rect 49222 -3462 49306 -3226
rect 49542 -3462 84986 -3226
rect 85222 -3462 85306 -3226
rect 85542 -3462 120986 -3226
rect 121222 -3462 121306 -3226
rect 121542 -3462 156986 -3226
rect 157222 -3462 157306 -3226
rect 157542 -3462 192986 -3226
rect 193222 -3462 193306 -3226
rect 193542 -3462 228986 -3226
rect 229222 -3462 229306 -3226
rect 229542 -3462 264986 -3226
rect 265222 -3462 265306 -3226
rect 265542 -3462 300986 -3226
rect 301222 -3462 301306 -3226
rect 301542 -3462 336986 -3226
rect 337222 -3462 337306 -3226
rect 337542 -3462 372986 -3226
rect 373222 -3462 373306 -3226
rect 373542 -3462 408986 -3226
rect 409222 -3462 409306 -3226
rect 409542 -3462 444986 -3226
rect 445222 -3462 445306 -3226
rect 445542 -3462 480986 -3226
rect 481222 -3462 481306 -3226
rect 481542 -3462 516986 -3226
rect 517222 -3462 517306 -3226
rect 517542 -3462 552986 -3226
rect 553222 -3462 553306 -3226
rect 553542 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 12986 -3546
rect 13222 -3782 13306 -3546
rect 13542 -3782 48986 -3546
rect 49222 -3782 49306 -3546
rect 49542 -3782 84986 -3546
rect 85222 -3782 85306 -3546
rect 85542 -3782 120986 -3546
rect 121222 -3782 121306 -3546
rect 121542 -3782 156986 -3546
rect 157222 -3782 157306 -3546
rect 157542 -3782 192986 -3546
rect 193222 -3782 193306 -3546
rect 193542 -3782 228986 -3546
rect 229222 -3782 229306 -3546
rect 229542 -3782 264986 -3546
rect 265222 -3782 265306 -3546
rect 265542 -3782 300986 -3546
rect 301222 -3782 301306 -3546
rect 301542 -3782 336986 -3546
rect 337222 -3782 337306 -3546
rect 337542 -3782 372986 -3546
rect 373222 -3782 373306 -3546
rect 373542 -3782 408986 -3546
rect 409222 -3782 409306 -3546
rect 409542 -3782 444986 -3546
rect 445222 -3782 445306 -3546
rect 445542 -3782 480986 -3546
rect 481222 -3782 481306 -3546
rect 481542 -3782 516986 -3546
rect 517222 -3782 517306 -3546
rect 517542 -3782 552986 -3546
rect 553222 -3782 553306 -3546
rect 553542 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 16706 -4186
rect 16942 -4422 17026 -4186
rect 17262 -4422 52706 -4186
rect 52942 -4422 53026 -4186
rect 53262 -4422 88706 -4186
rect 88942 -4422 89026 -4186
rect 89262 -4422 124706 -4186
rect 124942 -4422 125026 -4186
rect 125262 -4422 160706 -4186
rect 160942 -4422 161026 -4186
rect 161262 -4422 196706 -4186
rect 196942 -4422 197026 -4186
rect 197262 -4422 232706 -4186
rect 232942 -4422 233026 -4186
rect 233262 -4422 268706 -4186
rect 268942 -4422 269026 -4186
rect 269262 -4422 304706 -4186
rect 304942 -4422 305026 -4186
rect 305262 -4422 340706 -4186
rect 340942 -4422 341026 -4186
rect 341262 -4422 376706 -4186
rect 376942 -4422 377026 -4186
rect 377262 -4422 412706 -4186
rect 412942 -4422 413026 -4186
rect 413262 -4422 448706 -4186
rect 448942 -4422 449026 -4186
rect 449262 -4422 484706 -4186
rect 484942 -4422 485026 -4186
rect 485262 -4422 520706 -4186
rect 520942 -4422 521026 -4186
rect 521262 -4422 556706 -4186
rect 556942 -4422 557026 -4186
rect 557262 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 16706 -4506
rect 16942 -4742 17026 -4506
rect 17262 -4742 52706 -4506
rect 52942 -4742 53026 -4506
rect 53262 -4742 88706 -4506
rect 88942 -4742 89026 -4506
rect 89262 -4742 124706 -4506
rect 124942 -4742 125026 -4506
rect 125262 -4742 160706 -4506
rect 160942 -4742 161026 -4506
rect 161262 -4742 196706 -4506
rect 196942 -4742 197026 -4506
rect 197262 -4742 232706 -4506
rect 232942 -4742 233026 -4506
rect 233262 -4742 268706 -4506
rect 268942 -4742 269026 -4506
rect 269262 -4742 304706 -4506
rect 304942 -4742 305026 -4506
rect 305262 -4742 340706 -4506
rect 340942 -4742 341026 -4506
rect 341262 -4742 376706 -4506
rect 376942 -4742 377026 -4506
rect 377262 -4742 412706 -4506
rect 412942 -4742 413026 -4506
rect 413262 -4742 448706 -4506
rect 448942 -4742 449026 -4506
rect 449262 -4742 484706 -4506
rect 484942 -4742 485026 -4506
rect 485262 -4742 520706 -4506
rect 520942 -4742 521026 -4506
rect 521262 -4742 556706 -4506
rect 556942 -4742 557026 -4506
rect 557262 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 20426 -5146
rect 20662 -5382 20746 -5146
rect 20982 -5382 56426 -5146
rect 56662 -5382 56746 -5146
rect 56982 -5382 92426 -5146
rect 92662 -5382 92746 -5146
rect 92982 -5382 128426 -5146
rect 128662 -5382 128746 -5146
rect 128982 -5382 164426 -5146
rect 164662 -5382 164746 -5146
rect 164982 -5382 200426 -5146
rect 200662 -5382 200746 -5146
rect 200982 -5382 236426 -5146
rect 236662 -5382 236746 -5146
rect 236982 -5382 272426 -5146
rect 272662 -5382 272746 -5146
rect 272982 -5382 308426 -5146
rect 308662 -5382 308746 -5146
rect 308982 -5382 344426 -5146
rect 344662 -5382 344746 -5146
rect 344982 -5382 380426 -5146
rect 380662 -5382 380746 -5146
rect 380982 -5382 416426 -5146
rect 416662 -5382 416746 -5146
rect 416982 -5382 452426 -5146
rect 452662 -5382 452746 -5146
rect 452982 -5382 488426 -5146
rect 488662 -5382 488746 -5146
rect 488982 -5382 524426 -5146
rect 524662 -5382 524746 -5146
rect 524982 -5382 560426 -5146
rect 560662 -5382 560746 -5146
rect 560982 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 20426 -5466
rect 20662 -5702 20746 -5466
rect 20982 -5702 56426 -5466
rect 56662 -5702 56746 -5466
rect 56982 -5702 92426 -5466
rect 92662 -5702 92746 -5466
rect 92982 -5702 128426 -5466
rect 128662 -5702 128746 -5466
rect 128982 -5702 164426 -5466
rect 164662 -5702 164746 -5466
rect 164982 -5702 200426 -5466
rect 200662 -5702 200746 -5466
rect 200982 -5702 236426 -5466
rect 236662 -5702 236746 -5466
rect 236982 -5702 272426 -5466
rect 272662 -5702 272746 -5466
rect 272982 -5702 308426 -5466
rect 308662 -5702 308746 -5466
rect 308982 -5702 344426 -5466
rect 344662 -5702 344746 -5466
rect 344982 -5702 380426 -5466
rect 380662 -5702 380746 -5466
rect 380982 -5702 416426 -5466
rect 416662 -5702 416746 -5466
rect 416982 -5702 452426 -5466
rect 452662 -5702 452746 -5466
rect 452982 -5702 488426 -5466
rect 488662 -5702 488746 -5466
rect 488982 -5702 524426 -5466
rect 524662 -5702 524746 -5466
rect 524982 -5702 560426 -5466
rect 560662 -5702 560746 -5466
rect 560982 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 24146 -6106
rect 24382 -6342 24466 -6106
rect 24702 -6342 60146 -6106
rect 60382 -6342 60466 -6106
rect 60702 -6342 96146 -6106
rect 96382 -6342 96466 -6106
rect 96702 -6342 132146 -6106
rect 132382 -6342 132466 -6106
rect 132702 -6342 168146 -6106
rect 168382 -6342 168466 -6106
rect 168702 -6342 204146 -6106
rect 204382 -6342 204466 -6106
rect 204702 -6342 240146 -6106
rect 240382 -6342 240466 -6106
rect 240702 -6342 276146 -6106
rect 276382 -6342 276466 -6106
rect 276702 -6342 312146 -6106
rect 312382 -6342 312466 -6106
rect 312702 -6342 348146 -6106
rect 348382 -6342 348466 -6106
rect 348702 -6342 384146 -6106
rect 384382 -6342 384466 -6106
rect 384702 -6342 420146 -6106
rect 420382 -6342 420466 -6106
rect 420702 -6342 456146 -6106
rect 456382 -6342 456466 -6106
rect 456702 -6342 492146 -6106
rect 492382 -6342 492466 -6106
rect 492702 -6342 528146 -6106
rect 528382 -6342 528466 -6106
rect 528702 -6342 564146 -6106
rect 564382 -6342 564466 -6106
rect 564702 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 24146 -6426
rect 24382 -6662 24466 -6426
rect 24702 -6662 60146 -6426
rect 60382 -6662 60466 -6426
rect 60702 -6662 96146 -6426
rect 96382 -6662 96466 -6426
rect 96702 -6662 132146 -6426
rect 132382 -6662 132466 -6426
rect 132702 -6662 168146 -6426
rect 168382 -6662 168466 -6426
rect 168702 -6662 204146 -6426
rect 204382 -6662 204466 -6426
rect 204702 -6662 240146 -6426
rect 240382 -6662 240466 -6426
rect 240702 -6662 276146 -6426
rect 276382 -6662 276466 -6426
rect 276702 -6662 312146 -6426
rect 312382 -6662 312466 -6426
rect 312702 -6662 348146 -6426
rect 348382 -6662 348466 -6426
rect 348702 -6662 384146 -6426
rect 384382 -6662 384466 -6426
rect 384702 -6662 420146 -6426
rect 420382 -6662 420466 -6426
rect 420702 -6662 456146 -6426
rect 456382 -6662 456466 -6426
rect 456702 -6662 492146 -6426
rect 492382 -6662 492466 -6426
rect 492702 -6662 528146 -6426
rect 528382 -6662 528466 -6426
rect 528702 -6662 564146 -6426
rect 564382 -6662 564466 -6426
rect 564702 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 27866 -7066
rect 28102 -7302 28186 -7066
rect 28422 -7302 63866 -7066
rect 64102 -7302 64186 -7066
rect 64422 -7302 99866 -7066
rect 100102 -7302 100186 -7066
rect 100422 -7302 135866 -7066
rect 136102 -7302 136186 -7066
rect 136422 -7302 171866 -7066
rect 172102 -7302 172186 -7066
rect 172422 -7302 207866 -7066
rect 208102 -7302 208186 -7066
rect 208422 -7302 243866 -7066
rect 244102 -7302 244186 -7066
rect 244422 -7302 279866 -7066
rect 280102 -7302 280186 -7066
rect 280422 -7302 315866 -7066
rect 316102 -7302 316186 -7066
rect 316422 -7302 351866 -7066
rect 352102 -7302 352186 -7066
rect 352422 -7302 387866 -7066
rect 388102 -7302 388186 -7066
rect 388422 -7302 423866 -7066
rect 424102 -7302 424186 -7066
rect 424422 -7302 459866 -7066
rect 460102 -7302 460186 -7066
rect 460422 -7302 495866 -7066
rect 496102 -7302 496186 -7066
rect 496422 -7302 531866 -7066
rect 532102 -7302 532186 -7066
rect 532422 -7302 567866 -7066
rect 568102 -7302 568186 -7066
rect 568422 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 27866 -7386
rect 28102 -7622 28186 -7386
rect 28422 -7622 63866 -7386
rect 64102 -7622 64186 -7386
rect 64422 -7622 99866 -7386
rect 100102 -7622 100186 -7386
rect 100422 -7622 135866 -7386
rect 136102 -7622 136186 -7386
rect 136422 -7622 171866 -7386
rect 172102 -7622 172186 -7386
rect 172422 -7622 207866 -7386
rect 208102 -7622 208186 -7386
rect 208422 -7622 243866 -7386
rect 244102 -7622 244186 -7386
rect 244422 -7622 279866 -7386
rect 280102 -7622 280186 -7386
rect 280422 -7622 315866 -7386
rect 316102 -7622 316186 -7386
rect 316422 -7622 351866 -7386
rect 352102 -7622 352186 -7386
rect 352422 -7622 387866 -7386
rect 388102 -7622 388186 -7386
rect 388422 -7622 423866 -7386
rect 424102 -7622 424186 -7386
rect 424422 -7622 459866 -7386
rect 460102 -7622 460186 -7386
rect 460422 -7622 495866 -7386
rect 496102 -7622 496186 -7386
rect 496422 -7622 531866 -7386
rect 532102 -7622 532186 -7386
rect 532422 -7622 567866 -7386
rect 568102 -7622 568186 -7386
rect 568422 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use ci2406_z80  ci2406_z80
timestamp 0
transform 1 0 50000 0 1 240000
box 0 0 60000 60000
use execution_unit  eu0
timestamp 0
transform 1 0 60000 0 1 560000
box 0 0 75000 75000
use execution_unit  eu1
timestamp 0
transform 1 0 180000 0 1 560000
box 0 0 75000 75000
use execution_unit  eu2
timestamp 0
transform 1 0 300000 0 1 560000
box 0 0 75000 75000
use icache  icache
timestamp 0
transform 1 0 360000 0 1 180000
box 0 0 140000 170000
use multiplexer  multiplexer
timestamp 0
transform 1 0 240000 0 1 120000
box 0 0 40000 220000
use scrapcpu  scrapcpu
timestamp 0
transform 1 0 490000 0 1 600000
box 0 0 50000 55000
use unused_tie  unused_tie
timestamp 0
transform 1 0 50000 0 1 50000
box 0 0 35000 35000
use vliw  vliw
timestamp 0
transform 1 0 60000 0 1 390000
box 0 0 440000 130000
use wrapped_6502  wrapped_6502
timestamp 0
transform 1 0 360000 0 1 100000
box 0 0 45000 45000
use wrapped_as1802  wrapped_as1802
timestamp 0
transform 1 0 60000 0 1 120000
box 0 0 65000 65000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 1794 -7654 2414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 37794 -7654 38414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 -7654 74414 120207 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 183305 74414 238167 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 300449 74414 558575 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 73794 633233 74414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 -7654 110414 119988 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 300449 110414 389988 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 109794 634540 110414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 145794 -7654 146414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 -7654 182414 558575 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 181794 633233 182414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 -7654 218414 388711 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 217794 633233 218414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 -7654 254414 132447 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 253794 633233 254414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 -7654 290414 388711 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 289794 522121 290414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 -7654 326414 388711 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 325794 633233 326414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 -7654 362414 100479 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 361794 633233 362414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 -7654 398414 179799 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 397794 522121 398414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 -7654 434414 179799 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 433794 522121 434414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 -7654 470414 179799 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 469794 522121 470414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 -7654 506414 600207 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 505794 654737 506414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 541794 -7654 542414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 577794 -7654 578414 711590 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 2866 592650 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 38866 592650 39486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 74866 592650 75486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 110866 592650 111486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 146866 592650 147486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 182866 592650 183486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 218866 592650 219486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 254866 592650 255486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 290866 592650 291486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 326866 592650 327486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 362866 592650 363486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 398866 592650 399486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 434866 592650 435486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 470866 592650 471486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 506866 592650 507486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 542866 592650 543486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 578866 592650 579486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 614866 592650 615486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 650866 592650 651486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 686866 592650 687486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 9234 -7654 9854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 45234 -7654 45854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 -7654 81854 120207 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 183305 81854 238167 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 300449 81854 558575 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 81234 633233 81854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 -7654 117854 558575 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 117234 633233 117854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 153234 -7654 153854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 -7654 189854 558575 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 189234 633233 189854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 -7654 225854 388711 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 225234 633233 225854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 -7654 261854 132447 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 261234 522121 261854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 -7654 297854 388711 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 297234 522121 297854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 -7654 333854 388711 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 333234 633233 333854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 -7654 369854 100479 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 369234 633233 369854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 -7654 405854 179799 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 405234 522121 405854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 -7654 441854 179799 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 441234 522121 441854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 -7654 477854 179799 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 477234 522121 477854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 -7654 513854 600207 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 513234 654737 513854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 549234 -7654 549854 711590 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 10306 592650 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 46306 592650 46926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 82306 592650 82926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 118306 592650 118926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 154306 592650 154926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 190306 592650 190926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 226306 592650 226926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 262306 592650 262926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 298306 592650 298926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 334306 592650 334926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 370306 592650 370926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 406306 592650 406926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 442306 592650 442926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 478306 592650 478926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 514306 592650 514926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 550306 592650 550926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 586306 592650 586926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 622306 592650 622926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 658306 592650 658926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -8726 694306 592650 694926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 16674 -7654 17294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 52674 -7654 53294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 -7654 89294 120207 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 183305 89294 238167 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 300449 89294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 88674 633233 89294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 -7654 125294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 124674 633233 125294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 160674 -7654 161294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 -7654 197294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 196674 633233 197294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 -7654 233294 388711 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 522121 233294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 232674 633233 233294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 -7654 269294 132447 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 336713 269294 388711 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 268674 522121 269294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 -7654 305294 388711 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 522121 305294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 304674 633233 305294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 -7654 341294 388711 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 522121 341294 558575 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 340674 633233 341294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 -7654 377294 100479 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 376674 522121 377294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 -7654 413294 179799 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 412674 522121 413294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 -7654 449294 179799 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 448674 522121 449294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 -7654 485294 179799 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 484674 522121 485294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 -7654 521294 600207 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 520674 654737 521294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 556674 -7654 557294 711590 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 17746 592650 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 53746 592650 54366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 89746 592650 90366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 125746 592650 126366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 161746 592650 162366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 197746 592650 198366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 233746 592650 234366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 269746 592650 270366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 305746 592650 306366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 341746 592650 342366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 377746 592650 378366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 413746 592650 414366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 449746 592650 450366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 485746 592650 486366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 521746 592650 522366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 557746 592650 558366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 593746 592650 594366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 629746 592650 630366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -8726 665746 592650 666366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 24114 -7654 24734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 -7654 60734 120207 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 300449 60734 558575 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 60114 633233 60734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 -7654 96734 120207 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 300449 96734 558575 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 96114 633233 96734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 -7654 132734 558575 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 132114 633233 132734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 168114 -7654 168734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 -7654 204734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 204114 633233 204734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 -7654 240734 132447 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 336713 240734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 240114 633233 240734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 -7654 276734 132447 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 336713 276734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 276114 522121 276734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 -7654 312734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 312114 633233 312734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 -7654 348734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 348114 633233 348734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 -7654 384734 100479 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 348433 384734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 384114 522121 384734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 -7654 420734 179799 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 348433 420734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 420114 522121 420734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 -7654 456734 179799 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 349740 456734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 456114 522121 456734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 -7654 492734 179799 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 348433 492734 388711 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 492114 522121 492734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 -7654 528734 600207 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 528114 654737 528734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 564114 -7654 564734 711590 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 25186 592650 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 61186 592650 61806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 97186 592650 97806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 133186 592650 133806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 169186 592650 169806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 205186 592650 205806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 241186 592650 241806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 277186 592650 277806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 313186 592650 313806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 349186 592650 349806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 385186 592650 385806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 421186 592650 421806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 457186 592650 457806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 493186 592650 493806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 529186 592650 529806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 565186 592650 565806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 601186 592650 601806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 637186 592650 637806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -8726 673186 592650 673806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 20394 -7654 21014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 56394 -7654 57014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 -7654 93014 120207 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 183305 93014 238167 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 300449 93014 558575 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 92394 633233 93014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 -7654 129014 558575 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 128394 633233 129014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 164394 -7654 165014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 -7654 201014 388711 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 200394 633233 201014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 -7654 237014 388711 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 236394 633233 237014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 -7654 273014 132447 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 336713 273014 388711 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 272394 522121 273014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 -7654 309014 388711 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 308394 633233 309014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 -7654 345014 388711 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 344394 633233 345014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 -7654 381014 100479 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 380394 522121 381014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 -7654 417014 179799 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 416394 522121 417014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 -7654 453014 179799 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 452394 522121 453014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 -7654 489014 179799 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 488394 522121 489014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 -7654 525014 599988 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 524394 654956 525014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 560394 -7654 561014 711590 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 21466 592650 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 57466 592650 58086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 93466 592650 94086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 129466 592650 130086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 165466 592650 166086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 201466 592650 202086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 237466 592650 238086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 273466 592650 274086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 309466 592650 310086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 345466 592650 346086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 381466 592650 382086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 417466 592650 418086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 453466 592650 454086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 489466 592650 490086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 525466 592650 526086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 561466 592650 562086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 597466 592650 598086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 633466 592650 634086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -8726 669466 592650 670086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 27834 -7654 28454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 -7654 64454 119988 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 300449 64454 389988 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 63834 634540 64454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 -7654 100454 120207 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 300449 100454 558575 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 99834 633233 100454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 135834 -7654 136454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 -7654 172454 389988 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 171834 519484 172454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 -7654 208454 388711 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 207834 633233 208454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 -7654 244454 119988 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 243834 633233 244454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 -7654 280454 132447 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 279834 522121 280454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 -7654 316454 388711 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 315834 633233 316454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 -7654 352454 388711 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 351834 633233 352454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 -7654 388454 100479 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 387834 522121 388454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 -7654 424454 179799 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 423834 522121 424454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 -7654 460454 179799 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 459834 522121 460454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 -7654 496454 179799 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 522121 496454 600207 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 495834 654737 496454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 -7654 532454 600207 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 531834 654737 532454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 567834 -7654 568454 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 28906 592650 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 64906 592650 65526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 100906 592650 101526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 136906 592650 137526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 172906 592650 173526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 208906 592650 209526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 244906 592650 245526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 280906 592650 281526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 316906 592650 317526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 352906 592650 353526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 388906 592650 389526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 424906 592650 425526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 460906 592650 461526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 496906 592650 497526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 532906 592650 533526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 568906 592650 569526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 604906 592650 605526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 640906 592650 641526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 676906 592650 677526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 5514 -7654 6134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 41514 -7654 42134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 -7654 78134 120207 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 183305 78134 238167 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 300449 78134 558575 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 77514 633233 78134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 -7654 114134 120207 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 183305 114134 558575 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 113514 633233 114134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 149514 -7654 150134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 -7654 186134 558575 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 185514 633233 186134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 -7654 222134 388711 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 221514 633233 222134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 -7654 258134 132447 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 257514 522121 258134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 -7654 294134 388711 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 293514 522121 294134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 -7654 330134 388711 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 329514 633233 330134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 -7654 366134 100479 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 365514 634540 366134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 -7654 402134 179799 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 401514 522121 402134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 -7654 438134 179799 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 437514 522121 438134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 -7654 474134 179799 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 473514 522121 474134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 -7654 510134 599988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 509514 654956 510134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 545514 -7654 546134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 581514 -7654 582134 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 6586 592650 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 42586 592650 43206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 78586 592650 79206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 114586 592650 115206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 150586 592650 151206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 186586 592650 187206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 222586 592650 223206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 258586 592650 259206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 294586 592650 295206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 330586 592650 331206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 366586 592650 367206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 402586 592650 403206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 438586 592650 439206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 474586 592650 475206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 510586 592650 511206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 546586 592650 547206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 582586 592650 583206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 618586 592650 619206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 654586 592650 655206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 690586 592650 691206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 12954 -7654 13574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 48954 -7654 49574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 -7654 85574 120207 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 183305 85574 238167 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 300449 85574 558575 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 84954 633233 85574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 -7654 121574 558575 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 120954 633233 121574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 156954 -7654 157574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 -7654 193574 558575 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 192954 633233 193574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 -7654 229574 388711 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 228954 633233 229574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 -7654 265574 132447 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 336713 265574 388711 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 264954 522121 265574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 -7654 301574 388711 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 300954 633233 301574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 -7654 337574 388711 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 336954 633233 337574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 -7654 373574 100479 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 372954 633233 373574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 -7654 409574 179799 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 408954 522121 409574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 -7654 445574 179799 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 444954 522121 445574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 -7654 481574 179799 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 480954 522121 481574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 -7654 517574 600207 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 516954 654737 517574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 552954 -7654 553574 711590 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 14026 592650 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 50026 592650 50646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 86026 592650 86646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 122026 592650 122646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 158026 592650 158646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 194026 592650 194646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 230026 592650 230646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 266026 592650 266646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 302026 592650 302646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 338026 592650 338646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 374026 592650 374646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 410026 592650 410646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 446026 592650 446646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 482026 592650 482646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 518026 592650 518646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 554026 592650 554646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 590026 592650 590646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 626026 592650 626646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 662026 592650 662646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -8726 698026 592650 698646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
